// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 3 2022 09:53:11

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VR_READY_VCCINAUX,
    V33A_ENn,
    V1P8A_EN,
    VDDQ_EN,
    VCCST_OVERRIDE_3V3,
    V5S_OK,
    SLP_S3n,
    SLP_S0n,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    GPIO_FPGA_SoC_2,
    VCCIN_VR_PROCHOT_FPGA,
    SLP_SUSn,
    CPU_C10_GATE_N,
    VCCST_EN,
    V33DSW_OK,
    TPM_GPIO,
    SUSWARN_N,
    PLTRSTn,
    GPIO_FPGA_SoC_4,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    FPGA_OSC,
    VCCST_PWRGD,
    SYS_PWROK,
    SPI_FP_IO2,
    SATAXPCIE1_FPGA,
    GPIO_FPGA_EXP_1,
    VCCINAUX_VR_PROCHOT_FPGA,
    VCCINAUX_VR_PE,
    HDA_SDO_ATP,
    GPIO_FPGA_EXP_2,
    VPP_EN,
    VDDQ_OK,
    SUSACK_N,
    SLP_S4n,
    VCCST_CPU_OK,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    GPIO_FPGA_SoC_1,
    DSW_PWROK,
    V5A_EN,
    GPIO_FPGA_SoC_3,
    VR_PROCHOT_FPGA_OUT_N,
    VPP_OK,
    VCCIN_VR_PE,
    VCCIN_EN,
    SOC_SPKR,
    SLP_S5n,
    V12_MAIN_MON,
    SPI_FP_IO3,
    SATAXPCIE0_FPGA,
    V33A_OK,
    PCH_PWROK,
    FPGA_SLP_WLAN_N);

    input VR_READY_VCCINAUX;
    output V33A_ENn;
    output V1P8A_EN;
    output VDDQ_EN;
    input VCCST_OVERRIDE_3V3;
    input V5S_OK;
    input SLP_S3n;
    input SLP_S0n;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input GPIO_FPGA_SoC_2;
    input VCCIN_VR_PROCHOT_FPGA;
    input SLP_SUSn;
    input CPU_C10_GATE_N;
    output VCCST_EN;
    input V33DSW_OK;
    input TPM_GPIO;
    output SUSWARN_N;
    input PLTRSTn;
    input GPIO_FPGA_SoC_4;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output SYS_PWROK;
    input SPI_FP_IO2;
    input SATAXPCIE1_FPGA;
    input GPIO_FPGA_EXP_1;
    input VCCINAUX_VR_PROCHOT_FPGA;
    output VCCINAUX_VR_PE;
    output HDA_SDO_ATP;
    input GPIO_FPGA_EXP_2;
    output VPP_EN;
    input VDDQ_OK;
    input SUSACK_N;
    input SLP_S4n;
    input VCCST_CPU_OK;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input GPIO_FPGA_SoC_1;
    output DSW_PWROK;
    output V5A_EN;
    input GPIO_FPGA_SoC_3;
    input VR_PROCHOT_FPGA_OUT_N;
    input VPP_OK;
    output VCCIN_VR_PE;
    output VCCIN_EN;
    input SOC_SPKR;
    input SLP_S5n;
    input V12_MAIN_MON;
    input SPI_FP_IO3;
    input SATAXPCIE0_FPGA;
    input V33A_OK;
    output PCH_PWROK;
    input FPGA_SLP_WLAN_N;

    wire N__34571;
    wire N__34570;
    wire N__34569;
    wire N__34562;
    wire N__34561;
    wire N__34560;
    wire N__34553;
    wire N__34552;
    wire N__34551;
    wire N__34544;
    wire N__34543;
    wire N__34542;
    wire N__34535;
    wire N__34534;
    wire N__34533;
    wire N__34526;
    wire N__34525;
    wire N__34524;
    wire N__34517;
    wire N__34516;
    wire N__34515;
    wire N__34508;
    wire N__34507;
    wire N__34506;
    wire N__34499;
    wire N__34498;
    wire N__34497;
    wire N__34490;
    wire N__34489;
    wire N__34488;
    wire N__34481;
    wire N__34480;
    wire N__34479;
    wire N__34472;
    wire N__34471;
    wire N__34470;
    wire N__34463;
    wire N__34462;
    wire N__34461;
    wire N__34454;
    wire N__34453;
    wire N__34452;
    wire N__34445;
    wire N__34444;
    wire N__34443;
    wire N__34436;
    wire N__34435;
    wire N__34434;
    wire N__34427;
    wire N__34426;
    wire N__34425;
    wire N__34418;
    wire N__34417;
    wire N__34416;
    wire N__34409;
    wire N__34408;
    wire N__34407;
    wire N__34400;
    wire N__34399;
    wire N__34398;
    wire N__34391;
    wire N__34390;
    wire N__34389;
    wire N__34382;
    wire N__34381;
    wire N__34380;
    wire N__34373;
    wire N__34372;
    wire N__34371;
    wire N__34364;
    wire N__34363;
    wire N__34362;
    wire N__34355;
    wire N__34354;
    wire N__34353;
    wire N__34346;
    wire N__34345;
    wire N__34344;
    wire N__34337;
    wire N__34336;
    wire N__34335;
    wire N__34328;
    wire N__34327;
    wire N__34326;
    wire N__34319;
    wire N__34318;
    wire N__34317;
    wire N__34310;
    wire N__34309;
    wire N__34308;
    wire N__34301;
    wire N__34300;
    wire N__34299;
    wire N__34292;
    wire N__34291;
    wire N__34290;
    wire N__34283;
    wire N__34282;
    wire N__34281;
    wire N__34274;
    wire N__34273;
    wire N__34272;
    wire N__34265;
    wire N__34264;
    wire N__34263;
    wire N__34256;
    wire N__34255;
    wire N__34254;
    wire N__34247;
    wire N__34246;
    wire N__34245;
    wire N__34238;
    wire N__34237;
    wire N__34236;
    wire N__34229;
    wire N__34228;
    wire N__34227;
    wire N__34220;
    wire N__34219;
    wire N__34218;
    wire N__34211;
    wire N__34210;
    wire N__34209;
    wire N__34202;
    wire N__34201;
    wire N__34200;
    wire N__34193;
    wire N__34192;
    wire N__34191;
    wire N__34184;
    wire N__34183;
    wire N__34182;
    wire N__34175;
    wire N__34174;
    wire N__34173;
    wire N__34166;
    wire N__34165;
    wire N__34164;
    wire N__34157;
    wire N__34156;
    wire N__34155;
    wire N__34148;
    wire N__34147;
    wire N__34146;
    wire N__34139;
    wire N__34138;
    wire N__34137;
    wire N__34130;
    wire N__34129;
    wire N__34128;
    wire N__34121;
    wire N__34120;
    wire N__34119;
    wire N__34112;
    wire N__34111;
    wire N__34110;
    wire N__34103;
    wire N__34102;
    wire N__34101;
    wire N__34094;
    wire N__34093;
    wire N__34092;
    wire N__34085;
    wire N__34084;
    wire N__34083;
    wire N__34076;
    wire N__34075;
    wire N__34074;
    wire N__34067;
    wire N__34066;
    wire N__34065;
    wire N__34058;
    wire N__34057;
    wire N__34056;
    wire N__34049;
    wire N__34048;
    wire N__34047;
    wire N__34030;
    wire N__34027;
    wire N__34026;
    wire N__34025;
    wire N__34024;
    wire N__34023;
    wire N__34022;
    wire N__34021;
    wire N__34020;
    wire N__34011;
    wire N__34004;
    wire N__34003;
    wire N__34002;
    wire N__34001;
    wire N__34000;
    wire N__33999;
    wire N__33998;
    wire N__33995;
    wire N__33990;
    wire N__33989;
    wire N__33988;
    wire N__33987;
    wire N__33986;
    wire N__33985;
    wire N__33984;
    wire N__33983;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33965;
    wire N__33962;
    wire N__33953;
    wire N__33946;
    wire N__33945;
    wire N__33944;
    wire N__33943;
    wire N__33942;
    wire N__33941;
    wire N__33940;
    wire N__33939;
    wire N__33934;
    wire N__33933;
    wire N__33932;
    wire N__33931;
    wire N__33930;
    wire N__33929;
    wire N__33928;
    wire N__33925;
    wire N__33924;
    wire N__33923;
    wire N__33914;
    wire N__33911;
    wire N__33910;
    wire N__33909;
    wire N__33902;
    wire N__33901;
    wire N__33900;
    wire N__33893;
    wire N__33890;
    wire N__33887;
    wire N__33884;
    wire N__33881;
    wire N__33880;
    wire N__33879;
    wire N__33878;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33862;
    wire N__33861;
    wire N__33858;
    wire N__33855;
    wire N__33852;
    wire N__33851;
    wire N__33850;
    wire N__33849;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33827;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33810;
    wire N__33803;
    wire N__33798;
    wire N__33795;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33779;
    wire N__33770;
    wire N__33765;
    wire N__33762;
    wire N__33751;
    wire N__33748;
    wire N__33727;
    wire N__33726;
    wire N__33725;
    wire N__33724;
    wire N__33723;
    wire N__33722;
    wire N__33721;
    wire N__33720;
    wire N__33719;
    wire N__33718;
    wire N__33717;
    wire N__33716;
    wire N__33715;
    wire N__33714;
    wire N__33711;
    wire N__33710;
    wire N__33707;
    wire N__33706;
    wire N__33705;
    wire N__33702;
    wire N__33701;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33691;
    wire N__33688;
    wire N__33685;
    wire N__33684;
    wire N__33681;
    wire N__33678;
    wire N__33677;
    wire N__33676;
    wire N__33675;
    wire N__33666;
    wire N__33657;
    wire N__33656;
    wire N__33655;
    wire N__33654;
    wire N__33651;
    wire N__33650;
    wire N__33649;
    wire N__33642;
    wire N__33637;
    wire N__33634;
    wire N__33623;
    wire N__33622;
    wire N__33619;
    wire N__33618;
    wire N__33615;
    wire N__33614;
    wire N__33613;
    wire N__33610;
    wire N__33609;
    wire N__33608;
    wire N__33607;
    wire N__33606;
    wire N__33603;
    wire N__33600;
    wire N__33587;
    wire N__33584;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33562;
    wire N__33551;
    wire N__33548;
    wire N__33545;
    wire N__33540;
    wire N__33523;
    wire N__33522;
    wire N__33521;
    wire N__33520;
    wire N__33519;
    wire N__33518;
    wire N__33517;
    wire N__33514;
    wire N__33513;
    wire N__33512;
    wire N__33511;
    wire N__33510;
    wire N__33509;
    wire N__33506;
    wire N__33503;
    wire N__33498;
    wire N__33497;
    wire N__33496;
    wire N__33495;
    wire N__33494;
    wire N__33493;
    wire N__33492;
    wire N__33491;
    wire N__33490;
    wire N__33489;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33481;
    wire N__33478;
    wire N__33475;
    wire N__33466;
    wire N__33461;
    wire N__33460;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33452;
    wire N__33449;
    wire N__33442;
    wire N__33437;
    wire N__33436;
    wire N__33433;
    wire N__33430;
    wire N__33429;
    wire N__33428;
    wire N__33427;
    wire N__33418;
    wire N__33409;
    wire N__33406;
    wire N__33405;
    wire N__33402;
    wire N__33401;
    wire N__33396;
    wire N__33395;
    wire N__33392;
    wire N__33391;
    wire N__33388;
    wire N__33383;
    wire N__33370;
    wire N__33367;
    wire N__33366;
    wire N__33365;
    wire N__33364;
    wire N__33363;
    wire N__33360;
    wire N__33351;
    wire N__33348;
    wire N__33345;
    wire N__33340;
    wire N__33333;
    wire N__33330;
    wire N__33321;
    wire N__33314;
    wire N__33301;
    wire N__33300;
    wire N__33299;
    wire N__33298;
    wire N__33297;
    wire N__33296;
    wire N__33295;
    wire N__33294;
    wire N__33291;
    wire N__33290;
    wire N__33289;
    wire N__33288;
    wire N__33287;
    wire N__33286;
    wire N__33285;
    wire N__33284;
    wire N__33283;
    wire N__33282;
    wire N__33281;
    wire N__33270;
    wire N__33269;
    wire N__33268;
    wire N__33267;
    wire N__33266;
    wire N__33265;
    wire N__33264;
    wire N__33261;
    wire N__33248;
    wire N__33237;
    wire N__33236;
    wire N__33235;
    wire N__33234;
    wire N__33233;
    wire N__33232;
    wire N__33231;
    wire N__33230;
    wire N__33227;
    wire N__33224;
    wire N__33211;
    wire N__33204;
    wire N__33203;
    wire N__33202;
    wire N__33201;
    wire N__33192;
    wire N__33189;
    wire N__33188;
    wire N__33185;
    wire N__33184;
    wire N__33183;
    wire N__33180;
    wire N__33177;
    wire N__33170;
    wire N__33163;
    wire N__33158;
    wire N__33149;
    wire N__33136;
    wire N__33135;
    wire N__33134;
    wire N__33133;
    wire N__33128;
    wire N__33123;
    wire N__33122;
    wire N__33117;
    wire N__33116;
    wire N__33115;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33089;
    wire N__33088;
    wire N__33085;
    wire N__33080;
    wire N__33077;
    wire N__33070;
    wire N__33067;
    wire N__33064;
    wire N__33061;
    wire N__33060;
    wire N__33059;
    wire N__33058;
    wire N__33055;
    wire N__33052;
    wire N__33049;
    wire N__33046;
    wire N__33045;
    wire N__33044;
    wire N__33043;
    wire N__33042;
    wire N__33041;
    wire N__33040;
    wire N__33039;
    wire N__33038;
    wire N__33037;
    wire N__33032;
    wire N__33027;
    wire N__33024;
    wire N__33023;
    wire N__33022;
    wire N__33019;
    wire N__33018;
    wire N__33017;
    wire N__33016;
    wire N__33015;
    wire N__33012;
    wire N__33009;
    wire N__33006;
    wire N__33003;
    wire N__33000;
    wire N__32999;
    wire N__32996;
    wire N__32995;
    wire N__32994;
    wire N__32991;
    wire N__32990;
    wire N__32983;
    wire N__32980;
    wire N__32979;
    wire N__32978;
    wire N__32975;
    wire N__32974;
    wire N__32973;
    wire N__32972;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32964;
    wire N__32963;
    wire N__32962;
    wire N__32961;
    wire N__32958;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32948;
    wire N__32943;
    wire N__32942;
    wire N__32941;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32910;
    wire N__32907;
    wire N__32904;
    wire N__32903;
    wire N__32902;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32889;
    wire N__32886;
    wire N__32885;
    wire N__32884;
    wire N__32879;
    wire N__32876;
    wire N__32875;
    wire N__32874;
    wire N__32871;
    wire N__32870;
    wire N__32867;
    wire N__32864;
    wire N__32861;
    wire N__32858;
    wire N__32857;
    wire N__32852;
    wire N__32847;
    wire N__32844;
    wire N__32843;
    wire N__32840;
    wire N__32839;
    wire N__32832;
    wire N__32829;
    wire N__32822;
    wire N__32819;
    wire N__32818;
    wire N__32817;
    wire N__32812;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32800;
    wire N__32797;
    wire N__32794;
    wire N__32789;
    wire N__32786;
    wire N__32781;
    wire N__32778;
    wire N__32775;
    wire N__32770;
    wire N__32767;
    wire N__32766;
    wire N__32763;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32755;
    wire N__32754;
    wire N__32753;
    wire N__32752;
    wire N__32751;
    wire N__32748;
    wire N__32747;
    wire N__32744;
    wire N__32739;
    wire N__32736;
    wire N__32735;
    wire N__32732;
    wire N__32727;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32716;
    wire N__32715;
    wire N__32714;
    wire N__32709;
    wire N__32704;
    wire N__32701;
    wire N__32698;
    wire N__32689;
    wire N__32686;
    wire N__32681;
    wire N__32672;
    wire N__32669;
    wire N__32664;
    wire N__32661;
    wire N__32660;
    wire N__32659;
    wire N__32656;
    wire N__32653;
    wire N__32652;
    wire N__32651;
    wire N__32650;
    wire N__32647;
    wire N__32644;
    wire N__32641;
    wire N__32638;
    wire N__32637;
    wire N__32634;
    wire N__32631;
    wire N__32630;
    wire N__32629;
    wire N__32626;
    wire N__32623;
    wire N__32620;
    wire N__32617;
    wire N__32612;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32600;
    wire N__32597;
    wire N__32592;
    wire N__32589;
    wire N__32586;
    wire N__32583;
    wire N__32576;
    wire N__32573;
    wire N__32568;
    wire N__32565;
    wire N__32556;
    wire N__32553;
    wire N__32550;
    wire N__32549;
    wire N__32546;
    wire N__32543;
    wire N__32540;
    wire N__32537;
    wire N__32536;
    wire N__32535;
    wire N__32532;
    wire N__32523;
    wire N__32520;
    wire N__32515;
    wire N__32512;
    wire N__32509;
    wire N__32508;
    wire N__32507;
    wire N__32504;
    wire N__32499;
    wire N__32494;
    wire N__32491;
    wire N__32488;
    wire N__32483;
    wire N__32476;
    wire N__32471;
    wire N__32464;
    wire N__32455;
    wire N__32452;
    wire N__32445;
    wire N__32442;
    wire N__32439;
    wire N__32436;
    wire N__32429;
    wire N__32422;
    wire N__32419;
    wire N__32418;
    wire N__32415;
    wire N__32410;
    wire N__32405;
    wire N__32400;
    wire N__32395;
    wire N__32388;
    wire N__32379;
    wire N__32372;
    wire N__32369;
    wire N__32368;
    wire N__32367;
    wire N__32364;
    wire N__32359;
    wire N__32352;
    wire N__32349;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32323;
    wire N__32320;
    wire N__32319;
    wire N__32318;
    wire N__32317;
    wire N__32316;
    wire N__32315;
    wire N__32314;
    wire N__32311;
    wire N__32308;
    wire N__32305;
    wire N__32302;
    wire N__32299;
    wire N__32296;
    wire N__32293;
    wire N__32292;
    wire N__32291;
    wire N__32290;
    wire N__32289;
    wire N__32288;
    wire N__32287;
    wire N__32286;
    wire N__32285;
    wire N__32284;
    wire N__32281;
    wire N__32278;
    wire N__32275;
    wire N__32272;
    wire N__32269;
    wire N__32266;
    wire N__32263;
    wire N__32230;
    wire N__32227;
    wire N__32224;
    wire N__32223;
    wire N__32218;
    wire N__32215;
    wire N__32212;
    wire N__32209;
    wire N__32206;
    wire N__32203;
    wire N__32200;
    wire N__32197;
    wire N__32194;
    wire N__32191;
    wire N__32190;
    wire N__32187;
    wire N__32184;
    wire N__32181;
    wire N__32176;
    wire N__32173;
    wire N__32170;
    wire N__32169;
    wire N__32168;
    wire N__32165;
    wire N__32162;
    wire N__32159;
    wire N__32158;
    wire N__32155;
    wire N__32152;
    wire N__32147;
    wire N__32144;
    wire N__32137;
    wire N__32134;
    wire N__32131;
    wire N__32128;
    wire N__32125;
    wire N__32122;
    wire N__32119;
    wire N__32118;
    wire N__32113;
    wire N__32110;
    wire N__32109;
    wire N__32104;
    wire N__32101;
    wire N__32098;
    wire N__32095;
    wire N__32092;
    wire N__32089;
    wire N__32086;
    wire N__32083;
    wire N__32082;
    wire N__32081;
    wire N__32080;
    wire N__32079;
    wire N__32078;
    wire N__32077;
    wire N__32076;
    wire N__32075;
    wire N__32074;
    wire N__32073;
    wire N__32070;
    wire N__32065;
    wire N__32060;
    wire N__32059;
    wire N__32054;
    wire N__32051;
    wire N__32050;
    wire N__32045;
    wire N__32042;
    wire N__32035;
    wire N__32034;
    wire N__32033;
    wire N__32032;
    wire N__32029;
    wire N__32026;
    wire N__32021;
    wire N__32020;
    wire N__32017;
    wire N__32016;
    wire N__32011;
    wire N__32010;
    wire N__32009;
    wire N__32008;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31989;
    wire N__31988;
    wire N__31987;
    wire N__31986;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31971;
    wire N__31968;
    wire N__31965;
    wire N__31956;
    wire N__31951;
    wire N__31948;
    wire N__31945;
    wire N__31934;
    wire N__31925;
    wire N__31920;
    wire N__31917;
    wire N__31912;
    wire N__31909;
    wire N__31908;
    wire N__31905;
    wire N__31902;
    wire N__31897;
    wire N__31896;
    wire N__31895;
    wire N__31894;
    wire N__31893;
    wire N__31892;
    wire N__31891;
    wire N__31888;
    wire N__31885;
    wire N__31884;
    wire N__31883;
    wire N__31880;
    wire N__31879;
    wire N__31876;
    wire N__31875;
    wire N__31872;
    wire N__31869;
    wire N__31866;
    wire N__31861;
    wire N__31860;
    wire N__31857;
    wire N__31852;
    wire N__31851;
    wire N__31848;
    wire N__31845;
    wire N__31840;
    wire N__31833;
    wire N__31830;
    wire N__31827;
    wire N__31824;
    wire N__31821;
    wire N__31818;
    wire N__31809;
    wire N__31806;
    wire N__31795;
    wire N__31792;
    wire N__31791;
    wire N__31790;
    wire N__31789;
    wire N__31788;
    wire N__31787;
    wire N__31786;
    wire N__31783;
    wire N__31780;
    wire N__31777;
    wire N__31776;
    wire N__31775;
    wire N__31768;
    wire N__31765;
    wire N__31764;
    wire N__31757;
    wire N__31754;
    wire N__31753;
    wire N__31750;
    wire N__31749;
    wire N__31748;
    wire N__31745;
    wire N__31742;
    wire N__31739;
    wire N__31736;
    wire N__31733;
    wire N__31730;
    wire N__31727;
    wire N__31724;
    wire N__31721;
    wire N__31720;
    wire N__31717;
    wire N__31712;
    wire N__31703;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31687;
    wire N__31682;
    wire N__31679;
    wire N__31674;
    wire N__31669;
    wire N__31666;
    wire N__31663;
    wire N__31660;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31638;
    wire N__31635;
    wire N__31632;
    wire N__31629;
    wire N__31626;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31599;
    wire N__31596;
    wire N__31593;
    wire N__31588;
    wire N__31585;
    wire N__31582;
    wire N__31579;
    wire N__31576;
    wire N__31573;
    wire N__31570;
    wire N__31567;
    wire N__31564;
    wire N__31561;
    wire N__31560;
    wire N__31555;
    wire N__31552;
    wire N__31549;
    wire N__31548;
    wire N__31547;
    wire N__31544;
    wire N__31541;
    wire N__31538;
    wire N__31537;
    wire N__31534;
    wire N__31533;
    wire N__31528;
    wire N__31525;
    wire N__31524;
    wire N__31523;
    wire N__31522;
    wire N__31521;
    wire N__31520;
    wire N__31517;
    wire N__31514;
    wire N__31509;
    wire N__31506;
    wire N__31501;
    wire N__31498;
    wire N__31495;
    wire N__31480;
    wire N__31479;
    wire N__31478;
    wire N__31475;
    wire N__31472;
    wire N__31471;
    wire N__31470;
    wire N__31465;
    wire N__31464;
    wire N__31461;
    wire N__31460;
    wire N__31459;
    wire N__31456;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31443;
    wire N__31440;
    wire N__31437;
    wire N__31434;
    wire N__31431;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31405;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31393;
    wire N__31390;
    wire N__31387;
    wire N__31384;
    wire N__31381;
    wire N__31378;
    wire N__31377;
    wire N__31376;
    wire N__31375;
    wire N__31374;
    wire N__31373;
    wire N__31370;
    wire N__31369;
    wire N__31366;
    wire N__31365;
    wire N__31364;
    wire N__31361;
    wire N__31360;
    wire N__31359;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31351;
    wire N__31350;
    wire N__31349;
    wire N__31348;
    wire N__31347;
    wire N__31346;
    wire N__31345;
    wire N__31344;
    wire N__31343;
    wire N__31342;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31327;
    wire N__31324;
    wire N__31323;
    wire N__31322;
    wire N__31321;
    wire N__31320;
    wire N__31311;
    wire N__31302;
    wire N__31299;
    wire N__31296;
    wire N__31291;
    wire N__31290;
    wire N__31289;
    wire N__31288;
    wire N__31287;
    wire N__31284;
    wire N__31283;
    wire N__31278;
    wire N__31273;
    wire N__31264;
    wire N__31261;
    wire N__31256;
    wire N__31251;
    wire N__31246;
    wire N__31239;
    wire N__31234;
    wire N__31231;
    wire N__31224;
    wire N__31221;
    wire N__31214;
    wire N__31207;
    wire N__31204;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31182;
    wire N__31181;
    wire N__31180;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31168;
    wire N__31165;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31149;
    wire N__31148;
    wire N__31145;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31120;
    wire N__31117;
    wire N__31116;
    wire N__31115;
    wire N__31114;
    wire N__31111;
    wire N__31110;
    wire N__31109;
    wire N__31108;
    wire N__31105;
    wire N__31104;
    wire N__31103;
    wire N__31102;
    wire N__31099;
    wire N__31098;
    wire N__31097;
    wire N__31096;
    wire N__31095;
    wire N__31094;
    wire N__31089;
    wire N__31088;
    wire N__31087;
    wire N__31086;
    wire N__31083;
    wire N__31082;
    wire N__31081;
    wire N__31080;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31072;
    wire N__31069;
    wire N__31066;
    wire N__31065;
    wire N__31062;
    wire N__31061;
    wire N__31056;
    wire N__31053;
    wire N__31052;
    wire N__31051;
    wire N__31050;
    wire N__31049;
    wire N__31040;
    wire N__31037;
    wire N__31030;
    wire N__31027;
    wire N__31024;
    wire N__31021;
    wire N__31018;
    wire N__31017;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31003;
    wire N__31002;
    wire N__31001;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30983;
    wire N__30974;
    wire N__30967;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30937;
    wire N__30932;
    wire N__30929;
    wire N__30926;
    wire N__30923;
    wire N__30920;
    wire N__30915;
    wire N__30904;
    wire N__30895;
    wire N__30880;
    wire N__30879;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30871;
    wire N__30870;
    wire N__30869;
    wire N__30866;
    wire N__30865;
    wire N__30862;
    wire N__30861;
    wire N__30856;
    wire N__30853;
    wire N__30852;
    wire N__30849;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30833;
    wire N__30830;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30818;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30796;
    wire N__30793;
    wire N__30790;
    wire N__30787;
    wire N__30784;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30771;
    wire N__30770;
    wire N__30769;
    wire N__30768;
    wire N__30765;
    wire N__30764;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30749;
    wire N__30748;
    wire N__30745;
    wire N__30742;
    wire N__30739;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30725;
    wire N__30720;
    wire N__30717;
    wire N__30712;
    wire N__30707;
    wire N__30700;
    wire N__30699;
    wire N__30698;
    wire N__30695;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30684;
    wire N__30683;
    wire N__30680;
    wire N__30679;
    wire N__30678;
    wire N__30677;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30667;
    wire N__30662;
    wire N__30659;
    wire N__30654;
    wire N__30649;
    wire N__30646;
    wire N__30643;
    wire N__30638;
    wire N__30631;
    wire N__30628;
    wire N__30625;
    wire N__30620;
    wire N__30613;
    wire N__30612;
    wire N__30607;
    wire N__30604;
    wire N__30601;
    wire N__30600;
    wire N__30597;
    wire N__30596;
    wire N__30593;
    wire N__30590;
    wire N__30585;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30571;
    wire N__30570;
    wire N__30569;
    wire N__30568;
    wire N__30565;
    wire N__30560;
    wire N__30557;
    wire N__30556;
    wire N__30555;
    wire N__30552;
    wire N__30551;
    wire N__30550;
    wire N__30549;
    wire N__30548;
    wire N__30547;
    wire N__30546;
    wire N__30541;
    wire N__30538;
    wire N__30535;
    wire N__30534;
    wire N__30533;
    wire N__30532;
    wire N__30529;
    wire N__30528;
    wire N__30527;
    wire N__30524;
    wire N__30523;
    wire N__30522;
    wire N__30515;
    wire N__30510;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30494;
    wire N__30491;
    wire N__30488;
    wire N__30485;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30475;
    wire N__30470;
    wire N__30469;
    wire N__30466;
    wire N__30459;
    wire N__30452;
    wire N__30451;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30430;
    wire N__30427;
    wire N__30424;
    wire N__30419;
    wire N__30414;
    wire N__30411;
    wire N__30408;
    wire N__30405;
    wire N__30400;
    wire N__30391;
    wire N__30388;
    wire N__30387;
    wire N__30386;
    wire N__30385;
    wire N__30384;
    wire N__30383;
    wire N__30382;
    wire N__30381;
    wire N__30380;
    wire N__30377;
    wire N__30376;
    wire N__30375;
    wire N__30374;
    wire N__30373;
    wire N__30372;
    wire N__30371;
    wire N__30368;
    wire N__30367;
    wire N__30366;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30358;
    wire N__30355;
    wire N__30354;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30338;
    wire N__30333;
    wire N__30328;
    wire N__30325;
    wire N__30316;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30295;
    wire N__30292;
    wire N__30289;
    wire N__30284;
    wire N__30277;
    wire N__30276;
    wire N__30275;
    wire N__30274;
    wire N__30269;
    wire N__30262;
    wire N__30259;
    wire N__30250;
    wire N__30245;
    wire N__30244;
    wire N__30243;
    wire N__30240;
    wire N__30233;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30219;
    wire N__30218;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30206;
    wire N__30203;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30185;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30159;
    wire N__30158;
    wire N__30157;
    wire N__30154;
    wire N__30153;
    wire N__30150;
    wire N__30149;
    wire N__30148;
    wire N__30147;
    wire N__30146;
    wire N__30145;
    wire N__30144;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30123;
    wire N__30120;
    wire N__30119;
    wire N__30118;
    wire N__30117;
    wire N__30116;
    wire N__30115;
    wire N__30114;
    wire N__30113;
    wire N__30110;
    wire N__30109;
    wire N__30108;
    wire N__30105;
    wire N__30104;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30082;
    wire N__30077;
    wire N__30074;
    wire N__30069;
    wire N__30062;
    wire N__30057;
    wire N__30050;
    wire N__30045;
    wire N__30038;
    wire N__30019;
    wire N__30018;
    wire N__30017;
    wire N__30014;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30006;
    wire N__30005;
    wire N__30004;
    wire N__30003;
    wire N__30000;
    wire N__29999;
    wire N__29998;
    wire N__29997;
    wire N__29994;
    wire N__29993;
    wire N__29990;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29971;
    wire N__29968;
    wire N__29967;
    wire N__29966;
    wire N__29965;
    wire N__29958;
    wire N__29955;
    wire N__29954;
    wire N__29949;
    wire N__29946;
    wire N__29943;
    wire N__29940;
    wire N__29937;
    wire N__29934;
    wire N__29931;
    wire N__29928;
    wire N__29921;
    wire N__29918;
    wire N__29913;
    wire N__29908;
    wire N__29887;
    wire N__29886;
    wire N__29885;
    wire N__29884;
    wire N__29883;
    wire N__29882;
    wire N__29881;
    wire N__29880;
    wire N__29879;
    wire N__29876;
    wire N__29873;
    wire N__29872;
    wire N__29871;
    wire N__29870;
    wire N__29869;
    wire N__29868;
    wire N__29865;
    wire N__29864;
    wire N__29863;
    wire N__29860;
    wire N__29857;
    wire N__29856;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29831;
    wire N__29830;
    wire N__29829;
    wire N__29828;
    wire N__29827;
    wire N__29826;
    wire N__29825;
    wire N__29824;
    wire N__29823;
    wire N__29822;
    wire N__29819;
    wire N__29816;
    wire N__29815;
    wire N__29812;
    wire N__29809;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29792;
    wire N__29789;
    wire N__29782;
    wire N__29775;
    wire N__29772;
    wire N__29767;
    wire N__29760;
    wire N__29753;
    wire N__29752;
    wire N__29749;
    wire N__29748;
    wire N__29745;
    wire N__29740;
    wire N__29737;
    wire N__29734;
    wire N__29731;
    wire N__29728;
    wire N__29723;
    wire N__29712;
    wire N__29705;
    wire N__29700;
    wire N__29683;
    wire N__29682;
    wire N__29681;
    wire N__29678;
    wire N__29677;
    wire N__29676;
    wire N__29675;
    wire N__29674;
    wire N__29673;
    wire N__29672;
    wire N__29671;
    wire N__29668;
    wire N__29667;
    wire N__29662;
    wire N__29661;
    wire N__29660;
    wire N__29659;
    wire N__29652;
    wire N__29649;
    wire N__29648;
    wire N__29647;
    wire N__29640;
    wire N__29639;
    wire N__29636;
    wire N__29635;
    wire N__29632;
    wire N__29631;
    wire N__29628;
    wire N__29623;
    wire N__29620;
    wire N__29617;
    wire N__29616;
    wire N__29615;
    wire N__29614;
    wire N__29613;
    wire N__29612;
    wire N__29611;
    wire N__29610;
    wire N__29609;
    wire N__29608;
    wire N__29607;
    wire N__29606;
    wire N__29605;
    wire N__29604;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29583;
    wire N__29580;
    wire N__29571;
    wire N__29568;
    wire N__29561;
    wire N__29552;
    wire N__29545;
    wire N__29540;
    wire N__29537;
    wire N__29530;
    wire N__29509;
    wire N__29508;
    wire N__29503;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29490;
    wire N__29485;
    wire N__29484;
    wire N__29483;
    wire N__29480;
    wire N__29479;
    wire N__29478;
    wire N__29477;
    wire N__29476;
    wire N__29475;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29465;
    wire N__29460;
    wire N__29457;
    wire N__29454;
    wire N__29453;
    wire N__29450;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29438;
    wire N__29437;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29420;
    wire N__29415;
    wire N__29410;
    wire N__29405;
    wire N__29402;
    wire N__29389;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29381;
    wire N__29378;
    wire N__29377;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29360;
    wire N__29357;
    wire N__29354;
    wire N__29347;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29327;
    wire N__29324;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29308;
    wire N__29307;
    wire N__29306;
    wire N__29305;
    wire N__29304;
    wire N__29299;
    wire N__29298;
    wire N__29297;
    wire N__29296;
    wire N__29295;
    wire N__29294;
    wire N__29293;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29274;
    wire N__29273;
    wire N__29270;
    wire N__29267;
    wire N__29262;
    wire N__29261;
    wire N__29258;
    wire N__29257;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29249;
    wire N__29246;
    wire N__29245;
    wire N__29242;
    wire N__29239;
    wire N__29236;
    wire N__29233;
    wire N__29228;
    wire N__29225;
    wire N__29224;
    wire N__29221;
    wire N__29218;
    wire N__29215;
    wire N__29212;
    wire N__29207;
    wire N__29200;
    wire N__29195;
    wire N__29192;
    wire N__29187;
    wire N__29184;
    wire N__29179;
    wire N__29158;
    wire N__29157;
    wire N__29156;
    wire N__29155;
    wire N__29154;
    wire N__29153;
    wire N__29152;
    wire N__29151;
    wire N__29146;
    wire N__29145;
    wire N__29142;
    wire N__29141;
    wire N__29140;
    wire N__29139;
    wire N__29138;
    wire N__29137;
    wire N__29136;
    wire N__29133;
    wire N__29132;
    wire N__29131;
    wire N__29130;
    wire N__29129;
    wire N__29128;
    wire N__29127;
    wire N__29124;
    wire N__29123;
    wire N__29122;
    wire N__29119;
    wire N__29114;
    wire N__29111;
    wire N__29104;
    wire N__29103;
    wire N__29102;
    wire N__29093;
    wire N__29090;
    wire N__29087;
    wire N__29080;
    wire N__29079;
    wire N__29076;
    wire N__29075;
    wire N__29074;
    wire N__29071;
    wire N__29060;
    wire N__29055;
    wire N__29052;
    wire N__29049;
    wire N__29046;
    wire N__29043;
    wire N__29038;
    wire N__29035;
    wire N__29032;
    wire N__29031;
    wire N__29028;
    wire N__29027;
    wire N__29022;
    wire N__29017;
    wire N__29012;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28966;
    wire N__28965;
    wire N__28964;
    wire N__28963;
    wire N__28962;
    wire N__28959;
    wire N__28954;
    wire N__28953;
    wire N__28952;
    wire N__28951;
    wire N__28950;
    wire N__28945;
    wire N__28944;
    wire N__28943;
    wire N__28938;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28923;
    wire N__28922;
    wire N__28919;
    wire N__28916;
    wire N__28913;
    wire N__28910;
    wire N__28909;
    wire N__28902;
    wire N__28895;
    wire N__28892;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28876;
    wire N__28873;
    wire N__28864;
    wire N__28863;
    wire N__28862;
    wire N__28861;
    wire N__28860;
    wire N__28859;
    wire N__28858;
    wire N__28857;
    wire N__28856;
    wire N__28855;
    wire N__28852;
    wire N__28851;
    wire N__28850;
    wire N__28845;
    wire N__28844;
    wire N__28843;
    wire N__28838;
    wire N__28835;
    wire N__28834;
    wire N__28831;
    wire N__28830;
    wire N__28829;
    wire N__28826;
    wire N__28821;
    wire N__28820;
    wire N__28819;
    wire N__28818;
    wire N__28817;
    wire N__28816;
    wire N__28815;
    wire N__28808;
    wire N__28805;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28791;
    wire N__28788;
    wire N__28785;
    wire N__28784;
    wire N__28781;
    wire N__28780;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28762;
    wire N__28761;
    wire N__28760;
    wire N__28759;
    wire N__28758;
    wire N__28757;
    wire N__28756;
    wire N__28753;
    wire N__28746;
    wire N__28743;
    wire N__28738;
    wire N__28735;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28723;
    wire N__28720;
    wire N__28713;
    wire N__28706;
    wire N__28699;
    wire N__28694;
    wire N__28669;
    wire N__28668;
    wire N__28665;
    wire N__28660;
    wire N__28657;
    wire N__28654;
    wire N__28653;
    wire N__28650;
    wire N__28647;
    wire N__28644;
    wire N__28643;
    wire N__28642;
    wire N__28641;
    wire N__28640;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28615;
    wire N__28600;
    wire N__28599;
    wire N__28598;
    wire N__28597;
    wire N__28594;
    wire N__28591;
    wire N__28590;
    wire N__28589;
    wire N__28588;
    wire N__28587;
    wire N__28586;
    wire N__28583;
    wire N__28580;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28566;
    wire N__28565;
    wire N__28564;
    wire N__28563;
    wire N__28560;
    wire N__28559;
    wire N__28556;
    wire N__28555;
    wire N__28554;
    wire N__28553;
    wire N__28546;
    wire N__28539;
    wire N__28534;
    wire N__28529;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28512;
    wire N__28505;
    wire N__28502;
    wire N__28489;
    wire N__28486;
    wire N__28485;
    wire N__28484;
    wire N__28483;
    wire N__28482;
    wire N__28481;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28469;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28461;
    wire N__28458;
    wire N__28457;
    wire N__28454;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28436;
    wire N__28435;
    wire N__28432;
    wire N__28429;
    wire N__28424;
    wire N__28421;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28405;
    wire N__28400;
    wire N__28395;
    wire N__28384;
    wire N__28383;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28366;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28356;
    wire N__28355;
    wire N__28352;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28330;
    wire N__28329;
    wire N__28328;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28312;
    wire N__28303;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28279;
    wire N__28276;
    wire N__28273;
    wire N__28270;
    wire N__28269;
    wire N__28268;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28245;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28230;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28216;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28205;
    wire N__28202;
    wire N__28199;
    wire N__28198;
    wire N__28195;
    wire N__28190;
    wire N__28187;
    wire N__28180;
    wire N__28177;
    wire N__28176;
    wire N__28175;
    wire N__28174;
    wire N__28171;
    wire N__28170;
    wire N__28169;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28159;
    wire N__28156;
    wire N__28155;
    wire N__28152;
    wire N__28151;
    wire N__28150;
    wire N__28149;
    wire N__28148;
    wire N__28147;
    wire N__28144;
    wire N__28143;
    wire N__28142;
    wire N__28141;
    wire N__28140;
    wire N__28137;
    wire N__28130;
    wire N__28127;
    wire N__28118;
    wire N__28115;
    wire N__28112;
    wire N__28111;
    wire N__28108;
    wire N__28107;
    wire N__28106;
    wire N__28105;
    wire N__28100;
    wire N__28097;
    wire N__28092;
    wire N__28091;
    wire N__28088;
    wire N__28085;
    wire N__28080;
    wire N__28077;
    wire N__28072;
    wire N__28069;
    wire N__28068;
    wire N__28067;
    wire N__28064;
    wire N__28061;
    wire N__28058;
    wire N__28055;
    wire N__28052;
    wire N__28049;
    wire N__28046;
    wire N__28043;
    wire N__28040;
    wire N__28039;
    wire N__28036;
    wire N__28031;
    wire N__28030;
    wire N__28029;
    wire N__28028;
    wire N__28027;
    wire N__28026;
    wire N__28025;
    wire N__28022;
    wire N__28017;
    wire N__28012;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__27997;
    wire N__27992;
    wire N__27989;
    wire N__27984;
    wire N__27981;
    wire N__27976;
    wire N__27969;
    wire N__27962;
    wire N__27959;
    wire N__27934;
    wire N__27933;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27915;
    wire N__27914;
    wire N__27913;
    wire N__27912;
    wire N__27909;
    wire N__27906;
    wire N__27905;
    wire N__27902;
    wire N__27897;
    wire N__27892;
    wire N__27889;
    wire N__27880;
    wire N__27877;
    wire N__27874;
    wire N__27871;
    wire N__27870;
    wire N__27869;
    wire N__27866;
    wire N__27863;
    wire N__27860;
    wire N__27857;
    wire N__27852;
    wire N__27847;
    wire N__27844;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27826;
    wire N__27825;
    wire N__27824;
    wire N__27819;
    wire N__27816;
    wire N__27811;
    wire N__27810;
    wire N__27807;
    wire N__27804;
    wire N__27799;
    wire N__27796;
    wire N__27795;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27769;
    wire N__27766;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27739;
    wire N__27736;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27712;
    wire N__27711;
    wire N__27708;
    wire N__27705;
    wire N__27702;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27682;
    wire N__27679;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27667;
    wire N__27664;
    wire N__27661;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27649;
    wire N__27646;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27631;
    wire N__27628;
    wire N__27627;
    wire N__27624;
    wire N__27621;
    wire N__27618;
    wire N__27613;
    wire N__27610;
    wire N__27609;
    wire N__27606;
    wire N__27603;
    wire N__27600;
    wire N__27595;
    wire N__27592;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27577;
    wire N__27574;
    wire N__27573;
    wire N__27572;
    wire N__27571;
    wire N__27570;
    wire N__27569;
    wire N__27568;
    wire N__27567;
    wire N__27566;
    wire N__27565;
    wire N__27564;
    wire N__27563;
    wire N__27562;
    wire N__27561;
    wire N__27560;
    wire N__27559;
    wire N__27558;
    wire N__27557;
    wire N__27556;
    wire N__27555;
    wire N__27554;
    wire N__27553;
    wire N__27552;
    wire N__27551;
    wire N__27550;
    wire N__27549;
    wire N__27548;
    wire N__27547;
    wire N__27546;
    wire N__27545;
    wire N__27544;
    wire N__27543;
    wire N__27542;
    wire N__27541;
    wire N__27540;
    wire N__27539;
    wire N__27538;
    wire N__27537;
    wire N__27536;
    wire N__27535;
    wire N__27534;
    wire N__27533;
    wire N__27532;
    wire N__27531;
    wire N__27530;
    wire N__27529;
    wire N__27528;
    wire N__27527;
    wire N__27526;
    wire N__27525;
    wire N__27524;
    wire N__27523;
    wire N__27522;
    wire N__27513;
    wire N__27504;
    wire N__27495;
    wire N__27486;
    wire N__27479;
    wire N__27470;
    wire N__27461;
    wire N__27454;
    wire N__27445;
    wire N__27436;
    wire N__27427;
    wire N__27420;
    wire N__27415;
    wire N__27410;
    wire N__27407;
    wire N__27402;
    wire N__27399;
    wire N__27398;
    wire N__27395;
    wire N__27394;
    wire N__27391;
    wire N__27390;
    wire N__27389;
    wire N__27388;
    wire N__27387;
    wire N__27386;
    wire N__27385;
    wire N__27382;
    wire N__27381;
    wire N__27380;
    wire N__27377;
    wire N__27374;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27344;
    wire N__27341;
    wire N__27338;
    wire N__27283;
    wire N__27280;
    wire N__27277;
    wire N__27276;
    wire N__27273;
    wire N__27270;
    wire N__27267;
    wire N__27262;
    wire N__27259;
    wire N__27256;
    wire N__27255;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27244;
    wire N__27241;
    wire N__27238;
    wire N__27237;
    wire N__27236;
    wire N__27235;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27223;
    wire N__27220;
    wire N__27217;
    wire N__27214;
    wire N__27211;
    wire N__27208;
    wire N__27205;
    wire N__27200;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27138;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27127;
    wire N__27124;
    wire N__27119;
    wire N__27116;
    wire N__27111;
    wire N__27108;
    wire N__27103;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27091;
    wire N__27088;
    wire N__27087;
    wire N__27084;
    wire N__27081;
    wire N__27076;
    wire N__27073;
    wire N__27070;
    wire N__27069;
    wire N__27066;
    wire N__27063;
    wire N__27060;
    wire N__27055;
    wire N__27052;
    wire N__27051;
    wire N__27048;
    wire N__27045;
    wire N__27040;
    wire N__27037;
    wire N__27036;
    wire N__27033;
    wire N__27030;
    wire N__27025;
    wire N__27022;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27010;
    wire N__27007;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26995;
    wire N__26992;
    wire N__26991;
    wire N__26988;
    wire N__26985;
    wire N__26982;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26940;
    wire N__26939;
    wire N__26936;
    wire N__26933;
    wire N__26930;
    wire N__26927;
    wire N__26926;
    wire N__26925;
    wire N__26924;
    wire N__26917;
    wire N__26914;
    wire N__26909;
    wire N__26904;
    wire N__26899;
    wire N__26896;
    wire N__26893;
    wire N__26890;
    wire N__26887;
    wire N__26884;
    wire N__26883;
    wire N__26878;
    wire N__26875;
    wire N__26872;
    wire N__26869;
    wire N__26866;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26832;
    wire N__26829;
    wire N__26826;
    wire N__26823;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26809;
    wire N__26808;
    wire N__26803;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26779;
    wire N__26776;
    wire N__26773;
    wire N__26770;
    wire N__26767;
    wire N__26764;
    wire N__26761;
    wire N__26758;
    wire N__26755;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26731;
    wire N__26730;
    wire N__26727;
    wire N__26726;
    wire N__26723;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26698;
    wire N__26695;
    wire N__26692;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26680;
    wire N__26679;
    wire N__26676;
    wire N__26673;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26652;
    wire N__26651;
    wire N__26650;
    wire N__26649;
    wire N__26648;
    wire N__26645;
    wire N__26642;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26634;
    wire N__26633;
    wire N__26632;
    wire N__26631;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26615;
    wire N__26612;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26581;
    wire N__26578;
    wire N__26573;
    wire N__26570;
    wire N__26567;
    wire N__26564;
    wire N__26561;
    wire N__26556;
    wire N__26553;
    wire N__26548;
    wire N__26541;
    wire N__26538;
    wire N__26535;
    wire N__26532;
    wire N__26527;
    wire N__26518;
    wire N__26515;
    wire N__26512;
    wire N__26511;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26499;
    wire N__26494;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26484;
    wire N__26479;
    wire N__26476;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26466;
    wire N__26463;
    wire N__26460;
    wire N__26457;
    wire N__26454;
    wire N__26449;
    wire N__26446;
    wire N__26443;
    wire N__26440;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26427;
    wire N__26426;
    wire N__26425;
    wire N__26422;
    wire N__26421;
    wire N__26420;
    wire N__26419;
    wire N__26416;
    wire N__26415;
    wire N__26414;
    wire N__26411;
    wire N__26406;
    wire N__26403;
    wire N__26400;
    wire N__26397;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26382;
    wire N__26379;
    wire N__26376;
    wire N__26373;
    wire N__26370;
    wire N__26363;
    wire N__26360;
    wire N__26355;
    wire N__26344;
    wire N__26343;
    wire N__26340;
    wire N__26337;
    wire N__26334;
    wire N__26331;
    wire N__26328;
    wire N__26325;
    wire N__26322;
    wire N__26317;
    wire N__26314;
    wire N__26311;
    wire N__26310;
    wire N__26307;
    wire N__26304;
    wire N__26299;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26289;
    wire N__26284;
    wire N__26281;
    wire N__26278;
    wire N__26277;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26241;
    wire N__26236;
    wire N__26233;
    wire N__26232;
    wire N__26229;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26209;
    wire N__26208;
    wire N__26203;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26182;
    wire N__26179;
    wire N__26176;
    wire N__26173;
    wire N__26172;
    wire N__26169;
    wire N__26166;
    wire N__26163;
    wire N__26160;
    wire N__26155;
    wire N__26152;
    wire N__26149;
    wire N__26148;
    wire N__26145;
    wire N__26142;
    wire N__26137;
    wire N__26134;
    wire N__26133;
    wire N__26130;
    wire N__26127;
    wire N__26124;
    wire N__26119;
    wire N__26116;
    wire N__26115;
    wire N__26114;
    wire N__26111;
    wire N__26110;
    wire N__26107;
    wire N__26102;
    wire N__26099;
    wire N__26098;
    wire N__26097;
    wire N__26094;
    wire N__26091;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26081;
    wire N__26076;
    wire N__26073;
    wire N__26068;
    wire N__26059;
    wire N__26056;
    wire N__26053;
    wire N__26050;
    wire N__26047;
    wire N__26044;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26020;
    wire N__26017;
    wire N__26016;
    wire N__26011;
    wire N__26008;
    wire N__26007;
    wire N__26004;
    wire N__26001;
    wire N__25998;
    wire N__25995;
    wire N__25992;
    wire N__25987;
    wire N__25984;
    wire N__25981;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25960;
    wire N__25957;
    wire N__25954;
    wire N__25951;
    wire N__25948;
    wire N__25945;
    wire N__25942;
    wire N__25939;
    wire N__25936;
    wire N__25933;
    wire N__25930;
    wire N__25927;
    wire N__25924;
    wire N__25921;
    wire N__25918;
    wire N__25917;
    wire N__25914;
    wire N__25913;
    wire N__25908;
    wire N__25905;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25889;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25873;
    wire N__25870;
    wire N__25867;
    wire N__25864;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25851;
    wire N__25848;
    wire N__25847;
    wire N__25844;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25810;
    wire N__25807;
    wire N__25804;
    wire N__25803;
    wire N__25800;
    wire N__25799;
    wire N__25796;
    wire N__25795;
    wire N__25792;
    wire N__25787;
    wire N__25784;
    wire N__25777;
    wire N__25774;
    wire N__25773;
    wire N__25770;
    wire N__25769;
    wire N__25766;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25738;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25725;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25710;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25684;
    wire N__25681;
    wire N__25678;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25660;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25623;
    wire N__25622;
    wire N__25619;
    wire N__25618;
    wire N__25615;
    wire N__25614;
    wire N__25609;
    wire N__25606;
    wire N__25603;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25585;
    wire N__25582;
    wire N__25581;
    wire N__25576;
    wire N__25573;
    wire N__25570;
    wire N__25567;
    wire N__25564;
    wire N__25561;
    wire N__25560;
    wire N__25555;
    wire N__25552;
    wire N__25549;
    wire N__25548;
    wire N__25543;
    wire N__25540;
    wire N__25537;
    wire N__25534;
    wire N__25531;
    wire N__25528;
    wire N__25527;
    wire N__25522;
    wire N__25519;
    wire N__25516;
    wire N__25515;
    wire N__25510;
    wire N__25507;
    wire N__25504;
    wire N__25501;
    wire N__25498;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25488;
    wire N__25483;
    wire N__25480;
    wire N__25479;
    wire N__25474;
    wire N__25471;
    wire N__25468;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25456;
    wire N__25455;
    wire N__25450;
    wire N__25447;
    wire N__25444;
    wire N__25443;
    wire N__25440;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25428;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25414;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25381;
    wire N__25380;
    wire N__25377;
    wire N__25372;
    wire N__25369;
    wire N__25366;
    wire N__25363;
    wire N__25360;
    wire N__25357;
    wire N__25354;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25336;
    wire N__25333;
    wire N__25330;
    wire N__25329;
    wire N__25324;
    wire N__25321;
    wire N__25318;
    wire N__25315;
    wire N__25312;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25300;
    wire N__25297;
    wire N__25294;
    wire N__25293;
    wire N__25290;
    wire N__25287;
    wire N__25282;
    wire N__25279;
    wire N__25276;
    wire N__25273;
    wire N__25270;
    wire N__25267;
    wire N__25264;
    wire N__25261;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25243;
    wire N__25240;
    wire N__25239;
    wire N__25238;
    wire N__25237;
    wire N__25236;
    wire N__25235;
    wire N__25224;
    wire N__25221;
    wire N__25216;
    wire N__25215;
    wire N__25214;
    wire N__25213;
    wire N__25212;
    wire N__25211;
    wire N__25210;
    wire N__25199;
    wire N__25194;
    wire N__25189;
    wire N__25186;
    wire N__25185;
    wire N__25184;
    wire N__25181;
    wire N__25180;
    wire N__25179;
    wire N__25178;
    wire N__25177;
    wire N__25172;
    wire N__25165;
    wire N__25160;
    wire N__25153;
    wire N__25150;
    wire N__25147;
    wire N__25146;
    wire N__25145;
    wire N__25144;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25136;
    wire N__25133;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25125;
    wire N__25124;
    wire N__25119;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25086;
    wire N__25083;
    wire N__25080;
    wire N__25073;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25050;
    wire N__25047;
    wire N__25042;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25032;
    wire N__25029;
    wire N__25026;
    wire N__25021;
    wire N__25020;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25008;
    wire N__25005;
    wire N__25004;
    wire N__25001;
    wire N__25000;
    wire N__24999;
    wire N__24996;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24976;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24966;
    wire N__24963;
    wire N__24958;
    wire N__24955;
    wire N__24954;
    wire N__24953;
    wire N__24946;
    wire N__24943;
    wire N__24936;
    wire N__24935;
    wire N__24934;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24914;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24883;
    wire N__24880;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24843;
    wire N__24838;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24820;
    wire N__24817;
    wire N__24814;
    wire N__24813;
    wire N__24812;
    wire N__24809;
    wire N__24808;
    wire N__24807;
    wire N__24802;
    wire N__24799;
    wire N__24798;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24766;
    wire N__24757;
    wire N__24754;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24742;
    wire N__24741;
    wire N__24740;
    wire N__24739;
    wire N__24736;
    wire N__24733;
    wire N__24728;
    wire N__24725;
    wire N__24724;
    wire N__24723;
    wire N__24718;
    wire N__24715;
    wire N__24710;
    wire N__24707;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24684;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24658;
    wire N__24655;
    wire N__24654;
    wire N__24653;
    wire N__24648;
    wire N__24645;
    wire N__24642;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24627;
    wire N__24626;
    wire N__24623;
    wire N__24618;
    wire N__24615;
    wire N__24610;
    wire N__24609;
    wire N__24604;
    wire N__24601;
    wire N__24598;
    wire N__24595;
    wire N__24592;
    wire N__24589;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24559;
    wire N__24556;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24534;
    wire N__24529;
    wire N__24526;
    wire N__24525;
    wire N__24522;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24507;
    wire N__24506;
    wire N__24503;
    wire N__24502;
    wire N__24501;
    wire N__24500;
    wire N__24499;
    wire N__24496;
    wire N__24495;
    wire N__24494;
    wire N__24493;
    wire N__24492;
    wire N__24489;
    wire N__24476;
    wire N__24473;
    wire N__24472;
    wire N__24469;
    wire N__24468;
    wire N__24465;
    wire N__24464;
    wire N__24461;
    wire N__24456;
    wire N__24451;
    wire N__24440;
    wire N__24437;
    wire N__24432;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24420;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24375;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24325;
    wire N__24322;
    wire N__24319;
    wire N__24316;
    wire N__24315;
    wire N__24310;
    wire N__24307;
    wire N__24306;
    wire N__24301;
    wire N__24298;
    wire N__24295;
    wire N__24292;
    wire N__24289;
    wire N__24286;
    wire N__24285;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24241;
    wire N__24238;
    wire N__24235;
    wire N__24234;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24169;
    wire N__24166;
    wire N__24163;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24151;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24139;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24123;
    wire N__24118;
    wire N__24115;
    wire N__24112;
    wire N__24109;
    wire N__24108;
    wire N__24103;
    wire N__24100;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24085;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24064;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24046;
    wire N__24043;
    wire N__24040;
    wire N__24037;
    wire N__24034;
    wire N__24031;
    wire N__24028;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__24001;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23991;
    wire N__23990;
    wire N__23985;
    wire N__23982;
    wire N__23977;
    wire N__23974;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23949;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23922;
    wire N__23919;
    wire N__23918;
    wire N__23915;
    wire N__23908;
    wire N__23905;
    wire N__23904;
    wire N__23901;
    wire N__23898;
    wire N__23895;
    wire N__23892;
    wire N__23889;
    wire N__23884;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23872;
    wire N__23869;
    wire N__23866;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23854;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23841;
    wire N__23838;
    wire N__23837;
    wire N__23834;
    wire N__23833;
    wire N__23832;
    wire N__23829;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23809;
    wire N__23808;
    wire N__23805;
    wire N__23802;
    wire N__23797;
    wire N__23794;
    wire N__23791;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23767;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23743;
    wire N__23740;
    wire N__23737;
    wire N__23736;
    wire N__23733;
    wire N__23732;
    wire N__23729;
    wire N__23722;
    wire N__23719;
    wire N__23716;
    wire N__23713;
    wire N__23710;
    wire N__23707;
    wire N__23704;
    wire N__23703;
    wire N__23700;
    wire N__23699;
    wire N__23696;
    wire N__23695;
    wire N__23692;
    wire N__23687;
    wire N__23684;
    wire N__23677;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23665;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23653;
    wire N__23652;
    wire N__23649;
    wire N__23646;
    wire N__23643;
    wire N__23638;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23602;
    wire N__23601;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23569;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23512;
    wire N__23511;
    wire N__23508;
    wire N__23505;
    wire N__23500;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23488;
    wire N__23487;
    wire N__23484;
    wire N__23481;
    wire N__23478;
    wire N__23473;
    wire N__23472;
    wire N__23469;
    wire N__23466;
    wire N__23461;
    wire N__23460;
    wire N__23459;
    wire N__23458;
    wire N__23457;
    wire N__23456;
    wire N__23447;
    wire N__23442;
    wire N__23437;
    wire N__23434;
    wire N__23431;
    wire N__23430;
    wire N__23425;
    wire N__23422;
    wire N__23421;
    wire N__23420;
    wire N__23419;
    wire N__23418;
    wire N__23417;
    wire N__23412;
    wire N__23403;
    wire N__23398;
    wire N__23395;
    wire N__23392;
    wire N__23389;
    wire N__23386;
    wire N__23385;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23374;
    wire N__23371;
    wire N__23370;
    wire N__23369;
    wire N__23368;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23353;
    wire N__23348;
    wire N__23345;
    wire N__23340;
    wire N__23339;
    wire N__23338;
    wire N__23335;
    wire N__23332;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23308;
    wire N__23307;
    wire N__23306;
    wire N__23305;
    wire N__23304;
    wire N__23297;
    wire N__23292;
    wire N__23289;
    wire N__23284;
    wire N__23283;
    wire N__23280;
    wire N__23277;
    wire N__23272;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23260;
    wire N__23259;
    wire N__23256;
    wire N__23253;
    wire N__23250;
    wire N__23245;
    wire N__23244;
    wire N__23241;
    wire N__23238;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23218;
    wire N__23217;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23194;
    wire N__23193;
    wire N__23190;
    wire N__23187;
    wire N__23182;
    wire N__23181;
    wire N__23178;
    wire N__23175;
    wire N__23172;
    wire N__23167;
    wire N__23164;
    wire N__23163;
    wire N__23160;
    wire N__23157;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23104;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23058;
    wire N__23057;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23032;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23020;
    wire N__23019;
    wire N__23018;
    wire N__23017;
    wire N__23016;
    wire N__23015;
    wire N__23012;
    wire N__23005;
    wire N__23000;
    wire N__22993;
    wire N__22990;
    wire N__22989;
    wire N__22988;
    wire N__22987;
    wire N__22984;
    wire N__22983;
    wire N__22980;
    wire N__22977;
    wire N__22974;
    wire N__22969;
    wire N__22966;
    wire N__22961;
    wire N__22960;
    wire N__22957;
    wire N__22952;
    wire N__22949;
    wire N__22944;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22911;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22896;
    wire N__22895;
    wire N__22894;
    wire N__22893;
    wire N__22890;
    wire N__22889;
    wire N__22886;
    wire N__22885;
    wire N__22880;
    wire N__22875;
    wire N__22874;
    wire N__22871;
    wire N__22866;
    wire N__22863;
    wire N__22862;
    wire N__22861;
    wire N__22858;
    wire N__22857;
    wire N__22854;
    wire N__22849;
    wire N__22846;
    wire N__22841;
    wire N__22838;
    wire N__22833;
    wire N__22822;
    wire N__22819;
    wire N__22816;
    wire N__22813;
    wire N__22810;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22765;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22710;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22684;
    wire N__22681;
    wire N__22678;
    wire N__22675;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22663;
    wire N__22660;
    wire N__22657;
    wire N__22656;
    wire N__22651;
    wire N__22648;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22635;
    wire N__22632;
    wire N__22629;
    wire N__22624;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22558;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22497;
    wire N__22494;
    wire N__22493;
    wire N__22492;
    wire N__22491;
    wire N__22486;
    wire N__22483;
    wire N__22478;
    wire N__22471;
    wire N__22470;
    wire N__22469;
    wire N__22466;
    wire N__22465;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22451;
    wire N__22444;
    wire N__22443;
    wire N__22440;
    wire N__22439;
    wire N__22436;
    wire N__22429;
    wire N__22426;
    wire N__22425;
    wire N__22422;
    wire N__22421;
    wire N__22420;
    wire N__22417;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22383;
    wire N__22382;
    wire N__22381;
    wire N__22380;
    wire N__22377;
    wire N__22372;
    wire N__22367;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22353;
    wire N__22352;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22340;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22300;
    wire N__22299;
    wire N__22298;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22282;
    wire N__22281;
    wire N__22278;
    wire N__22277;
    wire N__22276;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22258;
    wire N__22255;
    wire N__22252;
    wire N__22251;
    wire N__22248;
    wire N__22247;
    wire N__22244;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22219;
    wire N__22218;
    wire N__22215;
    wire N__22214;
    wire N__22211;
    wire N__22204;
    wire N__22201;
    wire N__22200;
    wire N__22197;
    wire N__22194;
    wire N__22189;
    wire N__22186;
    wire N__22183;
    wire N__22180;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22090;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22072;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22053;
    wire N__22052;
    wire N__22049;
    wire N__22048;
    wire N__22045;
    wire N__22040;
    wire N__22037;
    wire N__22030;
    wire N__22027;
    wire N__22024;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21972;
    wire N__21969;
    wire N__21964;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21952;
    wire N__21949;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21901;
    wire N__21898;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21847;
    wire N__21844;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21832;
    wire N__21829;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21811;
    wire N__21808;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21790;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21775;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21757;
    wire N__21754;
    wire N__21753;
    wire N__21752;
    wire N__21751;
    wire N__21750;
    wire N__21749;
    wire N__21748;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21730;
    wire N__21727;
    wire N__21726;
    wire N__21725;
    wire N__21724;
    wire N__21723;
    wire N__21722;
    wire N__21719;
    wire N__21718;
    wire N__21713;
    wire N__21710;
    wire N__21705;
    wire N__21702;
    wire N__21697;
    wire N__21686;
    wire N__21681;
    wire N__21678;
    wire N__21667;
    wire N__21666;
    wire N__21663;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21603;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21582;
    wire N__21577;
    wire N__21574;
    wire N__21573;
    wire N__21570;
    wire N__21565;
    wire N__21562;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21547;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21436;
    wire N__21433;
    wire N__21432;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21385;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21358;
    wire N__21357;
    wire N__21354;
    wire N__21353;
    wire N__21350;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21324;
    wire N__21321;
    wire N__21320;
    wire N__21315;
    wire N__21314;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21301;
    wire N__21292;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21282;
    wire N__21279;
    wire N__21276;
    wire N__21271;
    wire N__21268;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21214;
    wire N__21211;
    wire N__21208;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21172;
    wire N__21169;
    wire N__21166;
    wire N__21163;
    wire N__21160;
    wire N__21157;
    wire N__21156;
    wire N__21155;
    wire N__21154;
    wire N__21153;
    wire N__21152;
    wire N__21151;
    wire N__21150;
    wire N__21147;
    wire N__21146;
    wire N__21145;
    wire N__21144;
    wire N__21139;
    wire N__21134;
    wire N__21127;
    wire N__21126;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21114;
    wire N__21113;
    wire N__21112;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21102;
    wire N__21101;
    wire N__21100;
    wire N__21099;
    wire N__21098;
    wire N__21097;
    wire N__21096;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21077;
    wire N__21076;
    wire N__21075;
    wire N__21074;
    wire N__21073;
    wire N__21072;
    wire N__21065;
    wire N__21062;
    wire N__21053;
    wire N__21048;
    wire N__21045;
    wire N__21036;
    wire N__21025;
    wire N__21010;
    wire N__21007;
    wire N__21006;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20998;
    wire N__20997;
    wire N__20996;
    wire N__20993;
    wire N__20988;
    wire N__20987;
    wire N__20986;
    wire N__20985;
    wire N__20984;
    wire N__20979;
    wire N__20978;
    wire N__20977;
    wire N__20976;
    wire N__20973;
    wire N__20972;
    wire N__20971;
    wire N__20970;
    wire N__20969;
    wire N__20968;
    wire N__20967;
    wire N__20966;
    wire N__20965;
    wire N__20962;
    wire N__20959;
    wire N__20950;
    wire N__20949;
    wire N__20948;
    wire N__20947;
    wire N__20944;
    wire N__20941;
    wire N__20938;
    wire N__20935;
    wire N__20932;
    wire N__20931;
    wire N__20930;
    wire N__20929;
    wire N__20926;
    wire N__20925;
    wire N__20922;
    wire N__20911;
    wire N__20908;
    wire N__20901;
    wire N__20896;
    wire N__20893;
    wire N__20892;
    wire N__20891;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20876;
    wire N__20875;
    wire N__20874;
    wire N__20873;
    wire N__20872;
    wire N__20869;
    wire N__20860;
    wire N__20855;
    wire N__20852;
    wire N__20847;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20829;
    wire N__20824;
    wire N__20815;
    wire N__20812;
    wire N__20801;
    wire N__20788;
    wire N__20785;
    wire N__20784;
    wire N__20781;
    wire N__20778;
    wire N__20773;
    wire N__20772;
    wire N__20771;
    wire N__20770;
    wire N__20767;
    wire N__20762;
    wire N__20759;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20695;
    wire N__20694;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20677;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20665;
    wire N__20662;
    wire N__20661;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20632;
    wire N__20629;
    wire N__20626;
    wire N__20625;
    wire N__20622;
    wire N__20621;
    wire N__20618;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20610;
    wire N__20607;
    wire N__20606;
    wire N__20605;
    wire N__20602;
    wire N__20597;
    wire N__20596;
    wire N__20595;
    wire N__20594;
    wire N__20593;
    wire N__20592;
    wire N__20591;
    wire N__20590;
    wire N__20589;
    wire N__20588;
    wire N__20587;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20559;
    wire N__20550;
    wire N__20547;
    wire N__20542;
    wire N__20541;
    wire N__20540;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20515;
    wire N__20508;
    wire N__20501;
    wire N__20496;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20446;
    wire N__20445;
    wire N__20440;
    wire N__20437;
    wire N__20434;
    wire N__20431;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20419;
    wire N__20418;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20395;
    wire N__20394;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20382;
    wire N__20381;
    wire N__20374;
    wire N__20373;
    wire N__20372;
    wire N__20371;
    wire N__20370;
    wire N__20369;
    wire N__20368;
    wire N__20367;
    wire N__20366;
    wire N__20365;
    wire N__20364;
    wire N__20361;
    wire N__20352;
    wire N__20351;
    wire N__20350;
    wire N__20349;
    wire N__20348;
    wire N__20343;
    wire N__20336;
    wire N__20333;
    wire N__20332;
    wire N__20327;
    wire N__20326;
    wire N__20317;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20291;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20266;
    wire N__20263;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20251;
    wire N__20250;
    wire N__20245;
    wire N__20242;
    wire N__20239;
    wire N__20236;
    wire N__20233;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20221;
    wire N__20218;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20197;
    wire N__20196;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20166;
    wire N__20161;
    wire N__20160;
    wire N__20155;
    wire N__20152;
    wire N__20149;
    wire N__20146;
    wire N__20143;
    wire N__20142;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20130;
    wire N__20125;
    wire N__20124;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20086;
    wire N__20083;
    wire N__20082;
    wire N__20077;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20067;
    wire N__20064;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20050;
    wire N__20049;
    wire N__20044;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20013;
    wire N__20012;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19990;
    wire N__19989;
    wire N__19986;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19966;
    wire N__19965;
    wire N__19962;
    wire N__19959;
    wire N__19954;
    wire N__19953;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19927;
    wire N__19926;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19905;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19897;
    wire N__19896;
    wire N__19895;
    wire N__19892;
    wire N__19891;
    wire N__19890;
    wire N__19889;
    wire N__19888;
    wire N__19887;
    wire N__19886;
    wire N__19883;
    wire N__19878;
    wire N__19875;
    wire N__19872;
    wire N__19867;
    wire N__19862;
    wire N__19859;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19841;
    wire N__19828;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19816;
    wire N__19813;
    wire N__19810;
    wire N__19807;
    wire N__19806;
    wire N__19803;
    wire N__19800;
    wire N__19795;
    wire N__19792;
    wire N__19789;
    wire N__19788;
    wire N__19783;
    wire N__19780;
    wire N__19779;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19749;
    wire N__19744;
    wire N__19741;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19729;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19708;
    wire N__19705;
    wire N__19702;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19669;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19656;
    wire N__19653;
    wire N__19652;
    wire N__19649;
    wire N__19642;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19614;
    wire N__19611;
    wire N__19610;
    wire N__19607;
    wire N__19606;
    wire N__19605;
    wire N__19602;
    wire N__19599;
    wire N__19592;
    wire N__19585;
    wire N__19582;
    wire N__19579;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19567;
    wire N__19564;
    wire N__19561;
    wire N__19560;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19548;
    wire N__19545;
    wire N__19544;
    wire N__19541;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19479;
    wire N__19478;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19441;
    wire N__19438;
    wire N__19437;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19423;
    wire N__19422;
    wire N__19421;
    wire N__19418;
    wire N__19417;
    wire N__19416;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19402;
    wire N__19399;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19317;
    wire N__19314;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19287;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19260;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19237;
    wire N__19234;
    wire N__19231;
    wire N__19228;
    wire N__19225;
    wire N__19224;
    wire N__19221;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19201;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19188;
    wire N__19185;
    wire N__19182;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19148;
    wire N__19143;
    wire N__19140;
    wire N__19135;
    wire N__19132;
    wire N__19129;
    wire N__19126;
    wire N__19125;
    wire N__19122;
    wire N__19119;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19077;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19060;
    wire N__19057;
    wire N__19054;
    wire N__19051;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19011;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18990;
    wire N__18985;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18960;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18937;
    wire N__18934;
    wire N__18931;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18918;
    wire N__18915;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18898;
    wire N__18895;
    wire N__18892;
    wire N__18889;
    wire N__18888;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18873;
    wire N__18868;
    wire N__18865;
    wire N__18862;
    wire N__18859;
    wire N__18856;
    wire N__18853;
    wire N__18852;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18835;
    wire N__18832;
    wire N__18829;
    wire N__18826;
    wire N__18823;
    wire N__18822;
    wire N__18817;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18807;
    wire N__18804;
    wire N__18801;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18789;
    wire N__18786;
    wire N__18781;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18751;
    wire N__18750;
    wire N__18747;
    wire N__18746;
    wire N__18745;
    wire N__18744;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18727;
    wire N__18724;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18702;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18678;
    wire N__18675;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18657;
    wire N__18652;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18636;
    wire N__18631;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18619;
    wire N__18618;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18591;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18568;
    wire N__18565;
    wire N__18562;
    wire N__18559;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18541;
    wire N__18538;
    wire N__18535;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18523;
    wire N__18520;
    wire N__18519;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18507;
    wire N__18502;
    wire N__18501;
    wire N__18500;
    wire N__18497;
    wire N__18492;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18456;
    wire N__18453;
    wire N__18450;
    wire N__18449;
    wire N__18444;
    wire N__18441;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18420;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18400;
    wire N__18397;
    wire N__18394;
    wire N__18391;
    wire N__18388;
    wire N__18385;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18373;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18361;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18349;
    wire N__18346;
    wire N__18343;
    wire N__18342;
    wire N__18339;
    wire N__18338;
    wire N__18335;
    wire N__18334;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18320;
    wire N__18313;
    wire N__18310;
    wire N__18309;
    wire N__18308;
    wire N__18307;
    wire N__18306;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18283;
    wire N__18282;
    wire N__18279;
    wire N__18278;
    wire N__18275;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18259;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18251;
    wire N__18246;
    wire N__18243;
    wire N__18238;
    wire N__18235;
    wire N__18234;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18208;
    wire N__18205;
    wire N__18202;
    wire N__18201;
    wire N__18198;
    wire N__18197;
    wire N__18194;
    wire N__18187;
    wire N__18184;
    wire N__18181;
    wire N__18178;
    wire N__18175;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18163;
    wire N__18160;
    wire N__18157;
    wire N__18154;
    wire N__18151;
    wire N__18148;
    wire N__18145;
    wire N__18142;
    wire N__18139;
    wire N__18136;
    wire N__18133;
    wire N__18130;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18103;
    wire N__18100;
    wire N__18097;
    wire N__18094;
    wire N__18091;
    wire N__18090;
    wire N__18087;
    wire N__18086;
    wire N__18083;
    wire N__18082;
    wire N__18081;
    wire N__18078;
    wire N__18073;
    wire N__18070;
    wire N__18067;
    wire N__18058;
    wire N__18055;
    wire N__18052;
    wire N__18049;
    wire N__18046;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18034;
    wire N__18031;
    wire N__18028;
    wire N__18025;
    wire N__18022;
    wire N__18019;
    wire N__18016;
    wire N__18013;
    wire N__18010;
    wire N__18007;
    wire N__18004;
    wire N__18001;
    wire N__17998;
    wire N__17997;
    wire N__17996;
    wire N__17993;
    wire N__17992;
    wire N__17991;
    wire N__17988;
    wire N__17985;
    wire N__17978;
    wire N__17971;
    wire N__17970;
    wire N__17967;
    wire N__17966;
    wire N__17963;
    wire N__17956;
    wire N__17953;
    wire N__17950;
    wire N__17947;
    wire N__17944;
    wire N__17941;
    wire N__17938;
    wire N__17935;
    wire N__17932;
    wire N__17929;
    wire N__17926;
    wire N__17923;
    wire N__17920;
    wire N__17919;
    wire N__17916;
    wire N__17915;
    wire N__17912;
    wire N__17911;
    wire N__17908;
    wire N__17903;
    wire N__17900;
    wire N__17893;
    wire N__17890;
    wire N__17887;
    wire N__17884;
    wire N__17881;
    wire N__17878;
    wire N__17875;
    wire N__17872;
    wire N__17869;
    wire N__17866;
    wire N__17863;
    wire N__17860;
    wire N__17857;
    wire N__17854;
    wire N__17853;
    wire N__17848;
    wire N__17845;
    wire N__17842;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17830;
    wire N__17827;
    wire N__17824;
    wire N__17823;
    wire N__17822;
    wire N__17821;
    wire N__17820;
    wire N__17819;
    wire N__17818;
    wire N__17817;
    wire N__17816;
    wire N__17813;
    wire N__17812;
    wire N__17803;
    wire N__17796;
    wire N__17795;
    wire N__17794;
    wire N__17793;
    wire N__17792;
    wire N__17791;
    wire N__17790;
    wire N__17789;
    wire N__17782;
    wire N__17777;
    wire N__17770;
    wire N__17761;
    wire N__17752;
    wire N__17749;
    wire N__17748;
    wire N__17745;
    wire N__17742;
    wire N__17737;
    wire N__17734;
    wire N__17731;
    wire N__17728;
    wire N__17725;
    wire N__17722;
    wire N__17721;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17706;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17692;
    wire N__17691;
    wire N__17688;
    wire N__17685;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17673;
    wire N__17670;
    wire N__17667;
    wire N__17662;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17646;
    wire N__17643;
    wire N__17640;
    wire N__17637;
    wire N__17632;
    wire N__17629;
    wire N__17628;
    wire N__17625;
    wire N__17622;
    wire N__17619;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17605;
    wire N__17602;
    wire N__17601;
    wire N__17598;
    wire N__17595;
    wire N__17592;
    wire N__17587;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17575;
    wire N__17574;
    wire N__17571;
    wire N__17568;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17551;
    wire N__17548;
    wire N__17545;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17533;
    wire N__17532;
    wire N__17529;
    wire N__17526;
    wire N__17523;
    wire N__17518;
    wire N__17515;
    wire N__17514;
    wire N__17511;
    wire N__17508;
    wire N__17505;
    wire N__17500;
    wire N__17497;
    wire N__17496;
    wire N__17493;
    wire N__17490;
    wire N__17487;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17461;
    wire N__17458;
    wire N__17457;
    wire N__17454;
    wire N__17451;
    wire N__17448;
    wire N__17443;
    wire N__17440;
    wire N__17437;
    wire N__17436;
    wire N__17433;
    wire N__17430;
    wire N__17427;
    wire N__17422;
    wire N__17419;
    wire N__17418;
    wire N__17415;
    wire N__17412;
    wire N__17409;
    wire N__17404;
    wire N__17401;
    wire N__17398;
    wire N__17397;
    wire N__17394;
    wire N__17391;
    wire N__17388;
    wire N__17383;
    wire N__17380;
    wire N__17379;
    wire N__17376;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17359;
    wire N__17356;
    wire N__17355;
    wire N__17354;
    wire N__17351;
    wire N__17346;
    wire N__17341;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17311;
    wire N__17308;
    wire N__17307;
    wire N__17304;
    wire N__17301;
    wire N__17300;
    wire N__17297;
    wire N__17292;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17277;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17254;
    wire N__17253;
    wire N__17250;
    wire N__17247;
    wire N__17244;
    wire N__17239;
    wire N__17236;
    wire N__17233;
    wire N__17230;
    wire N__17227;
    wire N__17226;
    wire N__17223;
    wire N__17220;
    wire N__17217;
    wire N__17212;
    wire N__17209;
    wire N__17208;
    wire N__17205;
    wire N__17202;
    wire N__17199;
    wire N__17194;
    wire N__17191;
    wire N__17190;
    wire N__17187;
    wire N__17184;
    wire N__17181;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17166;
    wire N__17163;
    wire N__17160;
    wire N__17157;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17142;
    wire N__17139;
    wire N__17136;
    wire N__17133;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17092;
    wire N__17089;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17047;
    wire N__17044;
    wire N__17041;
    wire N__17040;
    wire N__17037;
    wire N__17034;
    wire N__17033;
    wire N__17030;
    wire N__17025;
    wire N__17020;
    wire N__17017;
    wire N__17014;
    wire N__17011;
    wire N__17008;
    wire N__17005;
    wire N__17002;
    wire N__16999;
    wire N__16996;
    wire N__16993;
    wire N__16992;
    wire N__16989;
    wire N__16986;
    wire N__16983;
    wire N__16978;
    wire N__16975;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16935;
    wire N__16934;
    wire N__16933;
    wire N__16932;
    wire N__16931;
    wire N__16930;
    wire N__16929;
    wire N__16928;
    wire N__16927;
    wire N__16926;
    wire N__16925;
    wire N__16924;
    wire N__16923;
    wire N__16922;
    wire N__16921;
    wire N__16920;
    wire N__16919;
    wire N__16918;
    wire N__16917;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16897;
    wire N__16896;
    wire N__16893;
    wire N__16886;
    wire N__16883;
    wire N__16876;
    wire N__16873;
    wire N__16870;
    wire N__16861;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16831;
    wire N__16826;
    wire N__16815;
    wire N__16810;
    wire N__16807;
    wire N__16804;
    wire N__16795;
    wire N__16792;
    wire N__16789;
    wire N__16786;
    wire N__16783;
    wire N__16780;
    wire N__16777;
    wire N__16774;
    wire N__16771;
    wire N__16768;
    wire N__16765;
    wire N__16762;
    wire N__16759;
    wire N__16756;
    wire N__16755;
    wire N__16752;
    wire N__16751;
    wire N__16748;
    wire N__16741;
    wire N__16738;
    wire N__16735;
    wire N__16732;
    wire N__16729;
    wire N__16726;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16714;
    wire N__16711;
    wire N__16708;
    wire N__16705;
    wire N__16702;
    wire N__16699;
    wire N__16696;
    wire N__16693;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16681;
    wire N__16678;
    wire N__16675;
    wire N__16672;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16662;
    wire N__16659;
    wire N__16658;
    wire N__16655;
    wire N__16648;
    wire N__16645;
    wire N__16642;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16630;
    wire N__16627;
    wire N__16624;
    wire N__16621;
    wire N__16618;
    wire N__16615;
    wire N__16612;
    wire N__16609;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16597;
    wire N__16594;
    wire N__16593;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16576;
    wire N__16573;
    wire N__16572;
    wire N__16567;
    wire N__16564;
    wire N__16561;
    wire N__16558;
    wire N__16555;
    wire N__16552;
    wire N__16549;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16537;
    wire N__16536;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16516;
    wire N__16513;
    wire N__16510;
    wire N__16509;
    wire N__16508;
    wire N__16503;
    wire N__16500;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16486;
    wire N__16485;
    wire N__16484;
    wire N__16483;
    wire N__16480;
    wire N__16473;
    wire N__16468;
    wire N__16465;
    wire N__16462;
    wire N__16459;
    wire N__16456;
    wire N__16453;
    wire N__16450;
    wire N__16447;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16435;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16405;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16397;
    wire N__16394;
    wire N__16389;
    wire N__16384;
    wire N__16383;
    wire N__16380;
    wire N__16377;
    wire N__16372;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16360;
    wire N__16359;
    wire N__16356;
    wire N__16353;
    wire N__16350;
    wire N__16345;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16333;
    wire N__16332;
    wire N__16329;
    wire N__16326;
    wire N__16321;
    wire N__16320;
    wire N__16317;
    wire N__16314;
    wire N__16309;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16299;
    wire N__16294;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16282;
    wire N__16281;
    wire N__16278;
    wire N__16275;
    wire N__16270;
    wire N__16269;
    wire N__16266;
    wire N__16263;
    wire N__16258;
    wire N__16257;
    wire N__16254;
    wire N__16251;
    wire N__16248;
    wire N__16243;
    wire N__16242;
    wire N__16239;
    wire N__16236;
    wire N__16231;
    wire N__16228;
    wire N__16227;
    wire N__16222;
    wire N__16219;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16192;
    wire N__16191;
    wire N__16190;
    wire N__16189;
    wire N__16188;
    wire N__16181;
    wire N__16176;
    wire N__16171;
    wire N__16168;
    wire N__16165;
    wire N__16164;
    wire N__16163;
    wire N__16162;
    wire N__16161;
    wire N__16150;
    wire N__16147;
    wire N__16146;
    wire N__16145;
    wire N__16144;
    wire N__16141;
    wire N__16140;
    wire N__16129;
    wire N__16126;
    wire N__16123;
    wire N__16120;
    wire N__16119;
    wire N__16118;
    wire N__16117;
    wire N__16110;
    wire N__16107;
    wire N__16104;
    wire N__16099;
    wire N__16096;
    wire N__16095;
    wire N__16090;
    wire N__16087;
    wire N__16084;
    wire N__16081;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16069;
    wire N__16066;
    wire N__16063;
    wire N__16060;
    wire N__16059;
    wire N__16056;
    wire N__16053;
    wire N__16048;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16036;
    wire N__16035;
    wire N__16032;
    wire N__16029;
    wire N__16026;
    wire N__16021;
    wire N__16020;
    wire N__16017;
    wire N__16014;
    wire N__16009;
    wire N__16008;
    wire N__16005;
    wire N__16002;
    wire N__15997;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15985;
    wire N__15984;
    wire N__15981;
    wire N__15978;
    wire N__15975;
    wire N__15970;
    wire N__15969;
    wire N__15966;
    wire N__15963;
    wire N__15958;
    wire N__15957;
    wire N__15954;
    wire N__15951;
    wire N__15946;
    wire N__15945;
    wire N__15942;
    wire N__15939;
    wire N__15934;
    wire N__15933;
    wire N__15930;
    wire N__15927;
    wire N__15924;
    wire N__15919;
    wire N__15918;
    wire N__15915;
    wire N__15912;
    wire N__15907;
    wire N__15906;
    wire N__15905;
    wire N__15904;
    wire N__15903;
    wire N__15902;
    wire N__15901;
    wire N__15892;
    wire N__15885;
    wire N__15884;
    wire N__15883;
    wire N__15882;
    wire N__15879;
    wire N__15876;
    wire N__15875;
    wire N__15874;
    wire N__15873;
    wire N__15872;
    wire N__15871;
    wire N__15870;
    wire N__15869;
    wire N__15866;
    wire N__15863;
    wire N__15860;
    wire N__15855;
    wire N__15848;
    wire N__15839;
    wire N__15826;
    wire N__15825;
    wire N__15824;
    wire N__15823;
    wire N__15822;
    wire N__15819;
    wire N__15814;
    wire N__15811;
    wire N__15808;
    wire N__15799;
    wire N__15796;
    wire N__15793;
    wire N__15790;
    wire N__15789;
    wire N__15786;
    wire N__15785;
    wire N__15784;
    wire N__15783;
    wire N__15780;
    wire N__15777;
    wire N__15770;
    wire N__15763;
    wire N__15762;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15744;
    wire N__15739;
    wire N__15738;
    wire N__15735;
    wire N__15732;
    wire N__15727;
    wire N__15726;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15712;
    wire N__15709;
    wire N__15708;
    wire N__15705;
    wire N__15700;
    wire N__15699;
    wire N__15696;
    wire N__15693;
    wire N__15688;
    wire N__15687;
    wire N__15682;
    wire N__15679;
    wire N__15676;
    wire N__15673;
    wire N__15670;
    wire N__15669;
    wire N__15664;
    wire N__15663;
    wire N__15660;
    wire N__15657;
    wire N__15652;
    wire N__15651;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15607;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15595;
    wire N__15592;
    wire N__15591;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15579;
    wire N__15576;
    wire N__15573;
    wire N__15568;
    wire N__15567;
    wire N__15562;
    wire N__15559;
    wire N__15556;
    wire N__15553;
    wire N__15550;
    wire N__15547;
    wire N__15546;
    wire N__15541;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15528;
    wire N__15523;
    wire N__15520;
    wire N__15517;
    wire N__15514;
    wire N__15511;
    wire N__15508;
    wire N__15507;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15480;
    wire N__15479;
    wire N__15476;
    wire N__15471;
    wire N__15468;
    wire N__15463;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15429;
    wire N__15428;
    wire N__15425;
    wire N__15420;
    wire N__15415;
    wire N__15414;
    wire N__15413;
    wire N__15412;
    wire N__15409;
    wire N__15408;
    wire N__15407;
    wire N__15404;
    wire N__15401;
    wire N__15400;
    wire N__15399;
    wire N__15396;
    wire N__15395;
    wire N__15392;
    wire N__15389;
    wire N__15380;
    wire N__15377;
    wire N__15376;
    wire N__15373;
    wire N__15370;
    wire N__15367;
    wire N__15362;
    wire N__15357;
    wire N__15354;
    wire N__15343;
    wire N__15340;
    wire N__15339;
    wire N__15334;
    wire N__15331;
    wire N__15330;
    wire N__15325;
    wire N__15322;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15310;
    wire N__15309;
    wire N__15306;
    wire N__15305;
    wire N__15304;
    wire N__15303;
    wire N__15302;
    wire N__15301;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15293;
    wire N__15284;
    wire N__15277;
    wire N__15274;
    wire N__15271;
    wire N__15268;
    wire N__15259;
    wire N__15256;
    wire N__15255;
    wire N__15254;
    wire N__15251;
    wire N__15250;
    wire N__15247;
    wire N__15244;
    wire N__15243;
    wire N__15240;
    wire N__15237;
    wire N__15230;
    wire N__15223;
    wire N__15222;
    wire N__15221;
    wire N__15220;
    wire N__15219;
    wire N__15216;
    wire N__15207;
    wire N__15202;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15190;
    wire N__15187;
    wire N__15184;
    wire N__15181;
    wire N__15178;
    wire N__15175;
    wire N__15172;
    wire N__15169;
    wire N__15166;
    wire N__15163;
    wire N__15160;
    wire N__15157;
    wire N__15156;
    wire N__15153;
    wire N__15150;
    wire N__15145;
    wire N__15144;
    wire N__15141;
    wire N__15138;
    wire N__15133;
    wire N__15132;
    wire N__15129;
    wire N__15126;
    wire N__15123;
    wire N__15118;
    wire N__15117;
    wire N__15114;
    wire N__15111;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15093;
    wire N__15090;
    wire N__15087;
    wire N__15082;
    wire N__15081;
    wire N__15078;
    wire N__15075;
    wire N__15070;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15055;
    wire N__15054;
    wire N__15051;
    wire N__15050;
    wire N__15045;
    wire N__15042;
    wire N__15037;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15024;
    wire N__15021;
    wire N__15018;
    wire N__15017;
    wire N__15012;
    wire N__15011;
    wire N__15010;
    wire N__15009;
    wire N__15008;
    wire N__15007;
    wire N__15006;
    wire N__15005;
    wire N__15004;
    wire N__15003;
    wire N__15000;
    wire N__14999;
    wire N__14998;
    wire N__14997;
    wire N__14996;
    wire N__14995;
    wire N__14992;
    wire N__14983;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14957;
    wire N__14950;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14925;
    wire N__14924;
    wire N__14917;
    wire N__14914;
    wire N__14911;
    wire N__14908;
    wire N__14907;
    wire N__14904;
    wire N__14901;
    wire N__14898;
    wire N__14893;
    wire N__14890;
    wire N__14887;
    wire N__14884;
    wire N__14883;
    wire N__14878;
    wire N__14875;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14859;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14845;
    wire N__14844;
    wire N__14841;
    wire N__14838;
    wire N__14835;
    wire N__14830;
    wire N__14829;
    wire N__14826;
    wire N__14823;
    wire N__14818;
    wire N__14815;
    wire N__14814;
    wire N__14811;
    wire N__14808;
    wire N__14803;
    wire N__14802;
    wire N__14801;
    wire N__14798;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14776;
    wire N__14775;
    wire N__14772;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14752;
    wire N__14749;
    wire N__14748;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14725;
    wire N__14724;
    wire N__14723;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14709;
    wire N__14706;
    wire N__14703;
    wire N__14698;
    wire N__14695;
    wire N__14692;
    wire N__14689;
    wire N__14688;
    wire N__14685;
    wire N__14682;
    wire N__14677;
    wire N__14676;
    wire N__14673;
    wire N__14670;
    wire N__14665;
    wire N__14662;
    wire N__14661;
    wire N__14656;
    wire N__14653;
    wire N__14650;
    wire N__14649;
    wire N__14646;
    wire N__14643;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14619;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14609;
    wire N__14602;
    wire N__14601;
    wire N__14596;
    wire N__14593;
    wire N__14590;
    wire N__14587;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14577;
    wire N__14574;
    wire N__14571;
    wire N__14566;
    wire N__14565;
    wire N__14562;
    wire N__14559;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14530;
    wire N__14529;
    wire N__14528;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14514;
    wire N__14513;
    wire N__14508;
    wire N__14505;
    wire N__14500;
    wire N__14499;
    wire N__14496;
    wire N__14493;
    wire N__14488;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14478;
    wire N__14473;
    wire N__14470;
    wire N__14467;
    wire N__14464;
    wire N__14461;
    wire N__14460;
    wire N__14457;
    wire N__14454;
    wire N__14449;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14433;
    wire N__14432;
    wire N__14429;
    wire N__14424;
    wire N__14419;
    wire N__14416;
    wire N__14415;
    wire N__14412;
    wire N__14409;
    wire N__14404;
    wire N__14401;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14359;
    wire N__14356;
    wire N__14353;
    wire N__14350;
    wire N__14347;
    wire N__14344;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14332;
    wire N__14329;
    wire N__14326;
    wire N__14323;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14313;
    wire N__14310;
    wire N__14307;
    wire N__14304;
    wire N__14299;
    wire N__14298;
    wire N__14293;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14283;
    wire N__14280;
    wire N__14277;
    wire N__14274;
    wire N__14269;
    wire N__14268;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14254;
    wire N__14253;
    wire N__14250;
    wire N__14247;
    wire N__14244;
    wire N__14239;
    wire N__14238;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14224;
    wire N__14221;
    wire N__14220;
    wire N__14217;
    wire N__14214;
    wire N__14211;
    wire N__14206;
    wire N__14205;
    wire N__14202;
    wire N__14197;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14184;
    wire N__14181;
    wire N__14178;
    wire N__14173;
    wire N__14170;
    wire N__14167;
    wire N__14166;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14140;
    wire N__14139;
    wire N__14136;
    wire N__14133;
    wire N__14128;
    wire N__14125;
    wire N__14122;
    wire N__14121;
    wire N__14118;
    wire N__14115;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14103;
    wire N__14098;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14086;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14062;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14029;
    wire N__14028;
    wire N__14027;
    wire N__14024;
    wire N__14019;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__13999;
    wire N__13998;
    wire N__13995;
    wire N__13992;
    wire N__13989;
    wire N__13984;
    wire N__13981;
    wire N__13978;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13953;
    wire N__13952;
    wire N__13949;
    wire N__13944;
    wire N__13939;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13924;
    wire N__13923;
    wire N__13922;
    wire N__13919;
    wire N__13914;
    wire N__13909;
    wire N__13906;
    wire N__13903;
    wire N__13900;
    wire N__13897;
    wire N__13894;
    wire N__13891;
    wire N__13888;
    wire N__13885;
    wire N__13882;
    wire N__13879;
    wire N__13878;
    wire N__13875;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13858;
    wire N__13857;
    wire N__13854;
    wire N__13851;
    wire N__13846;
    wire N__13843;
    wire N__13842;
    wire N__13839;
    wire N__13836;
    wire N__13831;
    wire N__13828;
    wire N__13825;
    wire N__13824;
    wire N__13821;
    wire N__13818;
    wire N__13813;
    wire N__13810;
    wire N__13809;
    wire N__13806;
    wire N__13803;
    wire N__13798;
    wire N__13795;
    wire N__13794;
    wire N__13791;
    wire N__13788;
    wire N__13783;
    wire N__13780;
    wire N__13779;
    wire N__13774;
    wire N__13771;
    wire N__13768;
    wire N__13765;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13752;
    wire N__13747;
    wire N__13744;
    wire N__13741;
    wire N__13738;
    wire N__13735;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13723;
    wire N__13720;
    wire N__13717;
    wire N__13714;
    wire N__13713;
    wire N__13708;
    wire N__13705;
    wire N__13702;
    wire N__13699;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13687;
    wire N__13684;
    wire N__13681;
    wire N__13680;
    wire N__13677;
    wire N__13674;
    wire N__13673;
    wire N__13668;
    wire N__13665;
    wire N__13660;
    wire N__13659;
    wire N__13654;
    wire N__13651;
    wire N__13648;
    wire N__13645;
    wire N__13644;
    wire N__13641;
    wire N__13638;
    wire N__13633;
    wire N__13632;
    wire N__13627;
    wire N__13624;
    wire N__13621;
    wire N__13618;
    wire N__13615;
    wire N__13612;
    wire N__13609;
    wire N__13606;
    wire N__13603;
    wire N__13600;
    wire N__13599;
    wire N__13594;
    wire N__13591;
    wire N__13588;
    wire N__13585;
    wire N__13582;
    wire N__13579;
    wire VCCG0;
    wire \PCH_PWRGD.count_rst_6 ;
    wire \PCH_PWRGD.count_rst_6_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_8_cascade_ ;
    wire \PCH_PWRGD.count_0_8 ;
    wire \PCH_PWRGD.count_rst_7_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_7_cascade_ ;
    wire \PCH_PWRGD.count_0_7 ;
    wire bfn_1_2_0_;
    wire \PCH_PWRGD.un2_count_1_cry_1 ;
    wire \PCH_PWRGD.un2_count_1_cry_2 ;
    wire \PCH_PWRGD.un2_count_1_cry_3 ;
    wire \PCH_PWRGD.un2_count_1_cry_4 ;
    wire \PCH_PWRGD.un2_count_1_cry_5 ;
    wire \PCH_PWRGD.countZ0Z_7 ;
    wire \PCH_PWRGD.un2_count_1_cry_6_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_6 ;
    wire \PCH_PWRGD.un2_count_1_axb_8 ;
    wire \PCH_PWRGD.un2_count_1_cry_7_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_7 ;
    wire \PCH_PWRGD.un2_count_1_cry_8 ;
    wire bfn_1_3_0_;
    wire \PCH_PWRGD.un2_count_1_cry_9 ;
    wire \PCH_PWRGD.un2_count_1_cry_10 ;
    wire \PCH_PWRGD.un2_count_1_cry_11 ;
    wire \PCH_PWRGD.un2_count_1_cry_12 ;
    wire \PCH_PWRGD.un2_count_1_cry_13 ;
    wire \PCH_PWRGD.un2_count_1_cry_14 ;
    wire \PCH_PWRGD.un2_count_1_axb_14 ;
    wire \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8PZ0Z7 ;
    wire \PCH_PWRGD.count_0_13 ;
    wire \PCH_PWRGD.count_rst_11_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_cry_2_THRU_CO ;
    wire \PCH_PWRGD.countZ0Z_3_cascade_ ;
    wire \PCH_PWRGD.count_0_3 ;
    wire \PCH_PWRGD.count_rst_10_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_4_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_cry_3_THRU_CO ;
    wire \PCH_PWRGD.count_0_4 ;
    wire \HDA_STRAP.un4_count_9_cascade_ ;
    wire \HDA_STRAP.un4_count_10_cascade_ ;
    wire \HDA_STRAP.un4_count_13 ;
    wire \HDA_STRAP.un4_count_cascade_ ;
    wire \HDA_STRAP.countZ0Z_0 ;
    wire bfn_1_6_0_;
    wire \HDA_STRAP.countZ0Z_1 ;
    wire \HDA_STRAP.un1_count_1_cry_0 ;
    wire \HDA_STRAP.countZ0Z_2 ;
    wire \HDA_STRAP.un1_count_1_cry_1 ;
    wire \HDA_STRAP.countZ0Z_3 ;
    wire \HDA_STRAP.un1_count_1_cry_2 ;
    wire \HDA_STRAP.countZ0Z_4 ;
    wire \HDA_STRAP.un1_count_1_cry_3 ;
    wire \HDA_STRAP.countZ0Z_5 ;
    wire \HDA_STRAP.un1_count_1_cry_4 ;
    wire \HDA_STRAP.un1_count_1_cry_5 ;
    wire \HDA_STRAP.un1_count_1_cry_6 ;
    wire \HDA_STRAP.un1_count_1_cry_7 ;
    wire bfn_1_7_0_;
    wire \HDA_STRAP.un1_count_1_cry_8 ;
    wire \HDA_STRAP.countZ0Z_10 ;
    wire \HDA_STRAP.un1_count_1_cry_9_THRU_CO ;
    wire \HDA_STRAP.un1_count_1_cry_9 ;
    wire \HDA_STRAP.countZ0Z_11 ;
    wire \HDA_STRAP.un1_count_1_cry_10_THRU_CO ;
    wire \HDA_STRAP.un1_count_1_cry_10 ;
    wire \HDA_STRAP.un1_count_1_cry_11 ;
    wire \HDA_STRAP.un1_count_1_cry_12 ;
    wire \HDA_STRAP.un1_count_1_cry_13 ;
    wire \HDA_STRAP.un1_count_1_cry_14 ;
    wire \HDA_STRAP.un1_count_1_cry_15 ;
    wire \HDA_STRAP.countZ0Z_16 ;
    wire \HDA_STRAP.un1_count_1_cry_15_THRU_CO ;
    wire bfn_1_8_0_;
    wire \HDA_STRAP.un1_count_1_cry_16 ;
    wire \HDA_STRAP.countZ0Z_17 ;
    wire \POWERLED.count_clk_0_4 ;
    wire \POWERLED.count_clk_0_15 ;
    wire \POWERLED.count_clk_0_10 ;
    wire \POWERLED.un1_dutycycle_168_0_0_o2_1_4_cascade_ ;
    wire \POWERLED.count_clk_0_14 ;
    wire \POWERLED.count_clk_0_11 ;
    wire \POWERLED.count_clk_0_12 ;
    wire bfn_1_11_0_;
    wire \POWERLED.un1_count_clk_2_cry_1 ;
    wire \POWERLED.un1_count_clk_2_cry_2 ;
    wire \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_3 ;
    wire \POWERLED.un1_count_clk_2_cry_4 ;
    wire \POWERLED.un1_count_clk_2_cry_5 ;
    wire \POWERLED.un1_count_clk_2_cry_6 ;
    wire \POWERLED.un1_count_clk_2_cry_7 ;
    wire \POWERLED.un1_count_clk_2_cry_8_cZ0 ;
    wire bfn_1_12_0_;
    wire \POWERLED.count_clkZ0Z_10 ;
    wire \POWERLED.count_clk_1_10 ;
    wire \POWERLED.un1_count_clk_2_cry_9_cZ0 ;
    wire \POWERLED.count_clkZ0Z_11 ;
    wire \POWERLED.count_clk_1_11 ;
    wire \POWERLED.un1_count_clk_2_cry_10 ;
    wire \POWERLED.count_clkZ0Z_12 ;
    wire \POWERLED.count_clk_1_12 ;
    wire \POWERLED.un1_count_clk_2_cry_11 ;
    wire \POWERLED.un1_count_clk_2_cry_12 ;
    wire \POWERLED.count_clkZ0Z_14 ;
    wire \POWERLED.count_clk_1_14 ;
    wire \POWERLED.un1_count_clk_2_cry_13 ;
    wire \POWERLED.count_clkZ0Z_15 ;
    wire \POWERLED.un1_count_clk_2_cry_14 ;
    wire \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ;
    wire \POWERLED.count_clk_0_13 ;
    wire \POWERLED.count_clk_1_13 ;
    wire \POWERLED.count_clkZ0Z_13 ;
    wire bfn_1_13_0_;
    wire \COUNTER.counter_1_cry_1 ;
    wire \COUNTER.counter_1_cry_2 ;
    wire \COUNTER.counter_1_cry_3 ;
    wire \COUNTER.counter_1_cry_4 ;
    wire \COUNTER.counter_1_cry_5 ;
    wire \COUNTER.counter_1_cry_6 ;
    wire \COUNTER.counter_1_cry_7 ;
    wire \COUNTER.counter_1_cry_8 ;
    wire bfn_1_14_0_;
    wire \COUNTER.counter_1_cry_9 ;
    wire \COUNTER.counter_1_cry_10 ;
    wire \COUNTER.counter_1_cry_11 ;
    wire \COUNTER.counter_1_cry_12 ;
    wire \COUNTER.counter_1_cry_13 ;
    wire \COUNTER.counter_1_cry_14 ;
    wire \COUNTER.counter_1_cry_15 ;
    wire \COUNTER.counter_1_cry_16 ;
    wire bfn_1_15_0_;
    wire \COUNTER.counter_1_cry_17 ;
    wire \COUNTER.counter_1_cry_18 ;
    wire \COUNTER.counter_1_cry_19 ;
    wire \COUNTER.counter_1_cry_20 ;
    wire \COUNTER.counter_1_cry_21 ;
    wire \COUNTER.counter_1_cry_22 ;
    wire \COUNTER.counter_1_cry_23 ;
    wire \COUNTER.counter_1_cry_24 ;
    wire bfn_1_16_0_;
    wire \COUNTER.counter_1_cry_25 ;
    wire \COUNTER.counter_1_cry_26 ;
    wire \COUNTER.counter_1_cry_27 ;
    wire \COUNTER.counter_1_cry_28 ;
    wire \COUNTER.counter_1_cry_29 ;
    wire \COUNTER.counter_1_cry_30 ;
    wire \PCH_PWRGD.count_rst_13_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_1 ;
    wire \PCH_PWRGD.un2_count_1_axb_1_cascade_ ;
    wire \PCH_PWRGD.count_RNI6HKKGZ0Z_1_cascade_ ;
    wire \PCH_PWRGD.count_0_0 ;
    wire \PCH_PWRGD.countZ0Z_0 ;
    wire \PCH_PWRGD.countZ0Z_0_cascade_ ;
    wire \PCH_PWRGD.N_2093_i ;
    wire \PCH_PWRGD.N_2093_i_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_13 ;
    wire \PCH_PWRGD.count_0_1 ;
    wire \PCH_PWRGD.count_rst_13 ;
    wire \PCH_PWRGD.count_1_i_a2_3_0 ;
    wire \PCH_PWRGD.count_1_i_a2_6_0 ;
    wire \PCH_PWRGD.count_1_i_a2_4_0_cascade_ ;
    wire \PCH_PWRGD.count_1_i_a2_12_0 ;
    wire \PCH_PWRGD.count_rst_0 ;
    wire \PCH_PWRGD.count_0_14 ;
    wire \PCH_PWRGD.count_1_i_a2_5_0 ;
    wire \PCH_PWRGD.un2_count_1_axb_11_cascade_ ;
    wire \PCH_PWRGD.count_0_11 ;
    wire \PCH_PWRGD.un2_count_1_axb_11 ;
    wire \PCH_PWRGD.un2_count_1_cry_10_THRU_CO ;
    wire \PCH_PWRGD.count_rst_3 ;
    wire \PCH_PWRGD.un2_count_1_cry_4_THRU_CO ;
    wire \PCH_PWRGD.count_rst_9_cascade_ ;
    wire \PCH_PWRGD.count_0_5 ;
    wire \PCH_PWRGD.count_rst_5_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_9 ;
    wire \PCH_PWRGD.un2_count_1_cry_8_THRU_CO ;
    wire \PCH_PWRGD.countZ0Z_9_cascade_ ;
    wire \PCH_PWRGD.count_0_9 ;
    wire \PCH_PWRGD.count_0_2 ;
    wire \PCH_PWRGD.count_rst_12 ;
    wire \PCH_PWRGD.count_0_10 ;
    wire \PCH_PWRGD.curr_state_RNISDK72Z0Z_0_cascade_ ;
    wire \PCH_PWRGD.count_rst_4 ;
    wire \PCH_PWRGD.countZ0Z_10 ;
    wire \PCH_PWRGD.countZ0Z_2 ;
    wire \PCH_PWRGD.countZ0Z_6 ;
    wire \PCH_PWRGD.countZ0Z_10_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_12 ;
    wire \PCH_PWRGD.countZ0Z_5 ;
    wire \PCH_PWRGD.countZ0Z_3 ;
    wire \PCH_PWRGD.count_1_i_a2_8_0_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_4 ;
    wire \PCH_PWRGD.count_1_i_a2_11_0 ;
    wire \PCH_PWRGD.count_rst_2 ;
    wire \PCH_PWRGD.count_0_12 ;
    wire \PCH_PWRGD.curr_state_0_0 ;
    wire \PCH_PWRGD.curr_state_7_0_cascade_ ;
    wire \PCH_PWRGD.curr_stateZ0Z_0_cascade_ ;
    wire \PCH_PWRGD.N_540 ;
    wire \PCH_PWRGD.N_205 ;
    wire \PCH_PWRGD.curr_state_0_1 ;
    wire \PCH_PWRGD.N_205_cascade_ ;
    wire \PCH_PWRGD.curr_stateZ0Z_1 ;
    wire \PCH_PWRGD.curr_stateZ0Z_1_cascade_ ;
    wire \PCH_PWRGD.N_2110_i_cascade_ ;
    wire \PCH_PWRGD.N_562 ;
    wire \PCH_PWRGD.N_562_cascade_ ;
    wire \PCH_PWRGD.N_38_f0_cascade_ ;
    wire \PCH_PWRGD.delayed_vccin_okZ0 ;
    wire gpio_fpga_soc_1;
    wire \HDA_STRAP.m14_i_0_cascade_ ;
    wire \HDA_STRAP.countZ0Z_13 ;
    wire \HDA_STRAP.countZ0Z_9 ;
    wire \HDA_STRAP.countZ0Z_12 ;
    wire \HDA_STRAP.countZ0Z_7 ;
    wire \HDA_STRAP.un4_count_11 ;
    wire \HDA_STRAP.countZ0Z_14 ;
    wire \HDA_STRAP.countZ0Z_15 ;
    wire \HDA_STRAP.un4_count_12 ;
    wire \HDA_STRAP.un1_count_1_cry_5_THRU_CO ;
    wire \HDA_STRAP.countZ0Z_6 ;
    wire \HDA_STRAP.un1_count_1_cry_7_THRU_CO ;
    wire \HDA_STRAP.countZ0Z_8 ;
    wire \HDA_STRAP.curr_state_RNIH91A_0Z0Z_0 ;
    wire \HDA_STRAP.N_9_cascade_ ;
    wire \HDA_STRAP.N_336 ;
    wire \HDA_STRAP.curr_stateZ0Z_2 ;
    wire hda_sdo_atp;
    wire \HDA_STRAP.un4_count ;
    wire \HDA_STRAP.curr_stateZ0Z_0 ;
    wire \HDA_STRAP.curr_stateZ0Z_1 ;
    wire vr_ready_vccin;
    wire \POWERLED.un1_dutycycle_168_0_0_o3_4_cascade_ ;
    wire \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ;
    wire \POWERLED.count_clk_0_3 ;
    wire \POWERLED.count_clkZ0Z_3 ;
    wire \POWERLED.count_clkZ0Z_3_cascade_ ;
    wire \POWERLED.count_clkZ0Z_4 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_i_i_a2_5_0_cascade_ ;
    wire \POWERLED.N_515_cascade_ ;
    wire \POWERLED.N_515 ;
    wire \POWERLED.N_47_i_cascade_ ;
    wire \POWERLED.count_clk_RNI_0Z0Z_0_cascade_ ;
    wire \POWERLED.count_clkZ0Z_0_cascade_ ;
    wire \POWERLED.count_clk_0_0 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_i_i_0 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_i_i_1 ;
    wire \POWERLED.N_415 ;
    wire \POWERLED.count_clkZ0Z_9 ;
    wire \POWERLED.count_clkZ0Z_9_cascade_ ;
    wire \POWERLED.N_320 ;
    wire \POWERLED.count_clkZ0Z_5 ;
    wire \POWERLED.N_289 ;
    wire \POWERLED.count_clkZ0Z_5_cascade_ ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_i_i_a2_1_2 ;
    wire \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ;
    wire \POWERLED.count_clk_0_5 ;
    wire \POWERLED.N_47_i ;
    wire \POWERLED.count_clkZ0Z_0 ;
    wire \POWERLED.count_clk_0_1 ;
    wire \POWERLED.count_clk_RNIZ0Z_0_cascade_ ;
    wire \POWERLED.count_clkZ0Z_1 ;
    wire \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ;
    wire \POWERLED.count_clk_0_9 ;
    wire \POWERLED.count_clkZ0Z_6 ;
    wire \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ;
    wire \POWERLED.count_clk_0_6 ;
    wire \POWERLED.count_clkZ0Z_8 ;
    wire \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ;
    wire \POWERLED.count_clk_0_8 ;
    wire \POWERLED.count_clkZ0Z_2 ;
    wire \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ;
    wire \POWERLED.count_clk_0_2 ;
    wire \POWERLED.count_clkZ0Z_7 ;
    wire \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ;
    wire \POWERLED.count_clk_0_7 ;
    wire vpp_ok;
    wire vddq_en;
    wire \COUNTER.counterZ0Z_8 ;
    wire \COUNTER.counterZ0Z_11 ;
    wire \COUNTER.counterZ0Z_10 ;
    wire \COUNTER.counterZ0Z_9 ;
    wire \COUNTER.counterZ0Z_14 ;
    wire \COUNTER.counterZ0Z_13 ;
    wire \COUNTER.counterZ0Z_15 ;
    wire \COUNTER.counterZ0Z_12 ;
    wire \COUNTER.counterZ0Z_18 ;
    wire \COUNTER.counterZ0Z_17 ;
    wire \COUNTER.counterZ0Z_19 ;
    wire \COUNTER.counterZ0Z_16 ;
    wire v33dsw_ok;
    wire \DSW_PWRGD.curr_stateZ0Z_0 ;
    wire \DSW_PWRGD.curr_stateZ0Z_1 ;
    wire DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_;
    wire G_28_cascade_;
    wire \DSW_PWRGD.un4_count_11 ;
    wire \DSW_PWRGD.un4_count_10 ;
    wire \DSW_PWRGD.un4_count_9_cascade_ ;
    wire \DSW_PWRGD.un4_count_8 ;
    wire \DSW_PWRGD.N_1_i ;
    wire \COUNTER.counterZ0Z_22 ;
    wire \COUNTER.counterZ0Z_20 ;
    wire \COUNTER.counterZ0Z_23 ;
    wire \COUNTER.counterZ0Z_21 ;
    wire \COUNTER.counterZ0Z_28 ;
    wire \COUNTER.counterZ0Z_30 ;
    wire \COUNTER.counterZ0Z_29 ;
    wire \COUNTER.counterZ0Z_31 ;
    wire \COUNTER.counterZ0Z_25 ;
    wire \COUNTER.counterZ0Z_24 ;
    wire \COUNTER.counterZ0Z_26 ;
    wire \COUNTER.counterZ0Z_27 ;
    wire \POWERLED.g0_i_o3_0_cascade_ ;
    wire \POWERLED.pwm_outZ0 ;
    wire \POWERLED.g0_i_o3_0 ;
    wire pwrbtn_led;
    wire \POWERLED.curr_state_3_0_cascade_ ;
    wire \POWERLED.curr_stateZ0Z_0_cascade_ ;
    wire \POWERLED.count_0_sqmuxa_i_cascade_ ;
    wire \POWERLED.count_RNIZ0Z_0_cascade_ ;
    wire \POWERLED.count_RNIZ0Z_1_cascade_ ;
    wire \POWERLED.countZ0Z_1_cascade_ ;
    wire \POWERLED.count_0_1 ;
    wire \POWERLED.count_0_0 ;
    wire \POWERLED.count_0_3 ;
    wire \POWERLED.count_0_12 ;
    wire \PCH_PWRGD.countZ0Z_15 ;
    wire \PCH_PWRGD.count_rst ;
    wire \PCH_PWRGD.count_0_15 ;
    wire \PCH_PWRGD.N_2110_i ;
    wire \PCH_PWRGD.N_314 ;
    wire \PCH_PWRGD.curr_stateZ0Z_0 ;
    wire \PCH_PWRGD.N_2091_i ;
    wire \POWERLED.count_0_13 ;
    wire \POWERLED.count_0_4 ;
    wire \POWERLED.count_0_5 ;
    wire bfn_4_5_0_;
    wire \POWERLED.mult1_un138_sum_cry_2 ;
    wire \POWERLED.mult1_un138_sum_cry_3 ;
    wire \POWERLED.mult1_un138_sum_cry_4 ;
    wire \POWERLED.mult1_un138_sum_cry_5 ;
    wire \POWERLED.mult1_un138_sum_cry_6 ;
    wire \POWERLED.mult1_un138_sum_cry_7 ;
    wire bfn_4_6_0_;
    wire \POWERLED.mult1_un131_sum_cry_3_s ;
    wire \POWERLED.mult1_un131_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_cry_4_s ;
    wire \POWERLED.mult1_un131_sum_cry_3 ;
    wire \POWERLED.mult1_un131_sum_cry_5_s ;
    wire \POWERLED.mult1_un131_sum_cry_4 ;
    wire \POWERLED.mult1_un131_sum_cry_6_s ;
    wire \POWERLED.mult1_un131_sum_cry_5 ;
    wire \POWERLED.mult1_un124_sum_i_0_8 ;
    wire \POWERLED.mult1_un138_sum_axb_8 ;
    wire \POWERLED.mult1_un131_sum_cry_6 ;
    wire \POWERLED.mult1_un131_sum_cry_7 ;
    wire \POWERLED.mult1_un131_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un131_sum_i_0_8 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a3_0_0_cascade_ ;
    wire \POWERLED.N_96_cascade_ ;
    wire \POWERLED.count_off_0_4 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a3_1 ;
    wire \POWERLED.N_455_cascade_ ;
    wire \POWERLED.count_clk_en_0_cascade_ ;
    wire \POWERLED.func_state_RNI81TV4Z0Z_1 ;
    wire \POWERLED.N_480 ;
    wire \POWERLED.func_state_1_ss0_i_0_o3_1_cascade_ ;
    wire \POWERLED.N_217 ;
    wire \POWERLED.N_217_cascade_ ;
    wire \POWERLED.N_321_cascade_ ;
    wire \POWERLED.func_state_1_ss0_i_0_o3_0 ;
    wire vccst_en;
    wire \POWERLED.N_516 ;
    wire \POWERLED.N_516_cascade_ ;
    wire \POWERLED.N_403 ;
    wire bfn_4_12_0_;
    wire \COUNTER.un4_counter_0 ;
    wire \COUNTER.un4_counter_2_and ;
    wire \COUNTER.un4_counter_1 ;
    wire \COUNTER.un4_counter_3_and ;
    wire \COUNTER.un4_counter_2 ;
    wire \COUNTER.un4_counter_4_and ;
    wire \COUNTER.un4_counter_3 ;
    wire \COUNTER.un4_counter_5_and ;
    wire \COUNTER.un4_counter_4 ;
    wire \COUNTER.un4_counter_6_and ;
    wire \COUNTER.un4_counter_5 ;
    wire \COUNTER.un4_counter_7_and ;
    wire \COUNTER.un4_counter_6 ;
    wire COUNTER_un4_counter_7;
    wire bfn_4_13_0_;
    wire \COUNTER.counter_1_cry_4_THRU_CO ;
    wire \COUNTER.counter_1_cry_2_THRU_CO ;
    wire \COUNTER.counterZ0Z_3 ;
    wire \COUNTER.un4_counter_0_and ;
    wire \COUNTER.counterZ0Z_1 ;
    wire \COUNTER.counterZ0Z_5 ;
    wire \COUNTER.counterZ0Z_7 ;
    wire \COUNTER.un4_counter_1_and ;
    wire \COUNTER.counter_1_cry_3_THRU_CO ;
    wire \COUNTER.counterZ0Z_4 ;
    wire \COUNTER.counter_1_cry_5_THRU_CO ;
    wire \COUNTER.counterZ0Z_6 ;
    wire \DSW_PWRGD.un1_curr_state10_0 ;
    wire \DSW_PWRGD.countZ0Z_0 ;
    wire bfn_4_14_0_;
    wire \DSW_PWRGD.countZ0Z_1 ;
    wire \DSW_PWRGD.un1_count_1_cry_0 ;
    wire \DSW_PWRGD.countZ0Z_2 ;
    wire \DSW_PWRGD.un1_count_1_cry_1 ;
    wire \DSW_PWRGD.countZ0Z_3 ;
    wire \DSW_PWRGD.un1_count_1_cry_2 ;
    wire \DSW_PWRGD.countZ0Z_4 ;
    wire \DSW_PWRGD.un1_count_1_cry_3 ;
    wire \DSW_PWRGD.countZ0Z_5 ;
    wire \DSW_PWRGD.un1_count_1_cry_4 ;
    wire \DSW_PWRGD.countZ0Z_6 ;
    wire \DSW_PWRGD.un1_count_1_cry_5 ;
    wire \DSW_PWRGD.countZ0Z_7 ;
    wire \DSW_PWRGD.un1_count_1_cry_6 ;
    wire \DSW_PWRGD.un1_count_1_cry_7 ;
    wire \DSW_PWRGD.countZ0Z_8 ;
    wire bfn_4_15_0_;
    wire \DSW_PWRGD.countZ0Z_9 ;
    wire \DSW_PWRGD.un1_count_1_cry_8 ;
    wire \DSW_PWRGD.countZ0Z_10 ;
    wire \DSW_PWRGD.un1_count_1_cry_9 ;
    wire \DSW_PWRGD.countZ0Z_11 ;
    wire \DSW_PWRGD.un1_count_1_cry_10 ;
    wire \DSW_PWRGD.countZ0Z_12 ;
    wire \DSW_PWRGD.un1_count_1_cry_11 ;
    wire \DSW_PWRGD.countZ0Z_13 ;
    wire \DSW_PWRGD.un1_count_1_cry_12 ;
    wire \DSW_PWRGD.countZ0Z_14 ;
    wire \DSW_PWRGD.un1_count_1_cry_13 ;
    wire \DSW_PWRGD.un1_count_1_cry_14 ;
    wire \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_4_16_0_;
    wire \DSW_PWRGD.countZ0Z_15 ;
    wire \DSW_PWRGD.N_42_1 ;
    wire G_28;
    wire \POWERLED.un79_clk_100khzlt6_cascade_ ;
    wire \POWERLED.un79_clk_100khzlto15_5_cascade_ ;
    wire \POWERLED.un79_clk_100khzlto15_7_cascade_ ;
    wire \POWERLED.un79_clk_100khzlto15_3 ;
    wire \POWERLED.count_RNIZ0Z_8_cascade_ ;
    wire \POWERLED.pwm_out_1_sqmuxa ;
    wire \POWERLED.N_8 ;
    wire bfn_5_2_0_;
    wire \POWERLED.un1_count_cry_1 ;
    wire \POWERLED.un1_count_cry_2_c_RNICZ0Z419 ;
    wire \POWERLED.un1_count_cry_2 ;
    wire \POWERLED.un1_count_cry_3_c_RNIDZ0Z629 ;
    wire \POWERLED.un1_count_cry_3 ;
    wire \POWERLED.un1_count_cry_4_c_RNIEZ0Z839 ;
    wire \POWERLED.un1_count_cry_4 ;
    wire \POWERLED.un1_count_cry_5 ;
    wire \POWERLED.un1_count_cry_6 ;
    wire \POWERLED.un1_count_cry_7 ;
    wire \POWERLED.un1_count_cry_8 ;
    wire bfn_5_3_0_;
    wire \POWERLED.un1_count_cry_9 ;
    wire \POWERLED.un1_count_cry_10 ;
    wire \POWERLED.un1_count_cry_11_c_RNISEHZ0Z7 ;
    wire \POWERLED.un1_count_cry_11 ;
    wire \POWERLED.un1_count_cry_12_c_RNITGIZ0Z7 ;
    wire \POWERLED.un1_count_cry_12 ;
    wire \POWERLED.un1_count_cry_13 ;
    wire \POWERLED.count_0_sqmuxa_i ;
    wire \POWERLED.un1_count_cry_14 ;
    wire \POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7 ;
    wire \POWERLED.count_0_14 ;
    wire \POWERLED.mult1_un131_sum_s_8 ;
    wire vccst_pwrgd;
    wire bfn_5_5_0_;
    wire \POWERLED.mult1_un145_sum_cry_2 ;
    wire \POWERLED.mult1_un138_sum_cry_3_s ;
    wire \POWERLED.mult1_un145_sum_cry_3 ;
    wire \POWERLED.mult1_un138_sum_cry_4_s ;
    wire \POWERLED.mult1_un145_sum_cry_4 ;
    wire \POWERLED.mult1_un138_sum_cry_5_s ;
    wire \POWERLED.mult1_un145_sum_cry_5 ;
    wire \POWERLED.mult1_un138_sum_cry_6_s ;
    wire \POWERLED.mult1_un145_sum_cry_6 ;
    wire \POWERLED.mult1_un145_sum_axb_8 ;
    wire \POWERLED.mult1_un145_sum_cry_7 ;
    wire \POWERLED.mult1_un138_sum_s_8 ;
    wire \POWERLED.mult1_un138_sum_i_0_8 ;
    wire bfn_5_6_0_;
    wire \POWERLED.mult1_un124_sum_cry_3_s ;
    wire \POWERLED.mult1_un124_sum_cry_2 ;
    wire \POWERLED.mult1_un124_sum_cry_4_s ;
    wire \POWERLED.mult1_un124_sum_cry_3 ;
    wire \POWERLED.mult1_un124_sum_cry_5_s ;
    wire \POWERLED.mult1_un124_sum_cry_4 ;
    wire \POWERLED.mult1_un124_sum_cry_6_s ;
    wire \POWERLED.mult1_un124_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_axb_8 ;
    wire \POWERLED.mult1_un124_sum_cry_6 ;
    wire \POWERLED.mult1_un124_sum_cry_7 ;
    wire \POWERLED.mult1_un124_sum_s_8 ;
    wire \POWERLED.mult1_un124_sum_axb_7_l_fx ;
    wire bfn_5_8_0_;
    wire \POWERLED.mult1_un159_sum_cry_1 ;
    wire \POWERLED.mult1_un159_sum_cry_2 ;
    wire \POWERLED.mult1_un159_sum_cry_3 ;
    wire \POWERLED.mult1_un159_sum_cry_4 ;
    wire \POWERLED.mult1_un159_sum_cry_5 ;
    wire \POWERLED.mult1_un159_sum_cry_6 ;
    wire \POWERLED.mult1_un152_sum_i_0_8 ;
    wire bfn_5_9_0_;
    wire \POWERLED.mult1_un145_sum_i ;
    wire \POWERLED.mult1_un152_sum_cry_3_s ;
    wire \POWERLED.mult1_un152_sum_cry_2 ;
    wire \POWERLED.mult1_un145_sum_cry_3_s ;
    wire \POWERLED.mult1_un152_sum_cry_4_s ;
    wire \POWERLED.mult1_un152_sum_cry_3 ;
    wire \POWERLED.mult1_un145_sum_cry_4_s ;
    wire \POWERLED.mult1_un152_sum_cry_5_s ;
    wire \POWERLED.mult1_un152_sum_cry_4 ;
    wire \POWERLED.mult1_un145_sum_cry_5_s ;
    wire \POWERLED.mult1_un152_sum_cry_6_s ;
    wire \POWERLED.mult1_un152_sum_cry_5 ;
    wire \POWERLED.mult1_un145_sum_cry_6_s ;
    wire \POWERLED.mult1_un159_sum_axb_7 ;
    wire \POWERLED.mult1_un152_sum_cry_6 ;
    wire \POWERLED.mult1_un152_sum_axb_8 ;
    wire \POWERLED.mult1_un152_sum_cry_7 ;
    wire \POWERLED.mult1_un152_sum_s_8 ;
    wire \POWERLED.mult1_un145_sum_s_8 ;
    wire \POWERLED.mult1_un145_sum_i_0_8 ;
    wire \POWERLED.count_clk_RNIZ0Z_9 ;
    wire \POWERLED.un1_func_state25_6_0_o_N_423_N_cascade_ ;
    wire \POWERLED.N_348 ;
    wire \POWERLED.func_state_1_m0_0_0_0 ;
    wire \POWERLED.func_state_RNI5DLR_0Z0Z_0_cascade_ ;
    wire \POWERLED.func_state_1_m0_0_cascade_ ;
    wire \POWERLED.count_clk_RNIZ0Z_7 ;
    wire \POWERLED.un34_clk_100khz_11_cascade_ ;
    wire \POWERLED.un34_clk_100khz_8 ;
    wire \POWERLED.N_322 ;
    wire \POWERLED.un34_clk_100khz_9 ;
    wire \POWERLED.count_off_0_3 ;
    wire \POWERLED.count_off_1_0 ;
    wire \POWERLED.count_offZ0Z_0_cascade_ ;
    wire \POWERLED.count_off_0_0 ;
    wire \COUNTER.counterZ0Z_0 ;
    wire \POWERLED.count_off_RNIZ0Z_1 ;
    wire \POWERLED.count_off_0_1 ;
    wire \POWERLED.count_off_RNIZ0Z_1_cascade_ ;
    wire \POWERLED.un34_clk_100khz_10 ;
    wire \COUNTER.counter_1_cry_1_THRU_CO ;
    wire \COUNTER.counterZ0Z_2 ;
    wire \POWERLED.count_off_0_13 ;
    wire \POWERLED.count_off_0_5 ;
    wire \POWERLED.count_off_0_14 ;
    wire \POWERLED.count_off_0_6 ;
    wire \POWERLED.un1_count_cry_5_c_RNIFAZ0Z49 ;
    wire \POWERLED.count_0_6 ;
    wire \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ;
    wire \POWERLED.count_0_15 ;
    wire \POWERLED.un1_count_cry_6_c_RNIGCZ0Z59 ;
    wire \POWERLED.count_0_7 ;
    wire \POWERLED.un1_count_cry_7_c_RNIHEZ0Z69 ;
    wire \POWERLED.count_0_8 ;
    wire \POWERLED.un1_count_cry_8_c_RNIIGZ0Z79 ;
    wire \POWERLED.count_0_9 ;
    wire \POWERLED.un1_count_cry_9_c_RNIJIZ0Z89 ;
    wire \POWERLED.count_0_10 ;
    wire \POWERLED.un1_count_cry_1_c_RNIBZ0Z209 ;
    wire \POWERLED.count_0_2 ;
    wire \POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7 ;
    wire \POWERLED.count_0_11 ;
    wire \POWERLED.countZ0Z_0 ;
    wire \POWERLED.un1_count_cry_0_i ;
    wire bfn_6_3_0_;
    wire \POWERLED.countZ0Z_1 ;
    wire \POWERLED.N_4698_i ;
    wire \POWERLED.un85_clk_100khz_cry_0 ;
    wire \POWERLED.un85_clk_100khz_2 ;
    wire \POWERLED.countZ0Z_2 ;
    wire \POWERLED.N_4699_i ;
    wire \POWERLED.un85_clk_100khz_cry_1 ;
    wire \POWERLED.countZ0Z_3 ;
    wire \POWERLED.un85_clk_100khz_3 ;
    wire \POWERLED.N_4700_i ;
    wire \POWERLED.un85_clk_100khz_cry_2 ;
    wire \POWERLED.countZ0Z_4 ;
    wire \POWERLED.un85_clk_100khz_4 ;
    wire \POWERLED.N_4701_i ;
    wire \POWERLED.un85_clk_100khz_cry_3 ;
    wire \POWERLED.un85_clk_100khz_5 ;
    wire \POWERLED.countZ0Z_5 ;
    wire \POWERLED.N_4702_i ;
    wire \POWERLED.un85_clk_100khz_cry_4 ;
    wire \POWERLED.un85_clk_100khz_6 ;
    wire \POWERLED.countZ0Z_6 ;
    wire \POWERLED.N_4703_i ;
    wire \POWERLED.un85_clk_100khz_cry_5 ;
    wire \POWERLED.countZ0Z_7 ;
    wire \POWERLED.N_4704_i ;
    wire \POWERLED.un85_clk_100khz_cry_6 ;
    wire \POWERLED.un85_clk_100khz_cry_7 ;
    wire \POWERLED.countZ0Z_8 ;
    wire \POWERLED.N_4705_i ;
    wire bfn_6_4_0_;
    wire \POWERLED.countZ0Z_9 ;
    wire \POWERLED.N_4706_i ;
    wire \POWERLED.un85_clk_100khz_cry_8 ;
    wire \POWERLED.countZ0Z_10 ;
    wire \POWERLED.N_4707_i ;
    wire \POWERLED.un85_clk_100khz_cry_9 ;
    wire \POWERLED.countZ0Z_11 ;
    wire \POWERLED.N_4708_i ;
    wire \POWERLED.un85_clk_100khz_cry_10 ;
    wire \POWERLED.countZ0Z_12 ;
    wire \POWERLED.N_4709_i ;
    wire \POWERLED.un85_clk_100khz_cry_11 ;
    wire \POWERLED.countZ0Z_13 ;
    wire \POWERLED.N_4710_i ;
    wire \POWERLED.un85_clk_100khz_cry_12 ;
    wire \POWERLED.countZ0Z_14 ;
    wire \POWERLED.N_4711_i ;
    wire \POWERLED.un85_clk_100khz_cry_13 ;
    wire \POWERLED.countZ0Z_15 ;
    wire \POWERLED.N_4712_i ;
    wire \POWERLED.un85_clk_100khz_cry_14 ;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0 ;
    wire bfn_6_5_0_;
    wire \POWERLED.un85_clk_100khz_7 ;
    wire \POWERLED.mult1_un131_sum_i ;
    wire \POWERLED.mult1_un138_sum_i ;
    wire \POWERLED.mult1_un117_sum_i ;
    wire \POWERLED.mult1_un124_sum_i ;
    wire bfn_6_6_0_;
    wire \POWERLED.mult1_un110_sum_i ;
    wire \POWERLED.mult1_un117_sum_cry_2 ;
    wire \POWERLED.mult1_un117_sum_cry_4_s ;
    wire \POWERLED.mult1_un117_sum_cry_3 ;
    wire \POWERLED.mult1_un117_sum_cry_5_s ;
    wire \POWERLED.mult1_un117_sum_cry_4 ;
    wire \POWERLED.mult1_un117_sum_cry_6_s ;
    wire \POWERLED.mult1_un117_sum_cry_5 ;
    wire \POWERLED.mult1_un110_sum_i_0_8 ;
    wire \POWERLED.mult1_un124_sum_axb_8 ;
    wire \POWERLED.mult1_un117_sum_cry_6 ;
    wire \POWERLED.mult1_un117_sum_cry_7 ;
    wire \POWERLED.mult1_un117_sum_cry_3_s ;
    wire \POWERLED.mult1_un117_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un124_sum_axb_4_l_fx ;
    wire \PCH_PWRGD.N_38_f0 ;
    wire \PCH_PWRGD.curr_state_0_sqmuxa ;
    wire \PCH_PWRGD.delayed_vccin_ok_0 ;
    wire \POWERLED.mult1_un117_sum_s_8 ;
    wire \POWERLED.mult1_un117_sum_i_0_8 ;
    wire \POWERLED.N_341_cascade_ ;
    wire bfn_6_8_0_;
    wire \POWERLED.mult1_un166_sum_cry_0 ;
    wire \POWERLED.mult1_un159_sum_cry_2_s ;
    wire \POWERLED.mult1_un166_sum_cry_1 ;
    wire \POWERLED.mult1_un159_sum_cry_3_s ;
    wire \POWERLED.mult1_un166_sum_cry_2 ;
    wire \POWERLED.mult1_un159_sum_cry_4_s ;
    wire \POWERLED.mult1_un166_sum_cry_3 ;
    wire \POWERLED.mult1_un159_sum_cry_5_s ;
    wire G_2129;
    wire \POWERLED.mult1_un166_sum_cry_4 ;
    wire \POWERLED.mult1_un166_sum_axb_6 ;
    wire \POWERLED.mult1_un166_sum_cry_5 ;
    wire \POWERLED.un85_clk_100khz_0 ;
    wire \POWERLED.mult1_un159_sum_s_7 ;
    wire \POWERLED.un85_clk_100khz_1 ;
    wire \POWERLED.N_394_cascade_ ;
    wire \POWERLED.N_453 ;
    wire \POWERLED.func_state_RNI5DLR_1Z0Z_1 ;
    wire \POWERLED.un1_func_state25_6_0_0_a3_0_cascade_ ;
    wire \POWERLED.un1_func_state25_6_0_o_N_422_N ;
    wire \POWERLED.un1_func_state25_6_0_o_N_516_N ;
    wire \POWERLED.un1_func_state25_6_0_o_N_425_N ;
    wire \POWERLED.un1_func_state25_6_0_0_2 ;
    wire \POWERLED.un1_func_state25_6_0_0_0 ;
    wire m3_1;
    wire \POWERLED.count_off_RNI_0Z0Z_10 ;
    wire \POWERLED.func_state_RNI5DLR_0Z0Z_0 ;
    wire \POWERLED.func_state_1_m0_i_o2_2_1 ;
    wire \POWERLED.func_state_RNILFRF4Z0Z_0 ;
    wire \POWERLED.N_143_cascade_ ;
    wire \POWERLED.func_stateZ1Z_0 ;
    wire \POWERLED.func_state_RNIU8CJBZ0Z_0 ;
    wire \POWERLED.func_stateZ0Z_0_cascade_ ;
    wire \POWERLED.count_off_0_10 ;
    wire \POWERLED.count_off_0_11 ;
    wire \POWERLED.count_off_0_2 ;
    wire \POWERLED.count_off_0_12 ;
    wire \POWERLED.count_offZ0Z_0 ;
    wire \POWERLED.count_offZ0Z_1 ;
    wire bfn_6_12_0_;
    wire \POWERLED.count_offZ0Z_2 ;
    wire \POWERLED.count_off_1_2 ;
    wire \POWERLED.un3_count_off_1_cry_1 ;
    wire \POWERLED.count_offZ0Z_3 ;
    wire \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ;
    wire \POWERLED.un3_count_off_1_cry_2 ;
    wire \POWERLED.count_offZ0Z_4 ;
    wire \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ;
    wire \POWERLED.un3_count_off_1_cry_3 ;
    wire \POWERLED.count_offZ0Z_5 ;
    wire \POWERLED.count_off_1_5 ;
    wire \POWERLED.un3_count_off_1_cry_4 ;
    wire \POWERLED.count_offZ0Z_6 ;
    wire \POWERLED.count_off_1_6 ;
    wire \POWERLED.un3_count_off_1_cry_5 ;
    wire \POWERLED.un3_count_off_1_cry_6 ;
    wire \POWERLED.un3_count_off_1_cry_7 ;
    wire \POWERLED.un3_count_off_1_cry_8 ;
    wire bfn_6_13_0_;
    wire \POWERLED.count_offZ0Z_10 ;
    wire \POWERLED.count_off_1_10 ;
    wire \POWERLED.un3_count_off_1_cry_9 ;
    wire \POWERLED.count_offZ0Z_11 ;
    wire \POWERLED.count_off_1_11 ;
    wire \POWERLED.un3_count_off_1_cry_10 ;
    wire \POWERLED.count_offZ0Z_12 ;
    wire \POWERLED.count_off_1_12 ;
    wire \POWERLED.un3_count_off_1_cry_11 ;
    wire \POWERLED.count_offZ0Z_13 ;
    wire \POWERLED.count_off_1_13 ;
    wire \POWERLED.un3_count_off_1_cry_12 ;
    wire \POWERLED.count_offZ0Z_14 ;
    wire \POWERLED.count_off_1_14 ;
    wire \POWERLED.un3_count_off_1_cry_13 ;
    wire \POWERLED.N_96 ;
    wire \POWERLED.un3_count_off_1_cry_14 ;
    wire \POWERLED.count_offZ0Z_9 ;
    wire \POWERLED.count_offZ0Z_15 ;
    wire \POWERLED.un3_count_off_1_cry_14_c_RNIMONZ0Z33 ;
    wire \POWERLED.count_off_0_15 ;
    wire \POWERLED.count_offZ0Z_7 ;
    wire \POWERLED.count_off_1_7 ;
    wire \POWERLED.count_off_0_7 ;
    wire \POWERLED.count_offZ0Z_8 ;
    wire \POWERLED.count_off_1_8 ;
    wire \POWERLED.count_off_0_8 ;
    wire \POWERLED.count_off_1_9 ;
    wire \POWERLED.count_off_0_9 ;
    wire \POWERLED.count_off_enZ0 ;
    wire G_10;
    wire \POWERLED.un85_clk_100khz_11 ;
    wire \POWERLED.un85_clk_100khz_10 ;
    wire \PCH_PWRGD.count_rst_8 ;
    wire \PCH_PWRGD.count_0_6 ;
    wire \PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ;
    wire \PCH_PWRGD.count_0_sqmuxa ;
    wire N_355;
    wire pch_pwrok;
    wire \POWERLED.mult1_un68_sum_i_8 ;
    wire \POWERLED.mult1_un75_sum_i_8 ;
    wire \POWERLED.un85_clk_100khz_9 ;
    wire \POWERLED.un85_clk_100khz_8 ;
    wire bfn_7_4_0_;
    wire \POWERLED.mult1_un103_sum_i ;
    wire \POWERLED.mult1_un110_sum_cry_3_s ;
    wire \POWERLED.mult1_un110_sum_cry_2 ;
    wire \POWERLED.mult1_un110_sum_cry_4_s ;
    wire \POWERLED.mult1_un110_sum_cry_3 ;
    wire \POWERLED.mult1_un110_sum_cry_5_s ;
    wire \POWERLED.mult1_un110_sum_cry_4 ;
    wire \POWERLED.mult1_un110_sum_cry_6_s ;
    wire \POWERLED.mult1_un110_sum_cry_5 ;
    wire \POWERLED.mult1_un103_sum_i_0_8 ;
    wire \POWERLED.mult1_un117_sum_axb_8 ;
    wire \POWERLED.mult1_un110_sum_cry_6 ;
    wire \POWERLED.mult1_un110_sum_cry_7 ;
    wire \POWERLED.mult1_un110_sum_s_8 ;
    wire \POWERLED.un85_clk_100khz_12 ;
    wire \POWERLED.mult1_un145_sum ;
    wire bfn_7_5_0_;
    wire \POWERLED.mult1_un138_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_0_cZ0 ;
    wire \POWERLED.mult1_un131_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_1_cZ0 ;
    wire \POWERLED.mult1_un124_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_2_cZ0 ;
    wire \POWERLED.mult1_un117_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_3_cZ0 ;
    wire \POWERLED.mult1_un110_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_4_cZ0 ;
    wire \POWERLED.un1_dutycycle_53_cry_5_cZ0 ;
    wire \POWERLED.un1_dutycycle_53_cry_6_cZ0 ;
    wire \POWERLED.un1_dutycycle_53_cry_7_cZ0 ;
    wire bfn_7_6_0_;
    wire \POWERLED.un1_dutycycle_53_cry_8 ;
    wire \POWERLED.un1_dutycycle_53_cry_9 ;
    wire \POWERLED.un1_dutycycle_53_cry_10 ;
    wire \POWERLED.un1_dutycycle_53_cry_11 ;
    wire \POWERLED.un1_dutycycle_53_cry_12 ;
    wire \POWERLED.un1_dutycycle_53_cry_13 ;
    wire \POWERLED.un1_dutycycle_53_cry_14 ;
    wire \POWERLED.un1_dutycycle_53_cry_15 ;
    wire bfn_7_7_0_;
    wire \POWERLED.CO2 ;
    wire \POWERLED.N_76_f0 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_1 ;
    wire \POWERLED.mult1_un159_sum_i ;
    wire \POWERLED.mult1_un152_sum_i ;
    wire \POWERLED.func_state_1_m0_i_o2_0_1 ;
    wire N_21;
    wire func_state_RNITGMHB_0_1_cascade_;
    wire \POWERLED.dutycycle_RNIZ0Z_3 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_1 ;
    wire \POWERLED.dutycycle_RNIZ0Z_2 ;
    wire \POWERLED.func_state_RNICK8N9Z0Z_1 ;
    wire \POWERLED.func_stateZ0Z_1 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_3 ;
    wire \POWERLED.N_80_f0_cascade_ ;
    wire \POWERLED.dutycycle_RNI375F3Z0Z_7 ;
    wire \POWERLED.dutycycleZ1Z_7 ;
    wire \POWERLED.dutycycle_RNI375F3Z0Z_7_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_4_cascade_ ;
    wire \RSMRST_PWRGD.N_8_mux ;
    wire m57_i_o2_2_cascade_;
    wire \RSMRST_PWRGD.N_4713_0_0_0_cascade_ ;
    wire \POWERLED.N_569_N_cascade_ ;
    wire \POWERLED.N_220_N_cascade_ ;
    wire \POWERLED.N_282_N_cascade_ ;
    wire \POWERLED.dutycycle_eena_8_d_cascade_ ;
    wire \POWERLED.dutycycle_RNI79E14Z0Z_3_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_6_cascade_ ;
    wire \POWERLED.dutycycle_eena_8_c ;
    wire \POWERLED.dutycycle_RNI79E14Z0Z_3 ;
    wire \POWERLED.dutycycleZ0Z_3 ;
    wire \POWERLED.N_2168_i ;
    wire \POWERLED.N_231_i_cascade_ ;
    wire \POWERLED.N_321 ;
    wire \POWERLED.N_52_i_i_0 ;
    wire \POWERLED.N_410_cascade_ ;
    wire \POWERLED.func_state_RNI1J4E2Z0Z_1 ;
    wire COUNTER_un4_counter_7_THRU_CO;
    wire G_44_cascade_;
    wire N_365;
    wire \VPP_VDDQ.N_464_i ;
    wire bfn_7_14_0_;
    wire \VPP_VDDQ.un1_count_1_cry_0 ;
    wire \VPP_VDDQ.un1_count_1_cry_1 ;
    wire \VPP_VDDQ.un1_count_1_cry_2 ;
    wire \VPP_VDDQ.un1_count_1_cry_3 ;
    wire \VPP_VDDQ.un1_count_1_cry_4 ;
    wire \VPP_VDDQ.un1_count_1_cry_5 ;
    wire \VPP_VDDQ.un1_count_1_cry_6 ;
    wire \VPP_VDDQ.un1_count_1_cry_7 ;
    wire bfn_7_15_0_;
    wire \VPP_VDDQ.un1_count_1_cry_8 ;
    wire \VPP_VDDQ.un1_count_1_cry_9 ;
    wire \VPP_VDDQ.un1_count_1_cry_10 ;
    wire \VPP_VDDQ.un1_count_1_cry_11 ;
    wire \VPP_VDDQ.un1_count_1_cry_12 ;
    wire \VPP_VDDQ.un1_count_1_cry_13 ;
    wire \VPP_VDDQ.un1_count_1_cry_14 ;
    wire \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_7_16_0_;
    wire \VPP_VDDQ.N_42_0 ;
    wire G_44;
    wire \POWERLED.mult1_un89_sum ;
    wire bfn_8_1_0_;
    wire \POWERLED.mult1_un82_sum_i ;
    wire \POWERLED.mult1_un89_sum_cry_2 ;
    wire \POWERLED.mult1_un89_sum_cry_3 ;
    wire \POWERLED.mult1_un89_sum_cry_4 ;
    wire \POWERLED.mult1_un89_sum_cry_5 ;
    wire \POWERLED.mult1_un89_sum_cry_6 ;
    wire \POWERLED.mult1_un89_sum_cry_7 ;
    wire \POWERLED.mult1_un89_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un96_sum ;
    wire bfn_8_2_0_;
    wire \POWERLED.mult1_un89_sum_i ;
    wire \POWERLED.mult1_un96_sum_cry_2 ;
    wire \POWERLED.mult1_un89_sum_cry_3_s ;
    wire \POWERLED.mult1_un96_sum_cry_3 ;
    wire \POWERLED.mult1_un89_sum_cry_4_s ;
    wire \POWERLED.mult1_un96_sum_cry_4 ;
    wire \POWERLED.mult1_un89_sum_s_8 ;
    wire \POWERLED.mult1_un89_sum_cry_5_s ;
    wire \POWERLED.mult1_un96_sum_cry_5 ;
    wire \POWERLED.mult1_un89_sum_cry_6_s ;
    wire \POWERLED.mult1_un89_sum_i_0_8 ;
    wire \POWERLED.mult1_un96_sum_cry_6 ;
    wire \POWERLED.mult1_un96_sum_axb_8 ;
    wire \POWERLED.mult1_un96_sum_cry_7 ;
    wire \POWERLED.mult1_un82_sum_i_0_8 ;
    wire \POWERLED.mult1_un103_sum ;
    wire bfn_8_3_0_;
    wire \POWERLED.mult1_un96_sum_i ;
    wire \POWERLED.mult1_un103_sum_cry_3_s ;
    wire \POWERLED.mult1_un103_sum_cry_2 ;
    wire \POWERLED.mult1_un96_sum_cry_3_s ;
    wire \POWERLED.mult1_un103_sum_cry_4_s ;
    wire \POWERLED.mult1_un103_sum_cry_3 ;
    wire \POWERLED.mult1_un96_sum_cry_4_s ;
    wire \POWERLED.mult1_un103_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_cry_4 ;
    wire \POWERLED.mult1_un96_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_cry_6_s ;
    wire \POWERLED.mult1_un103_sum_cry_5 ;
    wire \POWERLED.mult1_un96_sum_cry_6_s ;
    wire \POWERLED.mult1_un110_sum_axb_8 ;
    wire \POWERLED.mult1_un103_sum_cry_6 ;
    wire \POWERLED.mult1_un103_sum_axb_8 ;
    wire \POWERLED.mult1_un103_sum_cry_7 ;
    wire \POWERLED.mult1_un103_sum_s_8 ;
    wire \POWERLED.mult1_un96_sum_s_8 ;
    wire \POWERLED.mult1_un96_sum_i_0_8 ;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ;
    wire \POWERLED.curr_stateZ0Z_0 ;
    wire \POWERLED.count_RNIZ0Z_8 ;
    wire \POWERLED.curr_state_2_0 ;
    wire \POWERLED.CO2_THRU_CO ;
    wire \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ;
    wire \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_1 ;
    wire \POWERLED.g0_1_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_3 ;
    wire \POWERLED.g0_1_1 ;
    wire \POWERLED.dutycycle_RNIZ0Z_7_cascade_ ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_7 ;
    wire \POWERLED.dutycycle_RNI_9Z0Z_7_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_11 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_13 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_12 ;
    wire \POWERLED.N_9_i_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_7 ;
    wire \POWERLED.dutycycleZ1Z_4 ;
    wire \POWERLED.dutycycle_en_6 ;
    wire \POWERLED.dutycycleZ0Z_8_cascade_ ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_4_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_axb_12_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_15 ;
    wire \POWERLED.dutycycle_RNI_8Z0Z_10 ;
    wire \POWERLED.dutycycleZ0Z_15 ;
    wire \POWERLED.dutycycleZ0Z_12_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_15 ;
    wire \POWERLED.m69_0_o2_7 ;
    wire \POWERLED.N_81_cascade_ ;
    wire \POWERLED.N_85 ;
    wire \POWERLED.dutycycleZ1Z_1 ;
    wire \POWERLED.N_85_cascade_ ;
    wire \POWERLED.dutycycle_cascade_ ;
    wire \POWERLED.dutycycle_eena_0 ;
    wire \POWERLED.dutycycle_eena ;
    wire \POWERLED.dutycycle_eena_cascade_ ;
    wire \POWERLED.N_81 ;
    wire \POWERLED.dutycycleZ1Z_0 ;
    wire \POWERLED.N_441_cascade_ ;
    wire \POWERLED.dutycycle_eena_13 ;
    wire \POWERLED.dutycycle_0_6 ;
    wire \POWERLED.dutycycle_eena_13_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_6_cascade_ ;
    wire \POWERLED.N_442 ;
    wire \POWERLED.N_429_cascade_ ;
    wire \POWERLED.dutycycle_RNI9NTJ2Z0Z_2 ;
    wire \POWERLED.dutycycle_RNI9NTJ2Z0Z_2_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_2 ;
    wire N_2145_i_cascade_;
    wire \POWERLED.dutycycle_RNI_3Z0Z_6_cascade_ ;
    wire \POWERLED.func_stateZ0Z_0 ;
    wire \RSMRST_PWRGD.N_13 ;
    wire POWERLED_dutycycle_eena_14_0;
    wire \POWERLED.dutycycle_0_5 ;
    wire POWERLED_dutycycle_eena_14_0_cascade_;
    wire dutycycle_RNIKBMSJ_0_5_cascade_;
    wire \POWERLED.func_state_RNI_0Z0Z_0 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_5_cascade_ ;
    wire \POWERLED.func_state_RNI_5Z0Z_0 ;
    wire SUSWARN_N_rep1;
    wire \POWERLED.dutycycle_eena_5_0_s_tzZ0Z_1_cascade_ ;
    wire \POWERLED.N_443 ;
    wire POWERLED_func_state_0_sqmuxa_cascade_;
    wire N_14;
    wire \VPP_VDDQ.count_2_1_4_cascade_ ;
    wire \VPP_VDDQ.count_2_0_4 ;
    wire \VPP_VDDQ.count_2_0_5 ;
    wire \VPP_VDDQ.count_2_1_5_cascade_ ;
    wire \VPP_VDDQ.count_2_0_8 ;
    wire \VPP_VDDQ.count_2_1_8 ;
    wire \VPP_VDDQ.count_2_0_2 ;
    wire \VPP_VDDQ.count_2_1_2_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_2_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2_0_15 ;
    wire \VPP_VDDQ.N_551 ;
    wire vpp_en;
    wire \VPP_VDDQ.count_2_1_14_cascade_ ;
    wire \VPP_VDDQ.countZ0Z_5 ;
    wire \VPP_VDDQ.countZ0Z_4 ;
    wire \VPP_VDDQ.countZ0Z_3 ;
    wire \VPP_VDDQ.countZ0Z_7 ;
    wire \VPP_VDDQ.curr_stateZ0Z_1 ;
    wire N_325;
    wire \VPP_VDDQ.delayed_vddq_pwrgdZ0 ;
    wire VPP_VDDQ_curr_state_0;
    wire N_325_cascade_;
    wire \VPP_VDDQ.delayed_vddq_pwrgd_0 ;
    wire VCCST_EN_i_0;
    wire \VPP_VDDQ.N_541 ;
    wire \VPP_VDDQ.countZ0Z_14 ;
    wire \VPP_VDDQ.countZ0Z_13 ;
    wire \VPP_VDDQ.countZ0Z_15 ;
    wire \VPP_VDDQ.countZ0Z_12 ;
    wire \VPP_VDDQ.un6_count_10 ;
    wire \VPP_VDDQ.un6_count_9_cascade_ ;
    wire \VPP_VDDQ.un6_count ;
    wire \VPP_VDDQ.countZ0Z_9 ;
    wire \VPP_VDDQ.countZ0Z_0 ;
    wire \VPP_VDDQ.countZ0Z_8 ;
    wire \VPP_VDDQ.countZ0Z_11 ;
    wire \VPP_VDDQ.un6_count_11 ;
    wire \VPP_VDDQ.countZ0Z_6 ;
    wire \VPP_VDDQ.countZ0Z_2 ;
    wire \VPP_VDDQ.countZ0Z_10 ;
    wire \VPP_VDDQ.countZ0Z_1 ;
    wire \VPP_VDDQ.un6_count_8 ;
    wire v1p8a_en;
    wire \POWERLED.mult1_un82_sum ;
    wire bfn_9_1_0_;
    wire \POWERLED.mult1_un75_sum_i ;
    wire \POWERLED.mult1_un82_sum_cry_3_s ;
    wire \POWERLED.mult1_un82_sum_cry_2_c ;
    wire \POWERLED.mult1_un82_sum_cry_4_s ;
    wire \POWERLED.mult1_un82_sum_cry_3_c ;
    wire \POWERLED.mult1_un82_sum_cry_5_s ;
    wire \POWERLED.mult1_un82_sum_cry_4_c ;
    wire \POWERLED.mult1_un82_sum_cry_6_s ;
    wire \POWERLED.mult1_un82_sum_cry_5_c ;
    wire \POWERLED.mult1_un89_sum_axb_8 ;
    wire \POWERLED.mult1_un82_sum_cry_6_c ;
    wire \POWERLED.mult1_un82_sum_cry_7 ;
    wire \POWERLED.mult1_un82_sum_s_8 ;
    wire \POWERLED.mult1_un75_sum ;
    wire bfn_9_2_0_;
    wire \POWERLED.mult1_un68_sum_i ;
    wire \POWERLED.mult1_un75_sum_cry_3_s ;
    wire \POWERLED.mult1_un75_sum_cry_2 ;
    wire \POWERLED.mult1_un75_sum_cry_4_s ;
    wire \POWERLED.mult1_un75_sum_cry_3 ;
    wire \POWERLED.mult1_un75_sum_cry_5_s ;
    wire \POWERLED.mult1_un75_sum_cry_4 ;
    wire \POWERLED.mult1_un75_sum_cry_6_s ;
    wire \POWERLED.mult1_un75_sum_cry_5 ;
    wire \POWERLED.mult1_un68_sum_i_0_8 ;
    wire \POWERLED.mult1_un82_sum_axb_8 ;
    wire \POWERLED.mult1_un75_sum_cry_6 ;
    wire \POWERLED.mult1_un75_sum_cry_7 ;
    wire \POWERLED.mult1_un75_sum_s_8 ;
    wire \POWERLED.mult1_un75_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un75_sum_i_0_8 ;
    wire \POWERLED.mult1_un54_sum ;
    wire bfn_9_3_0_;
    wire \POWERLED.un1_dutycycle_53_i_28 ;
    wire \POWERLED.mult1_un54_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6 ;
    wire \POWERLED.mult1_un54_sum_cry_7 ;
    wire \POWERLED.mult1_un47_sum_l_fx_6 ;
    wire \POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434 ;
    wire bfn_9_4_0_;
    wire \POWERLED.un1_dutycycle_53_i_29 ;
    wire \POWERLED.mult1_un47_sum_cry_2 ;
    wire \POWERLED.mult1_un47_sum_axb_4 ;
    wire \POWERLED.mult1_un47_sum_cry_4_s ;
    wire \POWERLED.mult1_un47_sum_cry_3 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_4 ;
    wire \POWERLED.mult1_un47_sum_cry_5_s ;
    wire \POWERLED.mult1_un47_sum_cry_4 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_5 ;
    wire \POWERLED.mult1_un47_sum_cry_6_s ;
    wire \POWERLED.mult1_un47_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_7_THRU_CO ;
    wire \POWERLED.mult1_un47_sum_cry_6 ;
    wire \POWERLED.mult1_un61_sum_i_8 ;
    wire \POWERLED.mult1_un47_sum_cry_3_s ;
    wire \POWERLED.mult1_un47_sum_l_fx_3 ;
    wire \POWERLED.dutycycleZ0Z_13_cascade_ ;
    wire \POWERLED.N_2293_i_cascade_ ;
    wire \POWERLED.dutycycle_eena_2 ;
    wire \POWERLED.dutycycleZ1Z_9 ;
    wire \POWERLED.dutycycle_eena_2_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_2_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_13 ;
    wire \POWERLED.un1_dutycycle_53_7_a0_0 ;
    wire \POWERLED.dutycycleZ0Z_9_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_13_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_14 ;
    wire \POWERLED.un1_dutycycle_53_12_0 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_13 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_14 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_7 ;
    wire \POWERLED.un1_dutycycle_53_57_a0_d_cascade_ ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_13 ;
    wire bfn_9_7_0_;
    wire \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_0 ;
    wire \POWERLED.un1_dutycycle_94_cry_1_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ;
    wire \POWERLED.un1_dutycycle_94_cry_2_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ;
    wire \POWERLED.un1_dutycycle_94_cry_3_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_4 ;
    wire \POWERLED.un1_dutycycle_94_cry_5_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ;
    wire \POWERLED.un1_dutycycle_94_cry_6_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_7_cZ0 ;
    wire bfn_9_8_0_;
    wire \POWERLED.un1_dutycycle_94_cry_8_c_RNI3B2UZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_8 ;
    wire \POWERLED.un1_dutycycle_94_cry_9 ;
    wire \POWERLED.un1_dutycycle_94_cry_10 ;
    wire \POWERLED.un1_dutycycle_94_cry_11 ;
    wire \POWERLED.un1_dutycycle_94_cry_12_c_RNIE4NBZ0Z1 ;
    wire \POWERLED.un1_dutycycle_94_cry_12 ;
    wire \POWERLED.N_341_i ;
    wire \POWERLED.un1_dutycycle_94_cry_13 ;
    wire \POWERLED.un1_dutycycle_94_cry_14 ;
    wire \POWERLED.un1_dutycycle_94_cry_14_c_RNIG8PBZ0Z1 ;
    wire \POWERLED.N_292 ;
    wire \POWERLED.dutycycle_1_0_iv_i_a3_0_2_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ;
    wire \POWERLED.N_145 ;
    wire m57_i_o2_3;
    wire \POWERLED.un1_dutycycle_94_cry_5_c_RNIZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_5_c_RNIEVTSZ0Z3 ;
    wire \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ;
    wire \POWERLED.dutycycle_set_1 ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_6 ;
    wire \POWERLED.N_258 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_5 ;
    wire \POWERLED.N_505 ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_5_cascade_ ;
    wire \POWERLED.dutycycle_RNI2O4A1Z0Z_6 ;
    wire \POWERLED.func_state_RNIOGRS_0Z0Z_1_cascade_ ;
    wire \POWERLED.N_487 ;
    wire \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ;
    wire \POWERLED.N_379_N ;
    wire G_22_i_a2_1;
    wire SUSWARN_N_fast;
    wire \POWERLED.N_564 ;
    wire v5s_ok;
    wire vccst_cpu_ok;
    wire v33s_ok;
    wire dsw_pwrok;
    wire v5s_enn;
    wire \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_ ;
    wire vccin_en;
    wire N_323;
    wire N_323_cascade_;
    wire v33a_ok;
    wire slp_susn;
    wire v1p8a_ok;
    wire v5a_ok;
    wire N_171_cascade_;
    wire vr_ready_vccinaux;
    wire N_283;
    wire RSMRST_PWRGD_curr_state_0;
    wire N_283_cascade_;
    wire \RSMRST_PWRGD.curr_stateZ0Z_1 ;
    wire rsmrstn;
    wire \VPP_VDDQ.un9_clk_100khz_9 ;
    wire \VPP_VDDQ.un9_clk_100khz_0_cascade_ ;
    wire bfn_9_13_0_;
    wire \VPP_VDDQ.count_2Z0Z_2 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_1 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_2 ;
    wire \VPP_VDDQ.count_2Z0Z_4 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_3 ;
    wire \VPP_VDDQ.count_2Z0Z_5 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_4 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_6 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_5 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_6 ;
    wire \VPP_VDDQ.count_2Z0Z_8 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_8 ;
    wire bfn_9_14_0_;
    wire \VPP_VDDQ.un1_count_2_1_cry_9 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_10 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_11 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_12 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_13 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ;
    wire \VPP_VDDQ.count_2Z0Z_15 ;
    wire \VPP_VDDQ.count_2Z0Z_14 ;
    wire \VPP_VDDQ.count_2_1_6 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661 ;
    wire \VPP_VDDQ.count_2Z0Z_6 ;
    wire \VPP_VDDQ.count_2_1_9_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ;
    wire \VPP_VDDQ.count_2_0_9 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ;
    wire \VPP_VDDQ.count_2_0_10 ;
    wire \VPP_VDDQ.count_2_1_10_cascade_ ;
    wire \VPP_VDDQ.count_2_1_12_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_12 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0 ;
    wire \VPP_VDDQ.count_2_0_12 ;
    wire \VPP_VDDQ.count_2_1_13_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_13 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ;
    wire \VPP_VDDQ.count_2_0_13 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ;
    wire \VPP_VDDQ.count_2_0_14 ;
    wire \POWERLED.mult1_un68_sum ;
    wire bfn_11_2_0_;
    wire \POWERLED.mult1_un61_sum_i ;
    wire \POWERLED.mult1_un68_sum_cry_3_s ;
    wire \POWERLED.mult1_un68_sum_cry_2 ;
    wire \POWERLED.mult1_un68_sum_cry_4_s ;
    wire \POWERLED.mult1_un68_sum_cry_3 ;
    wire \POWERLED.mult1_un68_sum_cry_5_s ;
    wire \POWERLED.mult1_un68_sum_cry_4 ;
    wire \POWERLED.mult1_un68_sum_cry_6_s ;
    wire \POWERLED.mult1_un68_sum_cry_5 ;
    wire \POWERLED.mult1_un75_sum_axb_8 ;
    wire \POWERLED.mult1_un68_sum_cry_6 ;
    wire \POWERLED.mult1_un68_sum_cry_7 ;
    wire \POWERLED.mult1_un68_sum_s_8 ;
    wire \POWERLED.mult1_un61_sum ;
    wire bfn_11_3_0_;
    wire \POWERLED.mult1_un54_sum_i ;
    wire \POWERLED.mult1_un61_sum_cry_3_s ;
    wire \POWERLED.mult1_un61_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3_s ;
    wire \POWERLED.mult1_un61_sum_cry_4_s ;
    wire \POWERLED.mult1_un61_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4_s ;
    wire \POWERLED.mult1_un61_sum_cry_5_s ;
    wire \POWERLED.mult1_un61_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_s_8 ;
    wire \POWERLED.mult1_un54_sum_cry_5_s ;
    wire \POWERLED.mult1_un61_sum_cry_6_s ;
    wire \POWERLED.mult1_un61_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6_s ;
    wire \POWERLED.mult1_un54_sum_i_8 ;
    wire \POWERLED.mult1_un68_sum_axb_8 ;
    wire \POWERLED.mult1_un61_sum_cry_6 ;
    wire \POWERLED.mult1_un61_sum_axb_8 ;
    wire \POWERLED.mult1_un61_sum_cry_7 ;
    wire \POWERLED.mult1_un61_sum_s_8 ;
    wire \POWERLED.mult1_un61_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un61_sum_i_0_8 ;
    wire \POWERLED.un1_dutycycle_94_cry_13_c_RNIF6OBZ0Z1 ;
    wire \POWERLED.dutycycle_eena_11 ;
    wire \POWERLED.dutycycleZ0Z_14 ;
    wire \POWERLED.un1_dutycycle_53_8_a3_1_0_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_9 ;
    wire \POWERLED.un1_dutycycle_53_7_4_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_13 ;
    wire \POWERLED.un1_N_5_mux ;
    wire \POWERLED.un1_dutycycle_53_8_6_tz_sx_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_8_2_0_tz ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_10 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_9 ;
    wire \POWERLED.dutycycleZ1Z_8 ;
    wire \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ;
    wire \POWERLED.dutycycleZ0Z_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_11_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_57_a0_1_1 ;
    wire \POWERLED.un1_dutycycle_53_2_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI_10Z0Z_10 ;
    wire \POWERLED.dutycycle_RNI_11Z0Z_10 ;
    wire \POWERLED.un1_dutycycle_53_13_a1_1_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_11 ;
    wire \POWERLED.un1_dutycycle_94_cry_10_c_RNIC0LBZ0Z1 ;
    wire \POWERLED.dutycycle_eena_7 ;
    wire \POWERLED.dutycycleZ0Z_7_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_46_a3_1 ;
    wire \POWERLED.un1_dutycycle_53_46_a3_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_6Z0Z_7 ;
    wire \POWERLED.un1_dutycycle_53_46_a3_d ;
    wire \POWERLED.dutycycle_eena_9_cascade_ ;
    wire \POWERLED.dutycycle_eena_5_0_s_tz_isoZ0 ;
    wire \POWERLED.dutycycle_eena_4 ;
    wire \POWERLED.dutycycleZ1Z_10 ;
    wire \POWERLED.dutycycle_eena_4_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_9_c_RNI4D3UZ0 ;
    wire \POWERLED.dutycycleZ0Z_5_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_12 ;
    wire \POWERLED.dutycycle_eena_9 ;
    wire \POWERLED.un1_dutycycle_94_cry_11_c_RNID2MBZ0Z1 ;
    wire \POWERLED.un1_dutycycle_53_7_3_0_1 ;
    wire \POWERLED.dutycycleZ0Z_10_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_7_3 ;
    wire dutycycle_RNINBHJ5_0_2;
    wire \POWERLED.dutycycle_RNI_5Z0Z_1 ;
    wire \POWERLED.un1_dutycycle_172_m2s4_1_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_6 ;
    wire \POWERLED.un1_dutycycle_172_m2s4_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_1 ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_3 ;
    wire \POWERLED.N_414 ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_3_cascade_ ;
    wire \POWERLED.g0_i_1_1_0 ;
    wire \POWERLED.func_state_RNI56A8Z0Z_0 ;
    wire \POWERLED.N_239 ;
    wire \POWERLED.N_462 ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_6 ;
    wire \POWERLED.un1_clk_100khz_52_and_i_0_m3_1_rn_1_cascade_ ;
    wire POWERLED_un1_clk_100khz_52_and_i_0_m3_1;
    wire \POWERLED.m69_0_o2_2 ;
    wire RSMRSTn_rep1;
    wire N_110_0;
    wire \RSMRST_PWRGD.un4_count_9_cascade_ ;
    wire \RSMRST_PWRGD.N_1_i ;
    wire \RSMRST_PWRGD.un4_count_8 ;
    wire \RSMRST_PWRGD.un4_count_10 ;
    wire \RSMRST_PWRGD.un4_count_11 ;
    wire \RSMRST_PWRGD.N_445_i ;
    wire \RSMRST_PWRGD.countZ0Z_0 ;
    wire bfn_11_12_0_;
    wire \RSMRST_PWRGD.countZ0Z_1 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_0 ;
    wire \RSMRST_PWRGD.countZ0Z_2 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_1 ;
    wire \RSMRST_PWRGD.countZ0Z_3 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_2 ;
    wire \RSMRST_PWRGD.countZ0Z_4 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_3 ;
    wire \RSMRST_PWRGD.countZ0Z_5 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_4 ;
    wire \RSMRST_PWRGD.countZ0Z_6 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_5 ;
    wire \RSMRST_PWRGD.countZ0Z_7 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_6 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_7 ;
    wire \RSMRST_PWRGD.countZ0Z_8 ;
    wire bfn_11_13_0_;
    wire \RSMRST_PWRGD.countZ0Z_9 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_8 ;
    wire \RSMRST_PWRGD.countZ0Z_10 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_9 ;
    wire \RSMRST_PWRGD.countZ0Z_11 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_10 ;
    wire \RSMRST_PWRGD.countZ0Z_12 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_11 ;
    wire \RSMRST_PWRGD.countZ0Z_13 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_12 ;
    wire N_42_g;
    wire \RSMRST_PWRGD.countZ0Z_14 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_13 ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \RSMRST_PWRGD.un1_count_1_cry_14 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_11_14_0_;
    wire \RSMRST_PWRGD.countZ0Z_15 ;
    wire \RSMRST_PWRGD.N_42_2 ;
    wire G_12;
    wire \VPP_VDDQ.curr_state_2_0_0 ;
    wire \VPP_VDDQ.N_190_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ;
    wire \VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2_0_3 ;
    wire \VPP_VDDQ.count_2_1_3_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_3 ;
    wire \VPP_VDDQ.N_537_0_cascade_ ;
    wire \VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0_cascade_ ;
    wire \VPP_VDDQ.N_537_0 ;
    wire \VPP_VDDQ.N_28_i ;
    wire \VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0 ;
    wire \VPP_VDDQ.delayed_vddq_okZ0 ;
    wire \VPP_VDDQ.delayed_vddq_ok_en ;
    wire VPP_VDDQ_delayed_vddq_ok;
    wire \POWERLED.dutycycle_RNI_2Z0Z_9_cascade_ ;
    wire \POWERLED.dutycycle_RNI_6Z0Z_9 ;
    wire \POWERLED.un1_dutycycle_53_4_a0_1 ;
    wire \POWERLED.un1_dutycycle_53_4_a0_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_7_2 ;
    wire \POWERLED.un1_dutycycle_53_8_1 ;
    wire \POWERLED.un1_dutycycle_53_8_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_9 ;
    wire \POWERLED.dutycycle_RNIZ0Z_5 ;
    wire \POWERLED.dutycycle_eena_10 ;
    wire \POWERLED.N_507 ;
    wire \POWERLED.N_84_f0_cascade_ ;
    wire G_156;
    wire \POWERLED.dutycycle_en_3 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_11 ;
    wire \POWERLED.N_12_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_3 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_4 ;
    wire \POWERLED.un1_dutycycle_53_25_0_tz ;
    wire \POWERLED.N_6 ;
    wire \POWERLED.dutycycleZ0Z_12 ;
    wire POWERLED_func_state_0_sqmuxa;
    wire \POWERLED.N_2191_i_cascade_ ;
    wire \POWERLED.N_282_N ;
    wire \POWERLED.dutycycle_eena_12 ;
    wire \POWERLED.g0_i_i_a6_0_2 ;
    wire \POWERLED.dutycycle_RNIZ0Z_4 ;
    wire \POWERLED.dutycycleZ0Z_13 ;
    wire \POWERLED.g0_i_i_1 ;
    wire \POWERLED.un1_dutycycle_53_axb_11_1 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_14 ;
    wire \POWERLED.N_2293_i ;
    wire \POWERLED.un1_dutycycle_53_4_1 ;
    wire \POWERLED.dutycycle_RNI_6Z0Z_4_cascade_ ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_4 ;
    wire \POWERLED.o2_cascade_ ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_10 ;
    wire \POWERLED.dutycycleZ0Z_7 ;
    wire \POWERLED.dutycycleZ0Z_5 ;
    wire \POWERLED.dutycycleZ0Z_2 ;
    wire \POWERLED.dutycycleZ0Z_1 ;
    wire \POWERLED.N_2191_i ;
    wire \POWERLED.dutycycleZ0Z_10 ;
    wire \POWERLED.N_2187_i ;
    wire \POWERLED.un2_count_clk_17_0_0_a2_5_cascade_ ;
    wire \POWERLED.un2_count_clk_17_0_0_a2_0 ;
    wire \POWERLED.N_501 ;
    wire \POWERLED.dutycycleZ0Z_8 ;
    wire \POWERLED.dutycycleZ0Z_4 ;
    wire \POWERLED.dutycycleZ0Z_6 ;
    wire func_state_RNITGMHB_0_1;
    wire \POWERLED.un2_count_clk_17_0_1 ;
    wire \POWERLED.un2_count_clk_17_0_1_cascade_ ;
    wire \POWERLED.dutycycle ;
    wire \POWERLED.dutycycleZ0Z_0 ;
    wire \POWERLED.N_493 ;
    wire \POWERLED.g1_0_7 ;
    wire \POWERLED.g1_0_2 ;
    wire \POWERLED.g1_0_8_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_6 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_6 ;
    wire RSMRSTn_fast;
    wire \RSMRST_PWRGD.N_8_0_0_cascade_ ;
    wire func_state_RNIOGRS_1;
    wire dutycycle_RNIKBMSJ_0_5;
    wire POWERLED_g1;
    wire \RSMRST_PWRGD.N_9_0_cascade_ ;
    wire N_46;
    wire \RSMRST_PWRGD.N_11 ;
    wire \POWERLED.N_341 ;
    wire \POWERLED.N_335 ;
    wire N_22_0;
    wire N_22_0_cascade_;
    wire N_2145_i;
    wire g0_0_1;
    wire slp_s4n;
    wire slp_s3n;
    wire func_state_RNI_3_0;
    wire gpio_fpga_soc_4;
    wire \POWERLED.dutycycle_1_0_iv_i_a2_sx_5 ;
    wire \VPP_VDDQ.N_2112_i ;
    wire \VPP_VDDQ.count_2Z0Z_9 ;
    wire \VPP_VDDQ.count_2_1_7_cascade_ ;
    wire \VPP_VDDQ.un9_clk_100khz_10 ;
    wire \VPP_VDDQ.count_2Z0Z_10 ;
    wire \VPP_VDDQ.un9_clk_100khz_7_cascade_ ;
    wire \VPP_VDDQ.un9_clk_100khz_13 ;
    wire \VPP_VDDQ.count_2_1_0_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2_0_0 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7 ;
    wire \VPP_VDDQ.count_2Z0Z_7 ;
    wire \VPP_VDDQ.count_2_1_7 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_7 ;
    wire \VPP_VDDQ.count_2_RNIZ0Z_1_cascade_ ;
    wire \VPP_VDDQ.count_2_1_1_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_axb_1 ;
    wire \VPP_VDDQ.count_2_1_1 ;
    wire \VPP_VDDQ.count_2Z0Z_0 ;
    wire \VPP_VDDQ.un9_clk_100khz_1 ;
    wire \VPP_VDDQ.count_2_RNIZ0Z_1 ;
    wire \VPP_VDDQ.count_2Z0Z_1 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ;
    wire \VPP_VDDQ.count_2_0_11 ;
    wire \VPP_VDDQ.count_2_1_11_cascade_ ;
    wire \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ;
    wire \VPP_VDDQ.count_2Z0Z_11 ;
    wire \VPP_VDDQ.N_178_cascade_ ;
    wire suswarn_n;
    wire \VPP_VDDQ.N_1_i ;
    wire \VPP_VDDQ.curr_state_2Z0Z_0 ;
    wire \VPP_VDDQ.curr_state_2Z0Z_1 ;
    wire vddq_ok;
    wire \VPP_VDDQ.curr_state_2_0_1 ;
    wire fpga_osc;
    wire N_587_g;
    wire _gnd_net_;

    defparam ipInertedIOPad_VR_READY_VCCINAUX_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VR_READY_VCCINAUX_iopad (
            .OE(N__34571),
            .DIN(N__34570),
            .DOUT(N__34569),
            .PACKAGEPIN(VR_READY_VCCINAUX));
    defparam ipInertedIOPad_VR_READY_VCCINAUX_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCINAUX_preio (
            .PADOEN(N__34571),
            .PADOUT(N__34570),
            .PADIN(N__34569),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccinaux),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_ENn_iopad (
            .OE(N__34562),
            .DIN(N__34561),
            .DOUT(N__34560),
            .PACKAGEPIN(V33A_ENn));
    defparam ipInertedIOPad_V33A_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33A_ENn_preio (
            .PADOEN(N__34562),
            .PADOUT(N__34561),
            .PADIN(N__34560),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V1P8A_EN_iopad (
            .OE(N__34553),
            .DIN(N__34552),
            .DOUT(N__34551),
            .PACKAGEPIN(V1P8A_EN));
    defparam ipInertedIOPad_V1P8A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V1P8A_EN_preio (
            .PADOEN(N__34553),
            .PADOUT(N__34552),
            .PADIN(N__34551),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23620),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDDQ_EN_iopad (
            .OE(N__34544),
            .DIN(N__34543),
            .DOUT(N__34542),
            .PACKAGEPIN(VDDQ_EN));
    defparam ipInertedIOPad_VDDQ_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDDQ_EN_preio (
            .PADOEN(N__34544),
            .PADOUT(N__34543),
            .PADIN(N__34542),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16072),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad (
            .OE(N__34535),
            .DIN(N__34534),
            .DOUT(N__34533),
            .PACKAGEPIN(VCCST_OVERRIDE_3V3));
    defparam ipInertedIOPad_VCCST_OVERRIDE_3V3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_OVERRIDE_3V3_preio (
            .PADOEN(N__34535),
            .PADOUT(N__34534),
            .PADIN(N__34533),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_OK_iopad (
            .OE(N__34526),
            .DIN(N__34525),
            .DOUT(N__34524),
            .PACKAGEPIN(V5S_OK));
    defparam ipInertedIOPad_V5S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5S_OK_preio (
            .PADOEN(N__34526),
            .PADOUT(N__34525),
            .PADIN(N__34524),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S3n_iopad (
            .OE(N__34517),
            .DIN(N__34516),
            .DOUT(N__34515),
            .PACKAGEPIN(SLP_S3n));
    defparam ipInertedIOPad_SLP_S3n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S3n_preio (
            .PADOEN(N__34517),
            .PADOUT(N__34516),
            .PADIN(N__34515),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s3n),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S0n_iopad (
            .OE(N__34508),
            .DIN(N__34507),
            .DOUT(N__34506),
            .PACKAGEPIN(SLP_S0n));
    defparam ipInertedIOPad_SLP_S0n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S0n_preio (
            .PADOEN(N__34508),
            .PADOUT(N__34507),
            .PADIN(N__34506),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_ENn_iopad (
            .OE(N__34499),
            .DIN(N__34498),
            .DOUT(N__34497),
            .PACKAGEPIN(V5S_ENn));
    defparam ipInertedIOPad_V5S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5S_ENn_preio (
            .PADOEN(N__34499),
            .PADOUT(N__34498),
            .PADIN(N__34497),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25004),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V1P8A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V1P8A_OK_iopad (
            .OE(N__34490),
            .DIN(N__34489),
            .DOUT(N__34488),
            .PACKAGEPIN(V1P8A_OK));
    defparam ipInertedIOPad_V1P8A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V1P8A_OK_preio (
            .PADOEN(N__34490),
            .PADOUT(N__34489),
            .PADIN(N__34488),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v1p8a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTNn_iopad (
            .OE(N__34481),
            .DIN(N__34480),
            .DOUT(N__34479),
            .PACKAGEPIN(PWRBTNn));
    defparam ipInertedIOPad_PWRBTNn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PWRBTNn_preio (
            .PADOEN(N__34481),
            .PADOUT(N__34480),
            .PADIN(N__34479),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTN_LED_iopad (
            .OE(N__34472),
            .DIN(N__34471),
            .DOUT(N__34470),
            .PACKAGEPIN(PWRBTN_LED));
    defparam ipInertedIOPad_PWRBTN_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PWRBTN_LED_preio (
            .PADOEN(N__34472),
            .PADOUT(N__34471),
            .PADIN(N__34470),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16213),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_2_iopad (
            .OE(N__34463),
            .DIN(N__34462),
            .DOUT(N__34461),
            .PACKAGEPIN(GPIO_FPGA_SoC_2));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_2_preio (
            .PADOEN(N__34463),
            .PADOUT(N__34462),
            .PADIN(N__34461),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad (
            .OE(N__34454),
            .DIN(N__34453),
            .DOUT(N__34452),
            .PACKAGEPIN(VCCIN_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__34454),
            .PADOUT(N__34453),
            .PADIN(N__34452),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_SUSn_iopad (
            .OE(N__34445),
            .DIN(N__34444),
            .DOUT(N__34443),
            .PACKAGEPIN(SLP_SUSn));
    defparam ipInertedIOPad_SLP_SUSn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_SUSn_preio (
            .PADOEN(N__34445),
            .PADOUT(N__34444),
            .PADIN(N__34443),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_susn),
            .DIN1());
    IO_PAD ipInertedIOPad_CPU_C10_GATE_N_iopad (
            .OE(N__34436),
            .DIN(N__34435),
            .DOUT(N__34434),
            .PACKAGEPIN(CPU_C10_GATE_N));
    defparam ipInertedIOPad_CPU_C10_GATE_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_CPU_C10_GATE_N_preio (
            .PADOEN(N__34436),
            .PADOUT(N__34435),
            .PADIN(N__34434),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_EN_iopad (
            .OE(N__34427),
            .DIN(N__34426),
            .DOUT(N__34425),
            .PACKAGEPIN(VCCST_EN));
    defparam ipInertedIOPad_VCCST_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_EN_preio (
            .PADOEN(N__34427),
            .PADOUT(N__34426),
            .PADIN(N__34425),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17002),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V33DSW_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V33DSW_OK_iopad (
            .OE(N__34418),
            .DIN(N__34417),
            .DOUT(N__34416),
            .PACKAGEPIN(V33DSW_OK));
    defparam ipInertedIOPad_V33DSW_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33DSW_OK_preio (
            .PADOEN(N__34418),
            .PADOUT(N__34417),
            .PADIN(N__34416),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33dsw_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_TPM_GPIO_iopad (
            .OE(N__34409),
            .DIN(N__34408),
            .DOUT(N__34407),
            .PACKAGEPIN(TPM_GPIO));
    defparam ipInertedIOPad_TPM_GPIO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_TPM_GPIO_preio (
            .PADOEN(N__34409),
            .PADOUT(N__34408),
            .PADIN(N__34407),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSWARN_N_iopad (
            .OE(N__34400),
            .DIN(N__34399),
            .DOUT(N__34398),
            .PACKAGEPIN(SUSWARN_N));
    defparam ipInertedIOPad_SUSWARN_N_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SUSWARN_N_preio (
            .PADOEN(N__34400),
            .PADOUT(N__34399),
            .PADIN(N__34398),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__33932),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PLTRSTn_iopad (
            .OE(N__34391),
            .DIN(N__34390),
            .DOUT(N__34389),
            .PACKAGEPIN(PLTRSTn));
    defparam ipInertedIOPad_PLTRSTn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PLTRSTn_preio (
            .PADOEN(N__34391),
            .PADOUT(N__34390),
            .PADIN(N__34389),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_4_iopad (
            .OE(N__34382),
            .DIN(N__34381),
            .DOUT(N__34380),
            .PACKAGEPIN(GPIO_FPGA_SoC_4));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_4_preio (
            .PADOEN(N__34382),
            .PADOUT(N__34381),
            .PADIN(N__34380),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_4),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_READY_VCCIN_iopad (
            .OE(N__34373),
            .DIN(N__34372),
            .DOUT(N__34371),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam ipInertedIOPad_VR_READY_VCCIN_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCIN_preio (
            .PADOEN(N__34373),
            .PADOUT(N__34372),
            .PADIN(N__34371),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccin),
            .DIN1());
    defparam ipInertedIOPad_V5A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V5A_OK_iopad (
            .OE(N__34364),
            .DIN(N__34363),
            .DOUT(N__34362),
            .PACKAGEPIN(V5A_OK));
    defparam ipInertedIOPad_V5A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5A_OK_preio (
            .PADOEN(N__34364),
            .PADOUT(N__34363),
            .PADIN(N__34362),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_RSMRSTn_iopad (
            .OE(N__34355),
            .DIN(N__34354),
            .DOUT(N__34353),
            .PACKAGEPIN(RSMRSTn));
    defparam ipInertedIOPad_RSMRSTn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RSMRSTn_preio (
            .PADOEN(N__34355),
            .PADOUT(N__34354),
            .PADIN(N__34353),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25153),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_OSC_iopad (
            .OE(N__34346),
            .DIN(N__34345),
            .DOUT(N__34344),
            .PACKAGEPIN(FPGA_OSC));
    defparam ipInertedIOPad_FPGA_OSC_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_OSC_preio (
            .PADOEN(N__34346),
            .PADOUT(N__34345),
            .PADIN(N__34344),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(fpga_osc),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_PWRGD_iopad (
            .OE(N__34337),
            .DIN(N__34336),
            .DOUT(N__34335),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam ipInertedIOPad_VCCST_PWRGD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_PWRGD_preio (
            .PADOEN(N__34337),
            .PADOUT(N__34336),
            .PADIN(N__34335),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17893),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SYS_PWROK_iopad (
            .OE(N__34328),
            .DIN(N__34327),
            .DOUT(N__34326),
            .PACKAGEPIN(SYS_PWROK));
    defparam ipInertedIOPad_SYS_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SYS_PWROK_preio (
            .PADOEN(N__34328),
            .PADOUT(N__34327),
            .PADIN(N__34326),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20752),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO2_iopad (
            .OE(N__34319),
            .DIN(N__34318),
            .DOUT(N__34317),
            .PACKAGEPIN(SPI_FP_IO2));
    defparam ipInertedIOPad_SPI_FP_IO2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO2_preio (
            .PADOEN(N__34319),
            .PADOUT(N__34318),
            .PADIN(N__34317),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE1_FPGA_iopad (
            .OE(N__34310),
            .DIN(N__34309),
            .DOUT(N__34308),
            .PACKAGEPIN(SATAXPCIE1_FPGA));
    defparam ipInertedIOPad_SATAXPCIE1_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE1_FPGA_preio (
            .PADOEN(N__34310),
            .PADOUT(N__34309),
            .PADIN(N__34308),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_1_iopad (
            .OE(N__34301),
            .DIN(N__34300),
            .DOUT(N__34299),
            .PACKAGEPIN(GPIO_FPGA_EXP_1));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_1_preio (
            .PADOEN(N__34301),
            .PADOUT(N__34300),
            .PADIN(N__34299),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad (
            .OE(N__34292),
            .DIN(N__34291),
            .DOUT(N__34290),
            .PACKAGEPIN(VCCINAUX_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__34292),
            .PADOUT(N__34291),
            .PADIN(N__34290),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PE_iopad (
            .OE(N__34283),
            .DIN(N__34282),
            .DOUT(N__34281),
            .PACKAGEPIN(VCCINAUX_VR_PE));
    defparam ipInertedIOPad_VCCINAUX_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PE_preio (
            .PADOEN(N__34283),
            .PADOUT(N__34282),
            .PADIN(N__34281),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27255),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_HDA_SDO_ATP_iopad (
            .OE(N__34274),
            .DIN(N__34273),
            .DOUT(N__34272),
            .PACKAGEPIN(HDA_SDO_ATP));
    defparam ipInertedIOPad_HDA_SDO_ATP_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_HDA_SDO_ATP_preio (
            .PADOEN(N__34274),
            .PADOUT(N__34273),
            .PADIN(N__34272),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__15322),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_2_iopad (
            .OE(N__34265),
            .DIN(N__34264),
            .DOUT(N__34263),
            .PACKAGEPIN(GPIO_FPGA_EXP_2));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_2_preio (
            .PADOEN(N__34265),
            .PADOUT(N__34264),
            .PADIN(N__34263),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VPP_EN_iopad (
            .OE(N__34256),
            .DIN(N__34255),
            .DOUT(N__34254),
            .PACKAGEPIN(VPP_EN));
    defparam ipInertedIOPad_VPP_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VPP_EN_preio (
            .PADOEN(N__34256),
            .PADOUT(N__34255),
            .PADIN(N__34254),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23128),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VDDQ_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VDDQ_OK_iopad (
            .OE(N__34247),
            .DIN(N__34246),
            .DOUT(N__34245),
            .PACKAGEPIN(VDDQ_OK));
    defparam ipInertedIOPad_VDDQ_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDDQ_OK_preio (
            .PADOEN(N__34247),
            .PADOUT(N__34246),
            .PADIN(N__34245),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vddq_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSACK_N_iopad (
            .OE(N__34238),
            .DIN(N__34237),
            .DOUT(N__34236),
            .PACKAGEPIN(SUSACK_N));
    defparam ipInertedIOPad_SUSACK_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSACK_N_preio (
            .PADOEN(N__34238),
            .PADOUT(N__34237),
            .PADIN(N__34236),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S4n_iopad (
            .OE(N__34229),
            .DIN(N__34228),
            .DOUT(N__34227),
            .PACKAGEPIN(SLP_S4n));
    defparam ipInertedIOPad_SLP_S4n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S4n_preio (
            .PADOEN(N__34229),
            .PADOUT(N__34228),
            .PADIN(N__34227),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s4n),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_CPU_OK_iopad (
            .OE(N__34220),
            .DIN(N__34219),
            .DOUT(N__34218),
            .PACKAGEPIN(VCCST_CPU_OK));
    defparam ipInertedIOPad_VCCST_CPU_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_CPU_OK_preio (
            .PADOEN(N__34220),
            .PADOUT(N__34219),
            .PADIN(N__34218),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vccst_cpu_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_EN_iopad (
            .OE(N__34211),
            .DIN(N__34210),
            .DOUT(N__34209),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam ipInertedIOPad_VCCINAUX_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_EN_preio (
            .PADOEN(N__34211),
            .PADOUT(N__34210),
            .PADIN(N__34209),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25306),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_OK_iopad (
            .OE(N__34202),
            .DIN(N__34201),
            .DOUT(N__34200),
            .PACKAGEPIN(V33S_OK));
    defparam ipInertedIOPad_V33S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33S_OK_preio (
            .PADOEN(N__34202),
            .PADOUT(N__34201),
            .PADIN(N__34200),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_ENn_iopad (
            .OE(N__34193),
            .DIN(N__34192),
            .DOUT(N__34191),
            .PACKAGEPIN(V33S_ENn));
    defparam ipInertedIOPad_V33S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33S_ENn_preio (
            .PADOEN(N__34193),
            .PADOUT(N__34192),
            .PADIN(N__34191),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25009),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_1_iopad (
            .OE(N__34184),
            .DIN(N__34183),
            .DOUT(N__34182),
            .PACKAGEPIN(GPIO_FPGA_SoC_1));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_1_preio (
            .PADOEN(N__34184),
            .PADOUT(N__34183),
            .PADIN(N__34182),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_1),
            .DIN1());
    IO_PAD ipInertedIOPad_DSW_PWROK_iopad (
            .OE(N__34175),
            .DIN(N__34174),
            .DOUT(N__34173),
            .PACKAGEPIN(DSW_PWROK));
    defparam ipInertedIOPad_DSW_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DSW_PWROK_preio (
            .PADOEN(N__34175),
            .PADOUT(N__34174),
            .PADIN(N__34173),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24556),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5A_EN_iopad (
            .OE(N__34166),
            .DIN(N__34165),
            .DOUT(N__34164),
            .PACKAGEPIN(V5A_EN));
    defparam ipInertedIOPad_V5A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5A_EN_preio (
            .PADOEN(N__34166),
            .PADOUT(N__34165),
            .PADIN(N__34164),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24877),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_3_iopad (
            .OE(N__34157),
            .DIN(N__34156),
            .DOUT(N__34155),
            .PACKAGEPIN(GPIO_FPGA_SoC_3));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_3_preio (
            .PADOEN(N__34157),
            .PADOUT(N__34156),
            .PADIN(N__34155),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad (
            .OE(N__34148),
            .DIN(N__34147),
            .DOUT(N__34146),
            .PACKAGEPIN(VR_PROCHOT_FPGA_OUT_N));
    defparam ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio (
            .PADOEN(N__34148),
            .PADOUT(N__34147),
            .PADIN(N__34146),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VPP_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VPP_OK_iopad (
            .OE(N__34139),
            .DIN(N__34138),
            .DOUT(N__34137),
            .PACKAGEPIN(VPP_OK));
    defparam ipInertedIOPad_VPP_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VPP_OK_preio (
            .PADOEN(N__34139),
            .PADOUT(N__34138),
            .PADIN(N__34137),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vpp_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PE_iopad (
            .OE(N__34130),
            .DIN(N__34129),
            .DOUT(N__34128),
            .PACKAGEPIN(VCCIN_VR_PE));
    defparam ipInertedIOPad_VCCIN_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PE_preio (
            .PADOEN(N__34130),
            .PADOUT(N__34129),
            .PADIN(N__34128),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_EN_iopad (
            .OE(N__34121),
            .DIN(N__34120),
            .DOUT(N__34119),
            .PACKAGEPIN(VCCIN_EN));
    defparam ipInertedIOPad_VCCIN_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_EN_preio (
            .PADOEN(N__34121),
            .PADOUT(N__34120),
            .PADIN(N__34119),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24898),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SOC_SPKR_iopad (
            .OE(N__34112),
            .DIN(N__34111),
            .DOUT(N__34110),
            .PACKAGEPIN(SOC_SPKR));
    defparam ipInertedIOPad_SOC_SPKR_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SOC_SPKR_preio (
            .PADOEN(N__34112),
            .PADOUT(N__34111),
            .PADIN(N__34110),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S5n_iopad (
            .OE(N__34103),
            .DIN(N__34102),
            .DOUT(N__34101),
            .PACKAGEPIN(SLP_S5n));
    defparam ipInertedIOPad_SLP_S5n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S5n_preio (
            .PADOEN(N__34103),
            .PADOUT(N__34102),
            .PADIN(N__34101),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V12_MAIN_MON_iopad (
            .OE(N__34094),
            .DIN(N__34093),
            .DOUT(N__34092),
            .PACKAGEPIN(V12_MAIN_MON));
    defparam ipInertedIOPad_V12_MAIN_MON_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V12_MAIN_MON_preio (
            .PADOEN(N__34094),
            .PADOUT(N__34093),
            .PADIN(N__34092),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO3_iopad (
            .OE(N__34085),
            .DIN(N__34084),
            .DOUT(N__34083),
            .PACKAGEPIN(SPI_FP_IO3));
    defparam ipInertedIOPad_SPI_FP_IO3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO3_preio (
            .PADOEN(N__34085),
            .PADOUT(N__34084),
            .PADIN(N__34083),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE0_FPGA_iopad (
            .OE(N__34076),
            .DIN(N__34075),
            .DOUT(N__34074),
            .PACKAGEPIN(SATAXPCIE0_FPGA));
    defparam ipInertedIOPad_SATAXPCIE0_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE0_FPGA_preio (
            .PADOEN(N__34076),
            .PADOUT(N__34075),
            .PADIN(N__34074),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_OK_iopad (
            .OE(N__34067),
            .DIN(N__34066),
            .DOUT(N__34065),
            .PACKAGEPIN(V33A_OK));
    defparam ipInertedIOPad_V33A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33A_OK_preio (
            .PADOEN(N__34067),
            .PADOUT(N__34066),
            .PADIN(N__34065),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PCH_PWROK_iopad (
            .OE(N__34058),
            .DIN(N__34057),
            .DOUT(N__34056),
            .PACKAGEPIN(PCH_PWROK));
    defparam ipInertedIOPad_PCH_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PCH_PWROK_preio (
            .PADOEN(N__34058),
            .PADOUT(N__34057),
            .PADIN(N__34056),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20739),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_SLP_WLAN_N_iopad (
            .OE(N__34049),
            .DIN(N__34048),
            .DOUT(N__34047),
            .PACKAGEPIN(FPGA_SLP_WLAN_N));
    defparam ipInertedIOPad_FPGA_SLP_WLAN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_SLP_WLAN_N_preio (
            .PADOEN(N__34049),
            .PADOUT(N__34048),
            .PADIN(N__34047),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    CascadeMux I__7964 (
            .O(N__34030),
            .I(\VPP_VDDQ.N_178_cascade_ ));
    InMux I__7963 (
            .O(N__34027),
            .I(N__34011));
    InMux I__7962 (
            .O(N__34026),
            .I(N__34011));
    InMux I__7961 (
            .O(N__34025),
            .I(N__34011));
    InMux I__7960 (
            .O(N__34024),
            .I(N__34011));
    InMux I__7959 (
            .O(N__34023),
            .I(N__34004));
    InMux I__7958 (
            .O(N__34022),
            .I(N__34004));
    InMux I__7957 (
            .O(N__34021),
            .I(N__34004));
    CascadeMux I__7956 (
            .O(N__34020),
            .I(N__33995));
    LocalMux I__7955 (
            .O(N__34011),
            .I(N__33990));
    LocalMux I__7954 (
            .O(N__34004),
            .I(N__33990));
    InMux I__7953 (
            .O(N__34003),
            .I(N__33976));
    InMux I__7952 (
            .O(N__34002),
            .I(N__33976));
    InMux I__7951 (
            .O(N__34001),
            .I(N__33976));
    InMux I__7950 (
            .O(N__34000),
            .I(N__33973));
    CascadeMux I__7949 (
            .O(N__33999),
            .I(N__33970));
    InMux I__7948 (
            .O(N__33998),
            .I(N__33965));
    InMux I__7947 (
            .O(N__33995),
            .I(N__33965));
    Span4Mux_v I__7946 (
            .O(N__33990),
            .I(N__33962));
    InMux I__7945 (
            .O(N__33989),
            .I(N__33953));
    InMux I__7944 (
            .O(N__33988),
            .I(N__33953));
    InMux I__7943 (
            .O(N__33987),
            .I(N__33953));
    InMux I__7942 (
            .O(N__33986),
            .I(N__33953));
    InMux I__7941 (
            .O(N__33985),
            .I(N__33946));
    InMux I__7940 (
            .O(N__33984),
            .I(N__33946));
    InMux I__7939 (
            .O(N__33983),
            .I(N__33946));
    LocalMux I__7938 (
            .O(N__33976),
            .I(N__33934));
    LocalMux I__7937 (
            .O(N__33973),
            .I(N__33934));
    InMux I__7936 (
            .O(N__33970),
            .I(N__33925));
    LocalMux I__7935 (
            .O(N__33965),
            .I(N__33914));
    Sp12to4 I__7934 (
            .O(N__33962),
            .I(N__33914));
    LocalMux I__7933 (
            .O(N__33953),
            .I(N__33914));
    LocalMux I__7932 (
            .O(N__33946),
            .I(N__33914));
    InMux I__7931 (
            .O(N__33945),
            .I(N__33911));
    InMux I__7930 (
            .O(N__33944),
            .I(N__33902));
    InMux I__7929 (
            .O(N__33943),
            .I(N__33902));
    InMux I__7928 (
            .O(N__33942),
            .I(N__33902));
    InMux I__7927 (
            .O(N__33941),
            .I(N__33893));
    InMux I__7926 (
            .O(N__33940),
            .I(N__33893));
    InMux I__7925 (
            .O(N__33939),
            .I(N__33893));
    Span4Mux_v I__7924 (
            .O(N__33934),
            .I(N__33890));
    InMux I__7923 (
            .O(N__33933),
            .I(N__33887));
    IoInMux I__7922 (
            .O(N__33932),
            .I(N__33884));
    InMux I__7921 (
            .O(N__33931),
            .I(N__33881));
    InMux I__7920 (
            .O(N__33930),
            .I(N__33874));
    InMux I__7919 (
            .O(N__33929),
            .I(N__33871));
    InMux I__7918 (
            .O(N__33928),
            .I(N__33868));
    LocalMux I__7917 (
            .O(N__33925),
            .I(N__33865));
    InMux I__7916 (
            .O(N__33924),
            .I(N__33862));
    CascadeMux I__7915 (
            .O(N__33923),
            .I(N__33858));
    Span12Mux_s7_h I__7914 (
            .O(N__33914),
            .I(N__33855));
    LocalMux I__7913 (
            .O(N__33911),
            .I(N__33852));
    InMux I__7912 (
            .O(N__33910),
            .I(N__33844));
    InMux I__7911 (
            .O(N__33909),
            .I(N__33844));
    LocalMux I__7910 (
            .O(N__33902),
            .I(N__33841));
    InMux I__7909 (
            .O(N__33901),
            .I(N__33838));
    InMux I__7908 (
            .O(N__33900),
            .I(N__33835));
    LocalMux I__7907 (
            .O(N__33893),
            .I(N__33832));
    Span4Mux_v I__7906 (
            .O(N__33890),
            .I(N__33827));
    LocalMux I__7905 (
            .O(N__33887),
            .I(N__33827));
    LocalMux I__7904 (
            .O(N__33884),
            .I(N__33823));
    LocalMux I__7903 (
            .O(N__33881),
            .I(N__33820));
    InMux I__7902 (
            .O(N__33880),
            .I(N__33817));
    InMux I__7901 (
            .O(N__33879),
            .I(N__33810));
    InMux I__7900 (
            .O(N__33878),
            .I(N__33810));
    InMux I__7899 (
            .O(N__33877),
            .I(N__33810));
    LocalMux I__7898 (
            .O(N__33874),
            .I(N__33803));
    LocalMux I__7897 (
            .O(N__33871),
            .I(N__33803));
    LocalMux I__7896 (
            .O(N__33868),
            .I(N__33803));
    Span4Mux_v I__7895 (
            .O(N__33865),
            .I(N__33798));
    LocalMux I__7894 (
            .O(N__33862),
            .I(N__33798));
    InMux I__7893 (
            .O(N__33861),
            .I(N__33795));
    InMux I__7892 (
            .O(N__33858),
            .I(N__33792));
    Span12Mux_v I__7891 (
            .O(N__33855),
            .I(N__33789));
    Span12Mux_s10_h I__7890 (
            .O(N__33852),
            .I(N__33786));
    InMux I__7889 (
            .O(N__33851),
            .I(N__33779));
    InMux I__7888 (
            .O(N__33850),
            .I(N__33779));
    InMux I__7887 (
            .O(N__33849),
            .I(N__33779));
    LocalMux I__7886 (
            .O(N__33844),
            .I(N__33770));
    Span4Mux_s1_h I__7885 (
            .O(N__33841),
            .I(N__33770));
    LocalMux I__7884 (
            .O(N__33838),
            .I(N__33770));
    LocalMux I__7883 (
            .O(N__33835),
            .I(N__33770));
    Span4Mux_v I__7882 (
            .O(N__33832),
            .I(N__33765));
    Span4Mux_v I__7881 (
            .O(N__33827),
            .I(N__33765));
    InMux I__7880 (
            .O(N__33826),
            .I(N__33762));
    Span12Mux_s1_h I__7879 (
            .O(N__33823),
            .I(N__33751));
    Span12Mux_s10_h I__7878 (
            .O(N__33820),
            .I(N__33751));
    LocalMux I__7877 (
            .O(N__33817),
            .I(N__33751));
    LocalMux I__7876 (
            .O(N__33810),
            .I(N__33751));
    Span12Mux_s10_h I__7875 (
            .O(N__33803),
            .I(N__33751));
    Span4Mux_h I__7874 (
            .O(N__33798),
            .I(N__33748));
    LocalMux I__7873 (
            .O(N__33795),
            .I(suswarn_n));
    LocalMux I__7872 (
            .O(N__33792),
            .I(suswarn_n));
    Odrv12 I__7871 (
            .O(N__33789),
            .I(suswarn_n));
    Odrv12 I__7870 (
            .O(N__33786),
            .I(suswarn_n));
    LocalMux I__7869 (
            .O(N__33779),
            .I(suswarn_n));
    Odrv4 I__7868 (
            .O(N__33770),
            .I(suswarn_n));
    Odrv4 I__7867 (
            .O(N__33765),
            .I(suswarn_n));
    LocalMux I__7866 (
            .O(N__33762),
            .I(suswarn_n));
    Odrv12 I__7865 (
            .O(N__33751),
            .I(suswarn_n));
    Odrv4 I__7864 (
            .O(N__33748),
            .I(suswarn_n));
    CascadeMux I__7863 (
            .O(N__33727),
            .I(N__33711));
    CascadeMux I__7862 (
            .O(N__33726),
            .I(N__33707));
    CascadeMux I__7861 (
            .O(N__33725),
            .I(N__33702));
    InMux I__7860 (
            .O(N__33724),
            .I(N__33697));
    InMux I__7859 (
            .O(N__33723),
            .I(N__33694));
    CascadeMux I__7858 (
            .O(N__33722),
            .I(N__33691));
    CascadeMux I__7857 (
            .O(N__33721),
            .I(N__33688));
    CascadeMux I__7856 (
            .O(N__33720),
            .I(N__33685));
    CascadeMux I__7855 (
            .O(N__33719),
            .I(N__33681));
    CascadeMux I__7854 (
            .O(N__33718),
            .I(N__33678));
    InMux I__7853 (
            .O(N__33717),
            .I(N__33666));
    InMux I__7852 (
            .O(N__33716),
            .I(N__33666));
    InMux I__7851 (
            .O(N__33715),
            .I(N__33666));
    InMux I__7850 (
            .O(N__33714),
            .I(N__33666));
    InMux I__7849 (
            .O(N__33711),
            .I(N__33657));
    InMux I__7848 (
            .O(N__33710),
            .I(N__33657));
    InMux I__7847 (
            .O(N__33707),
            .I(N__33657));
    InMux I__7846 (
            .O(N__33706),
            .I(N__33657));
    CascadeMux I__7845 (
            .O(N__33705),
            .I(N__33651));
    InMux I__7844 (
            .O(N__33702),
            .I(N__33642));
    InMux I__7843 (
            .O(N__33701),
            .I(N__33642));
    InMux I__7842 (
            .O(N__33700),
            .I(N__33642));
    LocalMux I__7841 (
            .O(N__33697),
            .I(N__33637));
    LocalMux I__7840 (
            .O(N__33694),
            .I(N__33637));
    InMux I__7839 (
            .O(N__33691),
            .I(N__33634));
    InMux I__7838 (
            .O(N__33688),
            .I(N__33623));
    InMux I__7837 (
            .O(N__33685),
            .I(N__33623));
    InMux I__7836 (
            .O(N__33684),
            .I(N__33623));
    InMux I__7835 (
            .O(N__33681),
            .I(N__33623));
    InMux I__7834 (
            .O(N__33678),
            .I(N__33623));
    CascadeMux I__7833 (
            .O(N__33677),
            .I(N__33619));
    CascadeMux I__7832 (
            .O(N__33676),
            .I(N__33615));
    CascadeMux I__7831 (
            .O(N__33675),
            .I(N__33610));
    LocalMux I__7830 (
            .O(N__33666),
            .I(N__33603));
    LocalMux I__7829 (
            .O(N__33657),
            .I(N__33600));
    InMux I__7828 (
            .O(N__33656),
            .I(N__33587));
    InMux I__7827 (
            .O(N__33655),
            .I(N__33587));
    InMux I__7826 (
            .O(N__33654),
            .I(N__33587));
    InMux I__7825 (
            .O(N__33651),
            .I(N__33587));
    InMux I__7824 (
            .O(N__33650),
            .I(N__33587));
    InMux I__7823 (
            .O(N__33649),
            .I(N__33587));
    LocalMux I__7822 (
            .O(N__33642),
            .I(N__33584));
    Span4Mux_v I__7821 (
            .O(N__33637),
            .I(N__33581));
    LocalMux I__7820 (
            .O(N__33634),
            .I(N__33578));
    LocalMux I__7819 (
            .O(N__33623),
            .I(N__33575));
    InMux I__7818 (
            .O(N__33622),
            .I(N__33562));
    InMux I__7817 (
            .O(N__33619),
            .I(N__33562));
    InMux I__7816 (
            .O(N__33618),
            .I(N__33562));
    InMux I__7815 (
            .O(N__33615),
            .I(N__33562));
    InMux I__7814 (
            .O(N__33614),
            .I(N__33562));
    InMux I__7813 (
            .O(N__33613),
            .I(N__33562));
    InMux I__7812 (
            .O(N__33610),
            .I(N__33551));
    InMux I__7811 (
            .O(N__33609),
            .I(N__33551));
    InMux I__7810 (
            .O(N__33608),
            .I(N__33551));
    InMux I__7809 (
            .O(N__33607),
            .I(N__33551));
    InMux I__7808 (
            .O(N__33606),
            .I(N__33551));
    Span4Mux_s2_h I__7807 (
            .O(N__33603),
            .I(N__33548));
    Span4Mux_s2_h I__7806 (
            .O(N__33600),
            .I(N__33545));
    LocalMux I__7805 (
            .O(N__33587),
            .I(N__33540));
    Span4Mux_s2_h I__7804 (
            .O(N__33584),
            .I(N__33540));
    Odrv4 I__7803 (
            .O(N__33581),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv4 I__7802 (
            .O(N__33578),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv12 I__7801 (
            .O(N__33575),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7800 (
            .O(N__33562),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7799 (
            .O(N__33551),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv4 I__7798 (
            .O(N__33548),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv4 I__7797 (
            .O(N__33545),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv4 I__7796 (
            .O(N__33540),
            .I(\VPP_VDDQ.N_1_i ));
    CascadeMux I__7795 (
            .O(N__33523),
            .I(N__33514));
    CascadeMux I__7794 (
            .O(N__33522),
            .I(N__33506));
    CascadeMux I__7793 (
            .O(N__33521),
            .I(N__33503));
    InMux I__7792 (
            .O(N__33520),
            .I(N__33498));
    InMux I__7791 (
            .O(N__33519),
            .I(N__33498));
    CascadeMux I__7790 (
            .O(N__33518),
            .I(N__33485));
    CascadeMux I__7789 (
            .O(N__33517),
            .I(N__33482));
    InMux I__7788 (
            .O(N__33514),
            .I(N__33478));
    InMux I__7787 (
            .O(N__33513),
            .I(N__33475));
    InMux I__7786 (
            .O(N__33512),
            .I(N__33466));
    InMux I__7785 (
            .O(N__33511),
            .I(N__33466));
    InMux I__7784 (
            .O(N__33510),
            .I(N__33466));
    InMux I__7783 (
            .O(N__33509),
            .I(N__33466));
    InMux I__7782 (
            .O(N__33506),
            .I(N__33461));
    InMux I__7781 (
            .O(N__33503),
            .I(N__33461));
    LocalMux I__7780 (
            .O(N__33498),
            .I(N__33456));
    InMux I__7779 (
            .O(N__33497),
            .I(N__33453));
    CascadeMux I__7778 (
            .O(N__33496),
            .I(N__33449));
    InMux I__7777 (
            .O(N__33495),
            .I(N__33442));
    InMux I__7776 (
            .O(N__33494),
            .I(N__33442));
    InMux I__7775 (
            .O(N__33493),
            .I(N__33442));
    InMux I__7774 (
            .O(N__33492),
            .I(N__33437));
    InMux I__7773 (
            .O(N__33491),
            .I(N__33437));
    CascadeMux I__7772 (
            .O(N__33490),
            .I(N__33433));
    CascadeMux I__7771 (
            .O(N__33489),
            .I(N__33430));
    InMux I__7770 (
            .O(N__33488),
            .I(N__33418));
    InMux I__7769 (
            .O(N__33485),
            .I(N__33418));
    InMux I__7768 (
            .O(N__33482),
            .I(N__33418));
    InMux I__7767 (
            .O(N__33481),
            .I(N__33418));
    LocalMux I__7766 (
            .O(N__33478),
            .I(N__33409));
    LocalMux I__7765 (
            .O(N__33475),
            .I(N__33409));
    LocalMux I__7764 (
            .O(N__33466),
            .I(N__33409));
    LocalMux I__7763 (
            .O(N__33461),
            .I(N__33409));
    CascadeMux I__7762 (
            .O(N__33460),
            .I(N__33406));
    CascadeMux I__7761 (
            .O(N__33459),
            .I(N__33402));
    Span4Mux_s0_h I__7760 (
            .O(N__33456),
            .I(N__33396));
    LocalMux I__7759 (
            .O(N__33453),
            .I(N__33396));
    CascadeMux I__7758 (
            .O(N__33452),
            .I(N__33392));
    InMux I__7757 (
            .O(N__33449),
            .I(N__33388));
    LocalMux I__7756 (
            .O(N__33442),
            .I(N__33383));
    LocalMux I__7755 (
            .O(N__33437),
            .I(N__33383));
    InMux I__7754 (
            .O(N__33436),
            .I(N__33370));
    InMux I__7753 (
            .O(N__33433),
            .I(N__33370));
    InMux I__7752 (
            .O(N__33430),
            .I(N__33370));
    InMux I__7751 (
            .O(N__33429),
            .I(N__33370));
    InMux I__7750 (
            .O(N__33428),
            .I(N__33370));
    InMux I__7749 (
            .O(N__33427),
            .I(N__33370));
    LocalMux I__7748 (
            .O(N__33418),
            .I(N__33367));
    Span4Mux_v I__7747 (
            .O(N__33409),
            .I(N__33360));
    InMux I__7746 (
            .O(N__33406),
            .I(N__33351));
    InMux I__7745 (
            .O(N__33405),
            .I(N__33351));
    InMux I__7744 (
            .O(N__33402),
            .I(N__33351));
    InMux I__7743 (
            .O(N__33401),
            .I(N__33351));
    Span4Mux_v I__7742 (
            .O(N__33396),
            .I(N__33348));
    InMux I__7741 (
            .O(N__33395),
            .I(N__33345));
    InMux I__7740 (
            .O(N__33392),
            .I(N__33340));
    InMux I__7739 (
            .O(N__33391),
            .I(N__33340));
    LocalMux I__7738 (
            .O(N__33388),
            .I(N__33333));
    Span4Mux_s1_v I__7737 (
            .O(N__33383),
            .I(N__33333));
    LocalMux I__7736 (
            .O(N__33370),
            .I(N__33333));
    Span4Mux_h I__7735 (
            .O(N__33367),
            .I(N__33330));
    InMux I__7734 (
            .O(N__33366),
            .I(N__33321));
    InMux I__7733 (
            .O(N__33365),
            .I(N__33321));
    InMux I__7732 (
            .O(N__33364),
            .I(N__33321));
    InMux I__7731 (
            .O(N__33363),
            .I(N__33321));
    Span4Mux_h I__7730 (
            .O(N__33360),
            .I(N__33314));
    LocalMux I__7729 (
            .O(N__33351),
            .I(N__33314));
    Span4Mux_v I__7728 (
            .O(N__33348),
            .I(N__33314));
    LocalMux I__7727 (
            .O(N__33345),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__7726 (
            .O(N__33340),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    Odrv4 I__7725 (
            .O(N__33333),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    Odrv4 I__7724 (
            .O(N__33330),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__7723 (
            .O(N__33321),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    Odrv4 I__7722 (
            .O(N__33314),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    CascadeMux I__7721 (
            .O(N__33301),
            .I(N__33291));
    InMux I__7720 (
            .O(N__33300),
            .I(N__33270));
    InMux I__7719 (
            .O(N__33299),
            .I(N__33270));
    InMux I__7718 (
            .O(N__33298),
            .I(N__33270));
    InMux I__7717 (
            .O(N__33297),
            .I(N__33270));
    InMux I__7716 (
            .O(N__33296),
            .I(N__33270));
    InMux I__7715 (
            .O(N__33295),
            .I(N__33261));
    InMux I__7714 (
            .O(N__33294),
            .I(N__33248));
    InMux I__7713 (
            .O(N__33291),
            .I(N__33248));
    InMux I__7712 (
            .O(N__33290),
            .I(N__33248));
    InMux I__7711 (
            .O(N__33289),
            .I(N__33248));
    InMux I__7710 (
            .O(N__33288),
            .I(N__33248));
    InMux I__7709 (
            .O(N__33287),
            .I(N__33248));
    InMux I__7708 (
            .O(N__33286),
            .I(N__33237));
    InMux I__7707 (
            .O(N__33285),
            .I(N__33237));
    InMux I__7706 (
            .O(N__33284),
            .I(N__33237));
    InMux I__7705 (
            .O(N__33283),
            .I(N__33237));
    InMux I__7704 (
            .O(N__33282),
            .I(N__33237));
    CascadeMux I__7703 (
            .O(N__33281),
            .I(N__33227));
    LocalMux I__7702 (
            .O(N__33270),
            .I(N__33224));
    InMux I__7701 (
            .O(N__33269),
            .I(N__33211));
    InMux I__7700 (
            .O(N__33268),
            .I(N__33211));
    InMux I__7699 (
            .O(N__33267),
            .I(N__33211));
    InMux I__7698 (
            .O(N__33266),
            .I(N__33211));
    InMux I__7697 (
            .O(N__33265),
            .I(N__33211));
    InMux I__7696 (
            .O(N__33264),
            .I(N__33211));
    LocalMux I__7695 (
            .O(N__33261),
            .I(N__33204));
    LocalMux I__7694 (
            .O(N__33248),
            .I(N__33204));
    LocalMux I__7693 (
            .O(N__33237),
            .I(N__33204));
    InMux I__7692 (
            .O(N__33236),
            .I(N__33192));
    InMux I__7691 (
            .O(N__33235),
            .I(N__33192));
    InMux I__7690 (
            .O(N__33234),
            .I(N__33192));
    InMux I__7689 (
            .O(N__33233),
            .I(N__33192));
    InMux I__7688 (
            .O(N__33232),
            .I(N__33189));
    CascadeMux I__7687 (
            .O(N__33231),
            .I(N__33185));
    InMux I__7686 (
            .O(N__33230),
            .I(N__33180));
    InMux I__7685 (
            .O(N__33227),
            .I(N__33177));
    Span4Mux_s1_v I__7684 (
            .O(N__33224),
            .I(N__33170));
    LocalMux I__7683 (
            .O(N__33211),
            .I(N__33170));
    Span4Mux_v I__7682 (
            .O(N__33204),
            .I(N__33170));
    InMux I__7681 (
            .O(N__33203),
            .I(N__33163));
    InMux I__7680 (
            .O(N__33202),
            .I(N__33163));
    InMux I__7679 (
            .O(N__33201),
            .I(N__33163));
    LocalMux I__7678 (
            .O(N__33192),
            .I(N__33158));
    LocalMux I__7677 (
            .O(N__33189),
            .I(N__33158));
    InMux I__7676 (
            .O(N__33188),
            .I(N__33149));
    InMux I__7675 (
            .O(N__33185),
            .I(N__33149));
    InMux I__7674 (
            .O(N__33184),
            .I(N__33149));
    InMux I__7673 (
            .O(N__33183),
            .I(N__33149));
    LocalMux I__7672 (
            .O(N__33180),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    LocalMux I__7671 (
            .O(N__33177),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    Odrv4 I__7670 (
            .O(N__33170),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    LocalMux I__7669 (
            .O(N__33163),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    Odrv4 I__7668 (
            .O(N__33158),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    LocalMux I__7667 (
            .O(N__33149),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    InMux I__7666 (
            .O(N__33136),
            .I(N__33128));
    InMux I__7665 (
            .O(N__33135),
            .I(N__33128));
    InMux I__7664 (
            .O(N__33134),
            .I(N__33123));
    InMux I__7663 (
            .O(N__33133),
            .I(N__33123));
    LocalMux I__7662 (
            .O(N__33128),
            .I(N__33117));
    LocalMux I__7661 (
            .O(N__33123),
            .I(N__33117));
    InMux I__7660 (
            .O(N__33122),
            .I(N__33111));
    Span4Mux_v I__7659 (
            .O(N__33117),
            .I(N__33108));
    InMux I__7658 (
            .O(N__33116),
            .I(N__33105));
    InMux I__7657 (
            .O(N__33115),
            .I(N__33100));
    InMux I__7656 (
            .O(N__33114),
            .I(N__33100));
    LocalMux I__7655 (
            .O(N__33111),
            .I(N__33097));
    Span4Mux_v I__7654 (
            .O(N__33108),
            .I(N__33094));
    LocalMux I__7653 (
            .O(N__33105),
            .I(N__33089));
    LocalMux I__7652 (
            .O(N__33100),
            .I(N__33089));
    Span4Mux_s2_v I__7651 (
            .O(N__33097),
            .I(N__33085));
    Span4Mux_v I__7650 (
            .O(N__33094),
            .I(N__33080));
    Span4Mux_s2_v I__7649 (
            .O(N__33089),
            .I(N__33080));
    InMux I__7648 (
            .O(N__33088),
            .I(N__33077));
    Odrv4 I__7647 (
            .O(N__33085),
            .I(vddq_ok));
    Odrv4 I__7646 (
            .O(N__33080),
            .I(vddq_ok));
    LocalMux I__7645 (
            .O(N__33077),
            .I(vddq_ok));
    InMux I__7644 (
            .O(N__33070),
            .I(N__33067));
    LocalMux I__7643 (
            .O(N__33067),
            .I(\VPP_VDDQ.curr_state_2_0_1 ));
    ClkMux I__7642 (
            .O(N__33064),
            .I(N__33061));
    LocalMux I__7641 (
            .O(N__33061),
            .I(N__33055));
    ClkMux I__7640 (
            .O(N__33060),
            .I(N__33052));
    ClkMux I__7639 (
            .O(N__33059),
            .I(N__33049));
    ClkMux I__7638 (
            .O(N__33058),
            .I(N__33046));
    Span4Mux_s3_v I__7637 (
            .O(N__33055),
            .I(N__33032));
    LocalMux I__7636 (
            .O(N__33052),
            .I(N__33032));
    LocalMux I__7635 (
            .O(N__33049),
            .I(N__33027));
    LocalMux I__7634 (
            .O(N__33046),
            .I(N__33027));
    ClkMux I__7633 (
            .O(N__33045),
            .I(N__33024));
    ClkMux I__7632 (
            .O(N__33044),
            .I(N__33019));
    ClkMux I__7631 (
            .O(N__33043),
            .I(N__33012));
    ClkMux I__7630 (
            .O(N__33042),
            .I(N__33009));
    ClkMux I__7629 (
            .O(N__33041),
            .I(N__33006));
    ClkMux I__7628 (
            .O(N__33040),
            .I(N__33003));
    ClkMux I__7627 (
            .O(N__33039),
            .I(N__33000));
    ClkMux I__7626 (
            .O(N__33038),
            .I(N__32996));
    ClkMux I__7625 (
            .O(N__33037),
            .I(N__32991));
    Span4Mux_h I__7624 (
            .O(N__33032),
            .I(N__32983));
    Span4Mux_s3_v I__7623 (
            .O(N__33027),
            .I(N__32983));
    LocalMux I__7622 (
            .O(N__33024),
            .I(N__32983));
    ClkMux I__7621 (
            .O(N__33023),
            .I(N__32980));
    ClkMux I__7620 (
            .O(N__33022),
            .I(N__32975));
    LocalMux I__7619 (
            .O(N__33019),
            .I(N__32968));
    ClkMux I__7618 (
            .O(N__33018),
            .I(N__32965));
    ClkMux I__7617 (
            .O(N__33017),
            .I(N__32958));
    ClkMux I__7616 (
            .O(N__33016),
            .I(N__32954));
    ClkMux I__7615 (
            .O(N__33015),
            .I(N__32951));
    LocalMux I__7614 (
            .O(N__33012),
            .I(N__32948));
    LocalMux I__7613 (
            .O(N__33009),
            .I(N__32943));
    LocalMux I__7612 (
            .O(N__33006),
            .I(N__32943));
    LocalMux I__7611 (
            .O(N__33003),
            .I(N__32938));
    LocalMux I__7610 (
            .O(N__33000),
            .I(N__32935));
    ClkMux I__7609 (
            .O(N__32999),
            .I(N__32932));
    LocalMux I__7608 (
            .O(N__32996),
            .I(N__32928));
    ClkMux I__7607 (
            .O(N__32995),
            .I(N__32925));
    ClkMux I__7606 (
            .O(N__32994),
            .I(N__32922));
    LocalMux I__7605 (
            .O(N__32991),
            .I(N__32918));
    ClkMux I__7604 (
            .O(N__32990),
            .I(N__32915));
    Span4Mux_v I__7603 (
            .O(N__32983),
            .I(N__32910));
    LocalMux I__7602 (
            .O(N__32980),
            .I(N__32910));
    ClkMux I__7601 (
            .O(N__32979),
            .I(N__32907));
    ClkMux I__7600 (
            .O(N__32978),
            .I(N__32904));
    LocalMux I__7599 (
            .O(N__32975),
            .I(N__32898));
    ClkMux I__7598 (
            .O(N__32974),
            .I(N__32895));
    ClkMux I__7597 (
            .O(N__32973),
            .I(N__32892));
    ClkMux I__7596 (
            .O(N__32972),
            .I(N__32889));
    ClkMux I__7595 (
            .O(N__32971),
            .I(N__32886));
    Span4Mux_v I__7594 (
            .O(N__32968),
            .I(N__32879));
    LocalMux I__7593 (
            .O(N__32965),
            .I(N__32879));
    ClkMux I__7592 (
            .O(N__32964),
            .I(N__32876));
    ClkMux I__7591 (
            .O(N__32963),
            .I(N__32871));
    ClkMux I__7590 (
            .O(N__32962),
            .I(N__32867));
    ClkMux I__7589 (
            .O(N__32961),
            .I(N__32864));
    LocalMux I__7588 (
            .O(N__32958),
            .I(N__32861));
    ClkMux I__7587 (
            .O(N__32957),
            .I(N__32858));
    LocalMux I__7586 (
            .O(N__32954),
            .I(N__32852));
    LocalMux I__7585 (
            .O(N__32951),
            .I(N__32852));
    Span4Mux_h I__7584 (
            .O(N__32948),
            .I(N__32847));
    Span4Mux_v I__7583 (
            .O(N__32943),
            .I(N__32847));
    ClkMux I__7582 (
            .O(N__32942),
            .I(N__32844));
    ClkMux I__7581 (
            .O(N__32941),
            .I(N__32840));
    Span4Mux_s3_v I__7580 (
            .O(N__32938),
            .I(N__32832));
    Span4Mux_s3_v I__7579 (
            .O(N__32935),
            .I(N__32832));
    LocalMux I__7578 (
            .O(N__32932),
            .I(N__32832));
    ClkMux I__7577 (
            .O(N__32931),
            .I(N__32829));
    Span4Mux_s3_h I__7576 (
            .O(N__32928),
            .I(N__32822));
    LocalMux I__7575 (
            .O(N__32925),
            .I(N__32822));
    LocalMux I__7574 (
            .O(N__32922),
            .I(N__32822));
    ClkMux I__7573 (
            .O(N__32921),
            .I(N__32819));
    Span4Mux_v I__7572 (
            .O(N__32918),
            .I(N__32812));
    LocalMux I__7571 (
            .O(N__32915),
            .I(N__32812));
    Span4Mux_h I__7570 (
            .O(N__32910),
            .I(N__32807));
    LocalMux I__7569 (
            .O(N__32907),
            .I(N__32807));
    LocalMux I__7568 (
            .O(N__32904),
            .I(N__32804));
    ClkMux I__7567 (
            .O(N__32903),
            .I(N__32801));
    ClkMux I__7566 (
            .O(N__32902),
            .I(N__32797));
    ClkMux I__7565 (
            .O(N__32901),
            .I(N__32794));
    Span4Mux_h I__7564 (
            .O(N__32898),
            .I(N__32789));
    LocalMux I__7563 (
            .O(N__32895),
            .I(N__32789));
    LocalMux I__7562 (
            .O(N__32892),
            .I(N__32786));
    LocalMux I__7561 (
            .O(N__32889),
            .I(N__32781));
    LocalMux I__7560 (
            .O(N__32886),
            .I(N__32781));
    ClkMux I__7559 (
            .O(N__32885),
            .I(N__32778));
    ClkMux I__7558 (
            .O(N__32884),
            .I(N__32775));
    Span4Mux_v I__7557 (
            .O(N__32879),
            .I(N__32770));
    LocalMux I__7556 (
            .O(N__32876),
            .I(N__32770));
    ClkMux I__7555 (
            .O(N__32875),
            .I(N__32767));
    ClkMux I__7554 (
            .O(N__32874),
            .I(N__32763));
    LocalMux I__7553 (
            .O(N__32871),
            .I(N__32759));
    ClkMux I__7552 (
            .O(N__32870),
            .I(N__32756));
    LocalMux I__7551 (
            .O(N__32867),
            .I(N__32748));
    LocalMux I__7550 (
            .O(N__32864),
            .I(N__32744));
    Span4Mux_s3_v I__7549 (
            .O(N__32861),
            .I(N__32739));
    LocalMux I__7548 (
            .O(N__32858),
            .I(N__32739));
    ClkMux I__7547 (
            .O(N__32857),
            .I(N__32736));
    Span4Mux_v I__7546 (
            .O(N__32852),
            .I(N__32732));
    Span4Mux_v I__7545 (
            .O(N__32847),
            .I(N__32727));
    LocalMux I__7544 (
            .O(N__32844),
            .I(N__32727));
    ClkMux I__7543 (
            .O(N__32843),
            .I(N__32723));
    LocalMux I__7542 (
            .O(N__32840),
            .I(N__32720));
    ClkMux I__7541 (
            .O(N__32839),
            .I(N__32717));
    Span4Mux_v I__7540 (
            .O(N__32832),
            .I(N__32709));
    LocalMux I__7539 (
            .O(N__32829),
            .I(N__32709));
    Span4Mux_v I__7538 (
            .O(N__32822),
            .I(N__32704));
    LocalMux I__7537 (
            .O(N__32819),
            .I(N__32704));
    ClkMux I__7536 (
            .O(N__32818),
            .I(N__32701));
    ClkMux I__7535 (
            .O(N__32817),
            .I(N__32698));
    Span4Mux_v I__7534 (
            .O(N__32812),
            .I(N__32689));
    Span4Mux_v I__7533 (
            .O(N__32807),
            .I(N__32689));
    Span4Mux_h I__7532 (
            .O(N__32804),
            .I(N__32689));
    LocalMux I__7531 (
            .O(N__32801),
            .I(N__32689));
    ClkMux I__7530 (
            .O(N__32800),
            .I(N__32686));
    LocalMux I__7529 (
            .O(N__32797),
            .I(N__32681));
    LocalMux I__7528 (
            .O(N__32794),
            .I(N__32681));
    Span4Mux_v I__7527 (
            .O(N__32789),
            .I(N__32672));
    Span4Mux_h I__7526 (
            .O(N__32786),
            .I(N__32672));
    Span4Mux_v I__7525 (
            .O(N__32781),
            .I(N__32672));
    LocalMux I__7524 (
            .O(N__32778),
            .I(N__32672));
    LocalMux I__7523 (
            .O(N__32775),
            .I(N__32669));
    Span4Mux_v I__7522 (
            .O(N__32770),
            .I(N__32664));
    LocalMux I__7521 (
            .O(N__32767),
            .I(N__32664));
    ClkMux I__7520 (
            .O(N__32766),
            .I(N__32661));
    LocalMux I__7519 (
            .O(N__32763),
            .I(N__32656));
    ClkMux I__7518 (
            .O(N__32762),
            .I(N__32653));
    Span4Mux_s2_h I__7517 (
            .O(N__32759),
            .I(N__32647));
    LocalMux I__7516 (
            .O(N__32756),
            .I(N__32644));
    ClkMux I__7515 (
            .O(N__32755),
            .I(N__32641));
    ClkMux I__7514 (
            .O(N__32754),
            .I(N__32638));
    ClkMux I__7513 (
            .O(N__32753),
            .I(N__32634));
    ClkMux I__7512 (
            .O(N__32752),
            .I(N__32631));
    ClkMux I__7511 (
            .O(N__32751),
            .I(N__32626));
    Span4Mux_v I__7510 (
            .O(N__32748),
            .I(N__32623));
    ClkMux I__7509 (
            .O(N__32747),
            .I(N__32620));
    Span4Mux_v I__7508 (
            .O(N__32744),
            .I(N__32617));
    Span4Mux_v I__7507 (
            .O(N__32739),
            .I(N__32612));
    LocalMux I__7506 (
            .O(N__32736),
            .I(N__32612));
    ClkMux I__7505 (
            .O(N__32735),
            .I(N__32609));
    Span4Mux_v I__7504 (
            .O(N__32732),
            .I(N__32606));
    Span4Mux_h I__7503 (
            .O(N__32727),
            .I(N__32603));
    ClkMux I__7502 (
            .O(N__32726),
            .I(N__32600));
    LocalMux I__7501 (
            .O(N__32723),
            .I(N__32597));
    Span4Mux_v I__7500 (
            .O(N__32720),
            .I(N__32592));
    LocalMux I__7499 (
            .O(N__32717),
            .I(N__32592));
    ClkMux I__7498 (
            .O(N__32716),
            .I(N__32589));
    ClkMux I__7497 (
            .O(N__32715),
            .I(N__32586));
    ClkMux I__7496 (
            .O(N__32714),
            .I(N__32583));
    Span4Mux_v I__7495 (
            .O(N__32709),
            .I(N__32576));
    Span4Mux_v I__7494 (
            .O(N__32704),
            .I(N__32576));
    LocalMux I__7493 (
            .O(N__32701),
            .I(N__32576));
    LocalMux I__7492 (
            .O(N__32698),
            .I(N__32573));
    Span4Mux_v I__7491 (
            .O(N__32689),
            .I(N__32568));
    LocalMux I__7490 (
            .O(N__32686),
            .I(N__32568));
    Span4Mux_v I__7489 (
            .O(N__32681),
            .I(N__32565));
    Span4Mux_v I__7488 (
            .O(N__32672),
            .I(N__32556));
    Span4Mux_h I__7487 (
            .O(N__32669),
            .I(N__32556));
    Span4Mux_h I__7486 (
            .O(N__32664),
            .I(N__32556));
    LocalMux I__7485 (
            .O(N__32661),
            .I(N__32556));
    ClkMux I__7484 (
            .O(N__32660),
            .I(N__32553));
    ClkMux I__7483 (
            .O(N__32659),
            .I(N__32550));
    Span4Mux_s2_h I__7482 (
            .O(N__32656),
            .I(N__32546));
    LocalMux I__7481 (
            .O(N__32653),
            .I(N__32543));
    ClkMux I__7480 (
            .O(N__32652),
            .I(N__32540));
    ClkMux I__7479 (
            .O(N__32651),
            .I(N__32537));
    ClkMux I__7478 (
            .O(N__32650),
            .I(N__32532));
    Span4Mux_h I__7477 (
            .O(N__32647),
            .I(N__32523));
    Span4Mux_s1_v I__7476 (
            .O(N__32644),
            .I(N__32523));
    LocalMux I__7475 (
            .O(N__32641),
            .I(N__32523));
    LocalMux I__7474 (
            .O(N__32638),
            .I(N__32523));
    ClkMux I__7473 (
            .O(N__32637),
            .I(N__32520));
    LocalMux I__7472 (
            .O(N__32634),
            .I(N__32515));
    LocalMux I__7471 (
            .O(N__32631),
            .I(N__32515));
    ClkMux I__7470 (
            .O(N__32630),
            .I(N__32512));
    ClkMux I__7469 (
            .O(N__32629),
            .I(N__32509));
    LocalMux I__7468 (
            .O(N__32626),
            .I(N__32504));
    Span4Mux_v I__7467 (
            .O(N__32623),
            .I(N__32499));
    LocalMux I__7466 (
            .O(N__32620),
            .I(N__32499));
    Span4Mux_v I__7465 (
            .O(N__32617),
            .I(N__32494));
    Span4Mux_v I__7464 (
            .O(N__32612),
            .I(N__32494));
    LocalMux I__7463 (
            .O(N__32609),
            .I(N__32491));
    Span4Mux_v I__7462 (
            .O(N__32606),
            .I(N__32488));
    Span4Mux_v I__7461 (
            .O(N__32603),
            .I(N__32483));
    LocalMux I__7460 (
            .O(N__32600),
            .I(N__32483));
    Span4Mux_v I__7459 (
            .O(N__32597),
            .I(N__32476));
    Span4Mux_v I__7458 (
            .O(N__32592),
            .I(N__32476));
    LocalMux I__7457 (
            .O(N__32589),
            .I(N__32476));
    LocalMux I__7456 (
            .O(N__32586),
            .I(N__32471));
    LocalMux I__7455 (
            .O(N__32583),
            .I(N__32471));
    Span4Mux_v I__7454 (
            .O(N__32576),
            .I(N__32464));
    Span4Mux_h I__7453 (
            .O(N__32573),
            .I(N__32464));
    Span4Mux_h I__7452 (
            .O(N__32568),
            .I(N__32464));
    Span4Mux_h I__7451 (
            .O(N__32565),
            .I(N__32455));
    Span4Mux_v I__7450 (
            .O(N__32556),
            .I(N__32455));
    LocalMux I__7449 (
            .O(N__32553),
            .I(N__32455));
    LocalMux I__7448 (
            .O(N__32550),
            .I(N__32455));
    ClkMux I__7447 (
            .O(N__32549),
            .I(N__32452));
    Span4Mux_v I__7446 (
            .O(N__32546),
            .I(N__32445));
    Span4Mux_s2_h I__7445 (
            .O(N__32543),
            .I(N__32445));
    LocalMux I__7444 (
            .O(N__32540),
            .I(N__32445));
    LocalMux I__7443 (
            .O(N__32537),
            .I(N__32442));
    ClkMux I__7442 (
            .O(N__32536),
            .I(N__32439));
    ClkMux I__7441 (
            .O(N__32535),
            .I(N__32436));
    LocalMux I__7440 (
            .O(N__32532),
            .I(N__32429));
    Span4Mux_v I__7439 (
            .O(N__32523),
            .I(N__32429));
    LocalMux I__7438 (
            .O(N__32520),
            .I(N__32429));
    Span4Mux_v I__7437 (
            .O(N__32515),
            .I(N__32422));
    LocalMux I__7436 (
            .O(N__32512),
            .I(N__32422));
    LocalMux I__7435 (
            .O(N__32509),
            .I(N__32422));
    ClkMux I__7434 (
            .O(N__32508),
            .I(N__32419));
    ClkMux I__7433 (
            .O(N__32507),
            .I(N__32415));
    Span4Mux_v I__7432 (
            .O(N__32504),
            .I(N__32410));
    Span4Mux_v I__7431 (
            .O(N__32499),
            .I(N__32410));
    Span4Mux_v I__7430 (
            .O(N__32494),
            .I(N__32405));
    Span4Mux_v I__7429 (
            .O(N__32491),
            .I(N__32405));
    IoSpan4Mux I__7428 (
            .O(N__32488),
            .I(N__32400));
    IoSpan4Mux I__7427 (
            .O(N__32483),
            .I(N__32400));
    Span4Mux_v I__7426 (
            .O(N__32476),
            .I(N__32395));
    Span4Mux_v I__7425 (
            .O(N__32471),
            .I(N__32395));
    Span4Mux_h I__7424 (
            .O(N__32464),
            .I(N__32388));
    IoSpan4Mux I__7423 (
            .O(N__32455),
            .I(N__32388));
    LocalMux I__7422 (
            .O(N__32452),
            .I(N__32388));
    Span4Mux_v I__7421 (
            .O(N__32445),
            .I(N__32379));
    Span4Mux_s2_h I__7420 (
            .O(N__32442),
            .I(N__32379));
    LocalMux I__7419 (
            .O(N__32439),
            .I(N__32379));
    LocalMux I__7418 (
            .O(N__32436),
            .I(N__32379));
    Span4Mux_v I__7417 (
            .O(N__32429),
            .I(N__32372));
    Span4Mux_v I__7416 (
            .O(N__32422),
            .I(N__32372));
    LocalMux I__7415 (
            .O(N__32419),
            .I(N__32372));
    ClkMux I__7414 (
            .O(N__32418),
            .I(N__32369));
    LocalMux I__7413 (
            .O(N__32415),
            .I(N__32364));
    IoSpan4Mux I__7412 (
            .O(N__32410),
            .I(N__32359));
    IoSpan4Mux I__7411 (
            .O(N__32405),
            .I(N__32359));
    IoSpan4Mux I__7410 (
            .O(N__32400),
            .I(N__32352));
    IoSpan4Mux I__7409 (
            .O(N__32395),
            .I(N__32352));
    IoSpan4Mux I__7408 (
            .O(N__32388),
            .I(N__32352));
    Span4Mux_h I__7407 (
            .O(N__32379),
            .I(N__32349));
    Span4Mux_v I__7406 (
            .O(N__32372),
            .I(N__32344));
    LocalMux I__7405 (
            .O(N__32369),
            .I(N__32344));
    ClkMux I__7404 (
            .O(N__32368),
            .I(N__32341));
    ClkMux I__7403 (
            .O(N__32367),
            .I(N__32338));
    Odrv12 I__7402 (
            .O(N__32364),
            .I(fpga_osc));
    Odrv4 I__7401 (
            .O(N__32359),
            .I(fpga_osc));
    Odrv4 I__7400 (
            .O(N__32352),
            .I(fpga_osc));
    Odrv4 I__7399 (
            .O(N__32349),
            .I(fpga_osc));
    Odrv4 I__7398 (
            .O(N__32344),
            .I(fpga_osc));
    LocalMux I__7397 (
            .O(N__32341),
            .I(fpga_osc));
    LocalMux I__7396 (
            .O(N__32338),
            .I(fpga_osc));
    CascadeMux I__7395 (
            .O(N__32323),
            .I(N__32320));
    InMux I__7394 (
            .O(N__32320),
            .I(N__32311));
    InMux I__7393 (
            .O(N__32319),
            .I(N__32308));
    InMux I__7392 (
            .O(N__32318),
            .I(N__32305));
    InMux I__7391 (
            .O(N__32317),
            .I(N__32302));
    InMux I__7390 (
            .O(N__32316),
            .I(N__32299));
    InMux I__7389 (
            .O(N__32315),
            .I(N__32296));
    InMux I__7388 (
            .O(N__32314),
            .I(N__32293));
    LocalMux I__7387 (
            .O(N__32311),
            .I(N__32281));
    LocalMux I__7386 (
            .O(N__32308),
            .I(N__32278));
    LocalMux I__7385 (
            .O(N__32305),
            .I(N__32275));
    LocalMux I__7384 (
            .O(N__32302),
            .I(N__32272));
    LocalMux I__7383 (
            .O(N__32299),
            .I(N__32269));
    LocalMux I__7382 (
            .O(N__32296),
            .I(N__32266));
    LocalMux I__7381 (
            .O(N__32293),
            .I(N__32263));
    CEMux I__7380 (
            .O(N__32292),
            .I(N__32230));
    CEMux I__7379 (
            .O(N__32291),
            .I(N__32230));
    CEMux I__7378 (
            .O(N__32290),
            .I(N__32230));
    CEMux I__7377 (
            .O(N__32289),
            .I(N__32230));
    CEMux I__7376 (
            .O(N__32288),
            .I(N__32230));
    CEMux I__7375 (
            .O(N__32287),
            .I(N__32230));
    CEMux I__7374 (
            .O(N__32286),
            .I(N__32230));
    CEMux I__7373 (
            .O(N__32285),
            .I(N__32230));
    CEMux I__7372 (
            .O(N__32284),
            .I(N__32230));
    Glb2LocalMux I__7371 (
            .O(N__32281),
            .I(N__32230));
    Glb2LocalMux I__7370 (
            .O(N__32278),
            .I(N__32230));
    Glb2LocalMux I__7369 (
            .O(N__32275),
            .I(N__32230));
    Glb2LocalMux I__7368 (
            .O(N__32272),
            .I(N__32230));
    Glb2LocalMux I__7367 (
            .O(N__32269),
            .I(N__32230));
    Glb2LocalMux I__7366 (
            .O(N__32266),
            .I(N__32230));
    Glb2LocalMux I__7365 (
            .O(N__32263),
            .I(N__32230));
    GlobalMux I__7364 (
            .O(N__32230),
            .I(N__32227));
    gio2CtrlBuf I__7363 (
            .O(N__32227),
            .I(N_587_g));
    InMux I__7362 (
            .O(N__32224),
            .I(N__32218));
    InMux I__7361 (
            .O(N__32223),
            .I(N__32218));
    LocalMux I__7360 (
            .O(N__32218),
            .I(\VPP_VDDQ.count_2Z0Z_7 ));
    InMux I__7359 (
            .O(N__32215),
            .I(N__32212));
    LocalMux I__7358 (
            .O(N__32212),
            .I(\VPP_VDDQ.count_2_1_7 ));
    InMux I__7357 (
            .O(N__32209),
            .I(N__32206));
    LocalMux I__7356 (
            .O(N__32206),
            .I(N__32203));
    Odrv4 I__7355 (
            .O(N__32203),
            .I(\VPP_VDDQ.un1_count_2_1_axb_7 ));
    CascadeMux I__7354 (
            .O(N__32200),
            .I(\VPP_VDDQ.count_2_RNIZ0Z_1_cascade_ ));
    CascadeMux I__7353 (
            .O(N__32197),
            .I(\VPP_VDDQ.count_2_1_1_cascade_ ));
    InMux I__7352 (
            .O(N__32194),
            .I(N__32191));
    LocalMux I__7351 (
            .O(N__32191),
            .I(N__32187));
    InMux I__7350 (
            .O(N__32190),
            .I(N__32184));
    Span4Mux_h I__7349 (
            .O(N__32187),
            .I(N__32181));
    LocalMux I__7348 (
            .O(N__32184),
            .I(\VPP_VDDQ.un1_count_2_1_axb_1 ));
    Odrv4 I__7347 (
            .O(N__32181),
            .I(\VPP_VDDQ.un1_count_2_1_axb_1 ));
    InMux I__7346 (
            .O(N__32176),
            .I(N__32173));
    LocalMux I__7345 (
            .O(N__32173),
            .I(\VPP_VDDQ.count_2_1_1 ));
    CascadeMux I__7344 (
            .O(N__32170),
            .I(N__32165));
    CascadeMux I__7343 (
            .O(N__32169),
            .I(N__32162));
    CascadeMux I__7342 (
            .O(N__32168),
            .I(N__32159));
    InMux I__7341 (
            .O(N__32165),
            .I(N__32155));
    InMux I__7340 (
            .O(N__32162),
            .I(N__32152));
    InMux I__7339 (
            .O(N__32159),
            .I(N__32147));
    InMux I__7338 (
            .O(N__32158),
            .I(N__32147));
    LocalMux I__7337 (
            .O(N__32155),
            .I(N__32144));
    LocalMux I__7336 (
            .O(N__32152),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    LocalMux I__7335 (
            .O(N__32147),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    Odrv12 I__7334 (
            .O(N__32144),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    InMux I__7333 (
            .O(N__32137),
            .I(N__32134));
    LocalMux I__7332 (
            .O(N__32134),
            .I(N__32131));
    Span4Mux_v I__7331 (
            .O(N__32131),
            .I(N__32128));
    Odrv4 I__7330 (
            .O(N__32128),
            .I(\VPP_VDDQ.un9_clk_100khz_1 ));
    InMux I__7329 (
            .O(N__32125),
            .I(N__32122));
    LocalMux I__7328 (
            .O(N__32122),
            .I(\VPP_VDDQ.count_2_RNIZ0Z_1 ));
    InMux I__7327 (
            .O(N__32119),
            .I(N__32113));
    InMux I__7326 (
            .O(N__32118),
            .I(N__32113));
    LocalMux I__7325 (
            .O(N__32113),
            .I(\VPP_VDDQ.count_2Z0Z_1 ));
    InMux I__7324 (
            .O(N__32110),
            .I(N__32104));
    InMux I__7323 (
            .O(N__32109),
            .I(N__32104));
    LocalMux I__7322 (
            .O(N__32104),
            .I(N__32101));
    Odrv4 I__7321 (
            .O(N__32101),
            .I(\VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ));
    InMux I__7320 (
            .O(N__32098),
            .I(N__32095));
    LocalMux I__7319 (
            .O(N__32095),
            .I(\VPP_VDDQ.count_2_0_11 ));
    CascadeMux I__7318 (
            .O(N__32092),
            .I(\VPP_VDDQ.count_2_1_11_cascade_ ));
    CEMux I__7317 (
            .O(N__32089),
            .I(N__32086));
    LocalMux I__7316 (
            .O(N__32086),
            .I(N__32083));
    Span4Mux_v I__7315 (
            .O(N__32083),
            .I(N__32070));
    InMux I__7314 (
            .O(N__32082),
            .I(N__32065));
    InMux I__7313 (
            .O(N__32081),
            .I(N__32065));
    InMux I__7312 (
            .O(N__32080),
            .I(N__32060));
    InMux I__7311 (
            .O(N__32079),
            .I(N__32060));
    InMux I__7310 (
            .O(N__32078),
            .I(N__32054));
    CEMux I__7309 (
            .O(N__32077),
            .I(N__32054));
    CascadeMux I__7308 (
            .O(N__32076),
            .I(N__32051));
    InMux I__7307 (
            .O(N__32075),
            .I(N__32045));
    CEMux I__7306 (
            .O(N__32074),
            .I(N__32045));
    CEMux I__7305 (
            .O(N__32073),
            .I(N__32042));
    Span4Mux_s0_v I__7304 (
            .O(N__32070),
            .I(N__32035));
    LocalMux I__7303 (
            .O(N__32065),
            .I(N__32035));
    LocalMux I__7302 (
            .O(N__32060),
            .I(N__32035));
    CEMux I__7301 (
            .O(N__32059),
            .I(N__32029));
    LocalMux I__7300 (
            .O(N__32054),
            .I(N__32026));
    InMux I__7299 (
            .O(N__32051),
            .I(N__32021));
    InMux I__7298 (
            .O(N__32050),
            .I(N__32021));
    LocalMux I__7297 (
            .O(N__32045),
            .I(N__32017));
    LocalMux I__7296 (
            .O(N__32042),
            .I(N__32011));
    Span4Mux_v I__7295 (
            .O(N__32035),
            .I(N__32011));
    InMux I__7294 (
            .O(N__32034),
            .I(N__32001));
    InMux I__7293 (
            .O(N__32033),
            .I(N__32001));
    CEMux I__7292 (
            .O(N__32032),
            .I(N__32001));
    LocalMux I__7291 (
            .O(N__32029),
            .I(N__31998));
    Span4Mux_v I__7290 (
            .O(N__32026),
            .I(N__31995));
    LocalMux I__7289 (
            .O(N__32021),
            .I(N__31992));
    InMux I__7288 (
            .O(N__32020),
            .I(N__31989));
    Span4Mux_v I__7287 (
            .O(N__32017),
            .I(N__31982));
    InMux I__7286 (
            .O(N__32016),
            .I(N__31979));
    Sp12to4 I__7285 (
            .O(N__32011),
            .I(N__31976));
    InMux I__7284 (
            .O(N__32010),
            .I(N__31971));
    InMux I__7283 (
            .O(N__32009),
            .I(N__31971));
    InMux I__7282 (
            .O(N__32008),
            .I(N__31968));
    LocalMux I__7281 (
            .O(N__32001),
            .I(N__31965));
    Span4Mux_h I__7280 (
            .O(N__31998),
            .I(N__31956));
    Span4Mux_s0_h I__7279 (
            .O(N__31995),
            .I(N__31956));
    Span4Mux_h I__7278 (
            .O(N__31992),
            .I(N__31956));
    LocalMux I__7277 (
            .O(N__31989),
            .I(N__31956));
    InMux I__7276 (
            .O(N__31988),
            .I(N__31951));
    InMux I__7275 (
            .O(N__31987),
            .I(N__31951));
    InMux I__7274 (
            .O(N__31986),
            .I(N__31948));
    InMux I__7273 (
            .O(N__31985),
            .I(N__31945));
    Sp12to4 I__7272 (
            .O(N__31982),
            .I(N__31934));
    LocalMux I__7271 (
            .O(N__31979),
            .I(N__31934));
    Span12Mux_s4_h I__7270 (
            .O(N__31976),
            .I(N__31934));
    LocalMux I__7269 (
            .O(N__31971),
            .I(N__31934));
    LocalMux I__7268 (
            .O(N__31968),
            .I(N__31934));
    Sp12to4 I__7267 (
            .O(N__31965),
            .I(N__31925));
    Sp12to4 I__7266 (
            .O(N__31956),
            .I(N__31925));
    LocalMux I__7265 (
            .O(N__31951),
            .I(N__31925));
    LocalMux I__7264 (
            .O(N__31948),
            .I(N__31925));
    LocalMux I__7263 (
            .O(N__31945),
            .I(N__31920));
    Span12Mux_v I__7262 (
            .O(N__31934),
            .I(N__31920));
    Span12Mux_s4_v I__7261 (
            .O(N__31925),
            .I(N__31917));
    Odrv12 I__7260 (
            .O(N__31920),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    Odrv12 I__7259 (
            .O(N__31917),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    InMux I__7258 (
            .O(N__31912),
            .I(N__31909));
    LocalMux I__7257 (
            .O(N__31909),
            .I(N__31905));
    InMux I__7256 (
            .O(N__31908),
            .I(N__31902));
    Odrv4 I__7255 (
            .O(N__31905),
            .I(\VPP_VDDQ.count_2Z0Z_11 ));
    LocalMux I__7254 (
            .O(N__31902),
            .I(\VPP_VDDQ.count_2Z0Z_11 ));
    InMux I__7253 (
            .O(N__31897),
            .I(N__31888));
    InMux I__7252 (
            .O(N__31896),
            .I(N__31885));
    CascadeMux I__7251 (
            .O(N__31895),
            .I(N__31880));
    InMux I__7250 (
            .O(N__31894),
            .I(N__31876));
    CascadeMux I__7249 (
            .O(N__31893),
            .I(N__31872));
    InMux I__7248 (
            .O(N__31892),
            .I(N__31869));
    InMux I__7247 (
            .O(N__31891),
            .I(N__31866));
    LocalMux I__7246 (
            .O(N__31888),
            .I(N__31861));
    LocalMux I__7245 (
            .O(N__31885),
            .I(N__31861));
    InMux I__7244 (
            .O(N__31884),
            .I(N__31857));
    InMux I__7243 (
            .O(N__31883),
            .I(N__31852));
    InMux I__7242 (
            .O(N__31880),
            .I(N__31852));
    InMux I__7241 (
            .O(N__31879),
            .I(N__31848));
    LocalMux I__7240 (
            .O(N__31876),
            .I(N__31845));
    InMux I__7239 (
            .O(N__31875),
            .I(N__31840));
    InMux I__7238 (
            .O(N__31872),
            .I(N__31840));
    LocalMux I__7237 (
            .O(N__31869),
            .I(N__31833));
    LocalMux I__7236 (
            .O(N__31866),
            .I(N__31833));
    Span4Mux_v I__7235 (
            .O(N__31861),
            .I(N__31833));
    InMux I__7234 (
            .O(N__31860),
            .I(N__31830));
    LocalMux I__7233 (
            .O(N__31857),
            .I(N__31827));
    LocalMux I__7232 (
            .O(N__31852),
            .I(N__31824));
    InMux I__7231 (
            .O(N__31851),
            .I(N__31821));
    LocalMux I__7230 (
            .O(N__31848),
            .I(N__31818));
    Span4Mux_v I__7229 (
            .O(N__31845),
            .I(N__31809));
    LocalMux I__7228 (
            .O(N__31840),
            .I(N__31809));
    Span4Mux_h I__7227 (
            .O(N__31833),
            .I(N__31809));
    LocalMux I__7226 (
            .O(N__31830),
            .I(N__31809));
    Span4Mux_h I__7225 (
            .O(N__31827),
            .I(N__31806));
    Odrv12 I__7224 (
            .O(N__31824),
            .I(func_state_RNI_3_0));
    LocalMux I__7223 (
            .O(N__31821),
            .I(func_state_RNI_3_0));
    Odrv12 I__7222 (
            .O(N__31818),
            .I(func_state_RNI_3_0));
    Odrv4 I__7221 (
            .O(N__31809),
            .I(func_state_RNI_3_0));
    Odrv4 I__7220 (
            .O(N__31806),
            .I(func_state_RNI_3_0));
    CascadeMux I__7219 (
            .O(N__31795),
            .I(N__31792));
    InMux I__7218 (
            .O(N__31792),
            .I(N__31783));
    InMux I__7217 (
            .O(N__31791),
            .I(N__31780));
    InMux I__7216 (
            .O(N__31790),
            .I(N__31777));
    InMux I__7215 (
            .O(N__31789),
            .I(N__31768));
    InMux I__7214 (
            .O(N__31788),
            .I(N__31768));
    InMux I__7213 (
            .O(N__31787),
            .I(N__31768));
    InMux I__7212 (
            .O(N__31786),
            .I(N__31765));
    LocalMux I__7211 (
            .O(N__31783),
            .I(N__31757));
    LocalMux I__7210 (
            .O(N__31780),
            .I(N__31757));
    LocalMux I__7209 (
            .O(N__31777),
            .I(N__31757));
    InMux I__7208 (
            .O(N__31776),
            .I(N__31754));
    CascadeMux I__7207 (
            .O(N__31775),
            .I(N__31750));
    LocalMux I__7206 (
            .O(N__31768),
            .I(N__31745));
    LocalMux I__7205 (
            .O(N__31765),
            .I(N__31742));
    InMux I__7204 (
            .O(N__31764),
            .I(N__31739));
    Span4Mux_v I__7203 (
            .O(N__31757),
            .I(N__31736));
    LocalMux I__7202 (
            .O(N__31754),
            .I(N__31733));
    InMux I__7201 (
            .O(N__31753),
            .I(N__31730));
    InMux I__7200 (
            .O(N__31750),
            .I(N__31727));
    InMux I__7199 (
            .O(N__31749),
            .I(N__31724));
    InMux I__7198 (
            .O(N__31748),
            .I(N__31721));
    Span4Mux_v I__7197 (
            .O(N__31745),
            .I(N__31717));
    Span4Mux_v I__7196 (
            .O(N__31742),
            .I(N__31712));
    LocalMux I__7195 (
            .O(N__31739),
            .I(N__31712));
    Span4Mux_h I__7194 (
            .O(N__31736),
            .I(N__31703));
    Span4Mux_v I__7193 (
            .O(N__31733),
            .I(N__31703));
    LocalMux I__7192 (
            .O(N__31730),
            .I(N__31703));
    LocalMux I__7191 (
            .O(N__31727),
            .I(N__31703));
    LocalMux I__7190 (
            .O(N__31724),
            .I(N__31698));
    LocalMux I__7189 (
            .O(N__31721),
            .I(N__31698));
    InMux I__7188 (
            .O(N__31720),
            .I(N__31695));
    Span4Mux_h I__7187 (
            .O(N__31717),
            .I(N__31692));
    Span4Mux_v I__7186 (
            .O(N__31712),
            .I(N__31687));
    Span4Mux_v I__7185 (
            .O(N__31703),
            .I(N__31687));
    Span4Mux_v I__7184 (
            .O(N__31698),
            .I(N__31682));
    LocalMux I__7183 (
            .O(N__31695),
            .I(N__31682));
    Span4Mux_v I__7182 (
            .O(N__31692),
            .I(N__31679));
    Span4Mux_h I__7181 (
            .O(N__31687),
            .I(N__31674));
    Span4Mux_v I__7180 (
            .O(N__31682),
            .I(N__31674));
    Odrv4 I__7179 (
            .O(N__31679),
            .I(gpio_fpga_soc_4));
    Odrv4 I__7178 (
            .O(N__31674),
            .I(gpio_fpga_soc_4));
    InMux I__7177 (
            .O(N__31669),
            .I(N__31666));
    LocalMux I__7176 (
            .O(N__31666),
            .I(N__31663));
    Odrv12 I__7175 (
            .O(N__31663),
            .I(\POWERLED.dutycycle_1_0_iv_i_a2_sx_5 ));
    InMux I__7174 (
            .O(N__31660),
            .I(N__31656));
    InMux I__7173 (
            .O(N__31659),
            .I(N__31653));
    LocalMux I__7172 (
            .O(N__31656),
            .I(N__31648));
    LocalMux I__7171 (
            .O(N__31653),
            .I(N__31648));
    Span12Mux_s7_v I__7170 (
            .O(N__31648),
            .I(N__31645));
    Odrv12 I__7169 (
            .O(N__31645),
            .I(\VPP_VDDQ.N_2112_i ));
    InMux I__7168 (
            .O(N__31642),
            .I(N__31639));
    LocalMux I__7167 (
            .O(N__31639),
            .I(N__31635));
    CascadeMux I__7166 (
            .O(N__31638),
            .I(N__31632));
    Span4Mux_v I__7165 (
            .O(N__31635),
            .I(N__31629));
    InMux I__7164 (
            .O(N__31632),
            .I(N__31626));
    Odrv4 I__7163 (
            .O(N__31629),
            .I(\VPP_VDDQ.count_2Z0Z_9 ));
    LocalMux I__7162 (
            .O(N__31626),
            .I(\VPP_VDDQ.count_2Z0Z_9 ));
    CascadeMux I__7161 (
            .O(N__31621),
            .I(\VPP_VDDQ.count_2_1_7_cascade_ ));
    InMux I__7160 (
            .O(N__31618),
            .I(N__31615));
    LocalMux I__7159 (
            .O(N__31615),
            .I(N__31612));
    Span4Mux_v I__7158 (
            .O(N__31612),
            .I(N__31609));
    Odrv4 I__7157 (
            .O(N__31609),
            .I(\VPP_VDDQ.un9_clk_100khz_10 ));
    InMux I__7156 (
            .O(N__31606),
            .I(N__31603));
    LocalMux I__7155 (
            .O(N__31603),
            .I(N__31600));
    Span4Mux_v I__7154 (
            .O(N__31600),
            .I(N__31596));
    InMux I__7153 (
            .O(N__31599),
            .I(N__31593));
    Odrv4 I__7152 (
            .O(N__31596),
            .I(\VPP_VDDQ.count_2Z0Z_10 ));
    LocalMux I__7151 (
            .O(N__31593),
            .I(\VPP_VDDQ.count_2Z0Z_10 ));
    CascadeMux I__7150 (
            .O(N__31588),
            .I(\VPP_VDDQ.un9_clk_100khz_7_cascade_ ));
    InMux I__7149 (
            .O(N__31585),
            .I(N__31582));
    LocalMux I__7148 (
            .O(N__31582),
            .I(N__31579));
    Span4Mux_h I__7147 (
            .O(N__31579),
            .I(N__31576));
    Odrv4 I__7146 (
            .O(N__31576),
            .I(\VPP_VDDQ.un9_clk_100khz_13 ));
    CascadeMux I__7145 (
            .O(N__31573),
            .I(\VPP_VDDQ.count_2_1_0_cascade_ ));
    CascadeMux I__7144 (
            .O(N__31570),
            .I(\VPP_VDDQ.count_2Z0Z_0_cascade_ ));
    InMux I__7143 (
            .O(N__31567),
            .I(N__31564));
    LocalMux I__7142 (
            .O(N__31564),
            .I(\VPP_VDDQ.count_2_0_0 ));
    InMux I__7141 (
            .O(N__31561),
            .I(N__31555));
    InMux I__7140 (
            .O(N__31560),
            .I(N__31555));
    LocalMux I__7139 (
            .O(N__31555),
            .I(N__31552));
    Odrv12 I__7138 (
            .O(N__31552),
            .I(\VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7 ));
    InMux I__7137 (
            .O(N__31549),
            .I(N__31544));
    InMux I__7136 (
            .O(N__31548),
            .I(N__31541));
    InMux I__7135 (
            .O(N__31547),
            .I(N__31538));
    LocalMux I__7134 (
            .O(N__31544),
            .I(N__31534));
    LocalMux I__7133 (
            .O(N__31541),
            .I(N__31528));
    LocalMux I__7132 (
            .O(N__31538),
            .I(N__31528));
    InMux I__7131 (
            .O(N__31537),
            .I(N__31525));
    Span4Mux_v I__7130 (
            .O(N__31534),
            .I(N__31517));
    InMux I__7129 (
            .O(N__31533),
            .I(N__31514));
    Span4Mux_h I__7128 (
            .O(N__31528),
            .I(N__31509));
    LocalMux I__7127 (
            .O(N__31525),
            .I(N__31509));
    InMux I__7126 (
            .O(N__31524),
            .I(N__31506));
    InMux I__7125 (
            .O(N__31523),
            .I(N__31501));
    InMux I__7124 (
            .O(N__31522),
            .I(N__31501));
    InMux I__7123 (
            .O(N__31521),
            .I(N__31498));
    InMux I__7122 (
            .O(N__31520),
            .I(N__31495));
    Odrv4 I__7121 (
            .O(N__31517),
            .I(\POWERLED.dutycycle ));
    LocalMux I__7120 (
            .O(N__31514),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__7119 (
            .O(N__31509),
            .I(\POWERLED.dutycycle ));
    LocalMux I__7118 (
            .O(N__31506),
            .I(\POWERLED.dutycycle ));
    LocalMux I__7117 (
            .O(N__31501),
            .I(\POWERLED.dutycycle ));
    LocalMux I__7116 (
            .O(N__31498),
            .I(\POWERLED.dutycycle ));
    LocalMux I__7115 (
            .O(N__31495),
            .I(\POWERLED.dutycycle ));
    CascadeMux I__7114 (
            .O(N__31480),
            .I(N__31475));
    InMux I__7113 (
            .O(N__31479),
            .I(N__31472));
    InMux I__7112 (
            .O(N__31478),
            .I(N__31465));
    InMux I__7111 (
            .O(N__31475),
            .I(N__31465));
    LocalMux I__7110 (
            .O(N__31472),
            .I(N__31461));
    CascadeMux I__7109 (
            .O(N__31471),
            .I(N__31456));
    InMux I__7108 (
            .O(N__31470),
            .I(N__31452));
    LocalMux I__7107 (
            .O(N__31465),
            .I(N__31449));
    CascadeMux I__7106 (
            .O(N__31464),
            .I(N__31446));
    Span4Mux_v I__7105 (
            .O(N__31461),
            .I(N__31443));
    InMux I__7104 (
            .O(N__31460),
            .I(N__31440));
    InMux I__7103 (
            .O(N__31459),
            .I(N__31437));
    InMux I__7102 (
            .O(N__31456),
            .I(N__31434));
    InMux I__7101 (
            .O(N__31455),
            .I(N__31431));
    LocalMux I__7100 (
            .O(N__31452),
            .I(N__31428));
    Sp12to4 I__7099 (
            .O(N__31449),
            .I(N__31425));
    InMux I__7098 (
            .O(N__31446),
            .I(N__31422));
    Odrv4 I__7097 (
            .O(N__31443),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__7096 (
            .O(N__31440),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__7095 (
            .O(N__31437),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__7094 (
            .O(N__31434),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__7093 (
            .O(N__31431),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__7092 (
            .O(N__31428),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv12 I__7091 (
            .O(N__31425),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__7090 (
            .O(N__31422),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    InMux I__7089 (
            .O(N__31405),
            .I(N__31401));
    InMux I__7088 (
            .O(N__31404),
            .I(N__31398));
    LocalMux I__7087 (
            .O(N__31401),
            .I(\POWERLED.N_493 ));
    LocalMux I__7086 (
            .O(N__31398),
            .I(\POWERLED.N_493 ));
    InMux I__7085 (
            .O(N__31393),
            .I(N__31390));
    LocalMux I__7084 (
            .O(N__31390),
            .I(\POWERLED.g1_0_7 ));
    InMux I__7083 (
            .O(N__31387),
            .I(N__31384));
    LocalMux I__7082 (
            .O(N__31384),
            .I(\POWERLED.g1_0_2 ));
    CascadeMux I__7081 (
            .O(N__31381),
            .I(\POWERLED.g1_0_8_cascade_ ));
    CascadeMux I__7080 (
            .O(N__31378),
            .I(N__31370));
    CascadeMux I__7079 (
            .O(N__31377),
            .I(N__31366));
    CascadeMux I__7078 (
            .O(N__31376),
            .I(N__31361));
    CascadeMux I__7077 (
            .O(N__31375),
            .I(N__31355));
    CascadeMux I__7076 (
            .O(N__31374),
            .I(N__31352));
    InMux I__7075 (
            .O(N__31373),
            .I(N__31338));
    InMux I__7074 (
            .O(N__31370),
            .I(N__31335));
    InMux I__7073 (
            .O(N__31369),
            .I(N__31332));
    InMux I__7072 (
            .O(N__31366),
            .I(N__31327));
    InMux I__7071 (
            .O(N__31365),
            .I(N__31327));
    CascadeMux I__7070 (
            .O(N__31364),
            .I(N__31324));
    InMux I__7069 (
            .O(N__31361),
            .I(N__31311));
    InMux I__7068 (
            .O(N__31360),
            .I(N__31311));
    InMux I__7067 (
            .O(N__31359),
            .I(N__31311));
    InMux I__7066 (
            .O(N__31358),
            .I(N__31311));
    InMux I__7065 (
            .O(N__31355),
            .I(N__31302));
    InMux I__7064 (
            .O(N__31352),
            .I(N__31302));
    InMux I__7063 (
            .O(N__31351),
            .I(N__31302));
    InMux I__7062 (
            .O(N__31350),
            .I(N__31302));
    InMux I__7061 (
            .O(N__31349),
            .I(N__31299));
    InMux I__7060 (
            .O(N__31348),
            .I(N__31296));
    InMux I__7059 (
            .O(N__31347),
            .I(N__31291));
    InMux I__7058 (
            .O(N__31346),
            .I(N__31291));
    CascadeMux I__7057 (
            .O(N__31345),
            .I(N__31284));
    InMux I__7056 (
            .O(N__31344),
            .I(N__31278));
    InMux I__7055 (
            .O(N__31343),
            .I(N__31278));
    InMux I__7054 (
            .O(N__31342),
            .I(N__31273));
    InMux I__7053 (
            .O(N__31341),
            .I(N__31273));
    LocalMux I__7052 (
            .O(N__31338),
            .I(N__31264));
    LocalMux I__7051 (
            .O(N__31335),
            .I(N__31264));
    LocalMux I__7050 (
            .O(N__31332),
            .I(N__31264));
    LocalMux I__7049 (
            .O(N__31327),
            .I(N__31264));
    InMux I__7048 (
            .O(N__31324),
            .I(N__31261));
    InMux I__7047 (
            .O(N__31323),
            .I(N__31256));
    InMux I__7046 (
            .O(N__31322),
            .I(N__31256));
    InMux I__7045 (
            .O(N__31321),
            .I(N__31251));
    InMux I__7044 (
            .O(N__31320),
            .I(N__31251));
    LocalMux I__7043 (
            .O(N__31311),
            .I(N__31246));
    LocalMux I__7042 (
            .O(N__31302),
            .I(N__31246));
    LocalMux I__7041 (
            .O(N__31299),
            .I(N__31239));
    LocalMux I__7040 (
            .O(N__31296),
            .I(N__31239));
    LocalMux I__7039 (
            .O(N__31291),
            .I(N__31239));
    InMux I__7038 (
            .O(N__31290),
            .I(N__31234));
    InMux I__7037 (
            .O(N__31289),
            .I(N__31234));
    InMux I__7036 (
            .O(N__31288),
            .I(N__31231));
    InMux I__7035 (
            .O(N__31287),
            .I(N__31224));
    InMux I__7034 (
            .O(N__31284),
            .I(N__31224));
    InMux I__7033 (
            .O(N__31283),
            .I(N__31224));
    LocalMux I__7032 (
            .O(N__31278),
            .I(N__31221));
    LocalMux I__7031 (
            .O(N__31273),
            .I(N__31214));
    Span4Mux_v I__7030 (
            .O(N__31264),
            .I(N__31214));
    LocalMux I__7029 (
            .O(N__31261),
            .I(N__31214));
    LocalMux I__7028 (
            .O(N__31256),
            .I(N__31207));
    LocalMux I__7027 (
            .O(N__31251),
            .I(N__31207));
    Span4Mux_s3_h I__7026 (
            .O(N__31246),
            .I(N__31207));
    Span12Mux_s4_h I__7025 (
            .O(N__31239),
            .I(N__31204));
    LocalMux I__7024 (
            .O(N__31234),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    LocalMux I__7023 (
            .O(N__31231),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    LocalMux I__7022 (
            .O(N__31224),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv12 I__7021 (
            .O(N__31221),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv4 I__7020 (
            .O(N__31214),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv4 I__7019 (
            .O(N__31207),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv12 I__7018 (
            .O(N__31204),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    InMux I__7017 (
            .O(N__31189),
            .I(N__31186));
    LocalMux I__7016 (
            .O(N__31186),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_6 ));
    InMux I__7015 (
            .O(N__31183),
            .I(N__31176));
    InMux I__7014 (
            .O(N__31182),
            .I(N__31173));
    InMux I__7013 (
            .O(N__31181),
            .I(N__31168));
    InMux I__7012 (
            .O(N__31180),
            .I(N__31168));
    InMux I__7011 (
            .O(N__31179),
            .I(N__31165));
    LocalMux I__7010 (
            .O(N__31176),
            .I(N__31161));
    LocalMux I__7009 (
            .O(N__31173),
            .I(N__31158));
    LocalMux I__7008 (
            .O(N__31168),
            .I(N__31155));
    LocalMux I__7007 (
            .O(N__31165),
            .I(N__31152));
    CascadeMux I__7006 (
            .O(N__31164),
            .I(N__31149));
    Span4Mux_h I__7005 (
            .O(N__31161),
            .I(N__31145));
    Span4Mux_s3_h I__7004 (
            .O(N__31158),
            .I(N__31140));
    Span4Mux_h I__7003 (
            .O(N__31155),
            .I(N__31140));
    Span4Mux_h I__7002 (
            .O(N__31152),
            .I(N__31137));
    InMux I__7001 (
            .O(N__31149),
            .I(N__31134));
    InMux I__7000 (
            .O(N__31148),
            .I(N__31131));
    Odrv4 I__6999 (
            .O(N__31145),
            .I(RSMRSTn_fast));
    Odrv4 I__6998 (
            .O(N__31140),
            .I(RSMRSTn_fast));
    Odrv4 I__6997 (
            .O(N__31137),
            .I(RSMRSTn_fast));
    LocalMux I__6996 (
            .O(N__31134),
            .I(RSMRSTn_fast));
    LocalMux I__6995 (
            .O(N__31131),
            .I(RSMRSTn_fast));
    CascadeMux I__6994 (
            .O(N__31120),
            .I(\RSMRST_PWRGD.N_8_0_0_cascade_ ));
    CascadeMux I__6993 (
            .O(N__31117),
            .I(N__31111));
    CascadeMux I__6992 (
            .O(N__31116),
            .I(N__31105));
    CascadeMux I__6991 (
            .O(N__31115),
            .I(N__31099));
    InMux I__6990 (
            .O(N__31114),
            .I(N__31089));
    InMux I__6989 (
            .O(N__31111),
            .I(N__31089));
    InMux I__6988 (
            .O(N__31110),
            .I(N__31083));
    CascadeMux I__6987 (
            .O(N__31109),
            .I(N__31076));
    InMux I__6986 (
            .O(N__31108),
            .I(N__31073));
    InMux I__6985 (
            .O(N__31105),
            .I(N__31069));
    CascadeMux I__6984 (
            .O(N__31104),
            .I(N__31066));
    CascadeMux I__6983 (
            .O(N__31103),
            .I(N__31062));
    InMux I__6982 (
            .O(N__31102),
            .I(N__31056));
    InMux I__6981 (
            .O(N__31099),
            .I(N__31056));
    InMux I__6980 (
            .O(N__31098),
            .I(N__31053));
    InMux I__6979 (
            .O(N__31097),
            .I(N__31040));
    InMux I__6978 (
            .O(N__31096),
            .I(N__31040));
    InMux I__6977 (
            .O(N__31095),
            .I(N__31040));
    InMux I__6976 (
            .O(N__31094),
            .I(N__31040));
    LocalMux I__6975 (
            .O(N__31089),
            .I(N__31037));
    InMux I__6974 (
            .O(N__31088),
            .I(N__31030));
    InMux I__6973 (
            .O(N__31087),
            .I(N__31030));
    InMux I__6972 (
            .O(N__31086),
            .I(N__31030));
    LocalMux I__6971 (
            .O(N__31083),
            .I(N__31027));
    InMux I__6970 (
            .O(N__31082),
            .I(N__31024));
    InMux I__6969 (
            .O(N__31081),
            .I(N__31021));
    InMux I__6968 (
            .O(N__31080),
            .I(N__31018));
    InMux I__6967 (
            .O(N__31079),
            .I(N__31012));
    InMux I__6966 (
            .O(N__31076),
            .I(N__31012));
    LocalMux I__6965 (
            .O(N__31073),
            .I(N__31009));
    InMux I__6964 (
            .O(N__31072),
            .I(N__31006));
    LocalMux I__6963 (
            .O(N__31069),
            .I(N__31003));
    InMux I__6962 (
            .O(N__31066),
            .I(N__30996));
    InMux I__6961 (
            .O(N__31065),
            .I(N__30996));
    InMux I__6960 (
            .O(N__31062),
            .I(N__30993));
    InMux I__6959 (
            .O(N__31061),
            .I(N__30990));
    LocalMux I__6958 (
            .O(N__31056),
            .I(N__30987));
    LocalMux I__6957 (
            .O(N__31053),
            .I(N__30984));
    InMux I__6956 (
            .O(N__31052),
            .I(N__30974));
    InMux I__6955 (
            .O(N__31051),
            .I(N__30974));
    InMux I__6954 (
            .O(N__31050),
            .I(N__30974));
    InMux I__6953 (
            .O(N__31049),
            .I(N__30974));
    LocalMux I__6952 (
            .O(N__31040),
            .I(N__30967));
    Span4Mux_s1_h I__6951 (
            .O(N__31037),
            .I(N__30967));
    LocalMux I__6950 (
            .O(N__31030),
            .I(N__30967));
    Span4Mux_s1_h I__6949 (
            .O(N__31027),
            .I(N__30962));
    LocalMux I__6948 (
            .O(N__31024),
            .I(N__30962));
    LocalMux I__6947 (
            .O(N__31021),
            .I(N__30959));
    LocalMux I__6946 (
            .O(N__31018),
            .I(N__30956));
    InMux I__6945 (
            .O(N__31017),
            .I(N__30953));
    LocalMux I__6944 (
            .O(N__31012),
            .I(N__30948));
    Span4Mux_s1_h I__6943 (
            .O(N__31009),
            .I(N__30948));
    LocalMux I__6942 (
            .O(N__31006),
            .I(N__30945));
    Span4Mux_s1_h I__6941 (
            .O(N__31003),
            .I(N__30942));
    InMux I__6940 (
            .O(N__31002),
            .I(N__30937));
    InMux I__6939 (
            .O(N__31001),
            .I(N__30937));
    LocalMux I__6938 (
            .O(N__30996),
            .I(N__30932));
    LocalMux I__6937 (
            .O(N__30993),
            .I(N__30932));
    LocalMux I__6936 (
            .O(N__30990),
            .I(N__30929));
    Span4Mux_h I__6935 (
            .O(N__30987),
            .I(N__30926));
    Span12Mux_s8_v I__6934 (
            .O(N__30984),
            .I(N__30923));
    InMux I__6933 (
            .O(N__30983),
            .I(N__30920));
    LocalMux I__6932 (
            .O(N__30974),
            .I(N__30915));
    Span4Mux_h I__6931 (
            .O(N__30967),
            .I(N__30915));
    Span4Mux_h I__6930 (
            .O(N__30962),
            .I(N__30904));
    Span4Mux_v I__6929 (
            .O(N__30959),
            .I(N__30904));
    Span4Mux_h I__6928 (
            .O(N__30956),
            .I(N__30904));
    LocalMux I__6927 (
            .O(N__30953),
            .I(N__30904));
    Span4Mux_h I__6926 (
            .O(N__30948),
            .I(N__30904));
    Span4Mux_s1_h I__6925 (
            .O(N__30945),
            .I(N__30895));
    Span4Mux_v I__6924 (
            .O(N__30942),
            .I(N__30895));
    LocalMux I__6923 (
            .O(N__30937),
            .I(N__30895));
    Span4Mux_v I__6922 (
            .O(N__30932),
            .I(N__30895));
    Odrv4 I__6921 (
            .O(N__30929),
            .I(func_state_RNIOGRS_1));
    Odrv4 I__6920 (
            .O(N__30926),
            .I(func_state_RNIOGRS_1));
    Odrv12 I__6919 (
            .O(N__30923),
            .I(func_state_RNIOGRS_1));
    LocalMux I__6918 (
            .O(N__30920),
            .I(func_state_RNIOGRS_1));
    Odrv4 I__6917 (
            .O(N__30915),
            .I(func_state_RNIOGRS_1));
    Odrv4 I__6916 (
            .O(N__30904),
            .I(func_state_RNIOGRS_1));
    Odrv4 I__6915 (
            .O(N__30895),
            .I(func_state_RNIOGRS_1));
    InMux I__6914 (
            .O(N__30880),
            .I(N__30875));
    CascadeMux I__6913 (
            .O(N__30879),
            .I(N__30872));
    CascadeMux I__6912 (
            .O(N__30878),
            .I(N__30866));
    LocalMux I__6911 (
            .O(N__30875),
            .I(N__30862));
    InMux I__6910 (
            .O(N__30872),
            .I(N__30856));
    InMux I__6909 (
            .O(N__30871),
            .I(N__30856));
    InMux I__6908 (
            .O(N__30870),
            .I(N__30853));
    CascadeMux I__6907 (
            .O(N__30869),
            .I(N__30849));
    InMux I__6906 (
            .O(N__30866),
            .I(N__30844));
    InMux I__6905 (
            .O(N__30865),
            .I(N__30844));
    Span4Mux_v I__6904 (
            .O(N__30862),
            .I(N__30841));
    InMux I__6903 (
            .O(N__30861),
            .I(N__30838));
    LocalMux I__6902 (
            .O(N__30856),
            .I(N__30833));
    LocalMux I__6901 (
            .O(N__30853),
            .I(N__30833));
    InMux I__6900 (
            .O(N__30852),
            .I(N__30830));
    InMux I__6899 (
            .O(N__30849),
            .I(N__30826));
    LocalMux I__6898 (
            .O(N__30844),
            .I(N__30823));
    Span4Mux_v I__6897 (
            .O(N__30841),
            .I(N__30818));
    LocalMux I__6896 (
            .O(N__30838),
            .I(N__30818));
    Span4Mux_v I__6895 (
            .O(N__30833),
            .I(N__30813));
    LocalMux I__6894 (
            .O(N__30830),
            .I(N__30813));
    InMux I__6893 (
            .O(N__30829),
            .I(N__30810));
    LocalMux I__6892 (
            .O(N__30826),
            .I(N__30807));
    Odrv12 I__6891 (
            .O(N__30823),
            .I(dutycycle_RNIKBMSJ_0_5));
    Odrv4 I__6890 (
            .O(N__30818),
            .I(dutycycle_RNIKBMSJ_0_5));
    Odrv4 I__6889 (
            .O(N__30813),
            .I(dutycycle_RNIKBMSJ_0_5));
    LocalMux I__6888 (
            .O(N__30810),
            .I(dutycycle_RNIKBMSJ_0_5));
    Odrv4 I__6887 (
            .O(N__30807),
            .I(dutycycle_RNIKBMSJ_0_5));
    InMux I__6886 (
            .O(N__30796),
            .I(N__30793));
    LocalMux I__6885 (
            .O(N__30793),
            .I(POWERLED_g1));
    CascadeMux I__6884 (
            .O(N__30790),
            .I(\RSMRST_PWRGD.N_9_0_cascade_ ));
    InMux I__6883 (
            .O(N__30787),
            .I(N__30784));
    LocalMux I__6882 (
            .O(N__30784),
            .I(N_46));
    InMux I__6881 (
            .O(N__30781),
            .I(N__30778));
    LocalMux I__6880 (
            .O(N__30778),
            .I(N__30775));
    Odrv12 I__6879 (
            .O(N__30775),
            .I(\RSMRST_PWRGD.N_11 ));
    InMux I__6878 (
            .O(N__30772),
            .I(N__30765));
    InMux I__6877 (
            .O(N__30771),
            .I(N__30761));
    InMux I__6876 (
            .O(N__30770),
            .I(N__30758));
    InMux I__6875 (
            .O(N__30769),
            .I(N__30755));
    InMux I__6874 (
            .O(N__30768),
            .I(N__30752));
    LocalMux I__6873 (
            .O(N__30765),
            .I(N__30749));
    InMux I__6872 (
            .O(N__30764),
            .I(N__30745));
    LocalMux I__6871 (
            .O(N__30761),
            .I(N__30742));
    LocalMux I__6870 (
            .O(N__30758),
            .I(N__30739));
    LocalMux I__6869 (
            .O(N__30755),
            .I(N__30734));
    LocalMux I__6868 (
            .O(N__30752),
            .I(N__30734));
    Span4Mux_s2_h I__6867 (
            .O(N__30749),
            .I(N__30731));
    InMux I__6866 (
            .O(N__30748),
            .I(N__30728));
    LocalMux I__6865 (
            .O(N__30745),
            .I(N__30725));
    Span4Mux_s1_h I__6864 (
            .O(N__30742),
            .I(N__30720));
    Span4Mux_s1_h I__6863 (
            .O(N__30739),
            .I(N__30720));
    Span4Mux_v I__6862 (
            .O(N__30734),
            .I(N__30717));
    Span4Mux_h I__6861 (
            .O(N__30731),
            .I(N__30712));
    LocalMux I__6860 (
            .O(N__30728),
            .I(N__30712));
    Span4Mux_v I__6859 (
            .O(N__30725),
            .I(N__30707));
    Span4Mux_h I__6858 (
            .O(N__30720),
            .I(N__30707));
    Odrv4 I__6857 (
            .O(N__30717),
            .I(\POWERLED.N_341 ));
    Odrv4 I__6856 (
            .O(N__30712),
            .I(\POWERLED.N_341 ));
    Odrv4 I__6855 (
            .O(N__30707),
            .I(\POWERLED.N_341 ));
    InMux I__6854 (
            .O(N__30700),
            .I(N__30695));
    InMux I__6853 (
            .O(N__30699),
            .I(N__30691));
    CascadeMux I__6852 (
            .O(N__30698),
            .I(N__30688));
    LocalMux I__6851 (
            .O(N__30695),
            .I(N__30685));
    CascadeMux I__6850 (
            .O(N__30694),
            .I(N__30680));
    LocalMux I__6849 (
            .O(N__30691),
            .I(N__30673));
    InMux I__6848 (
            .O(N__30688),
            .I(N__30670));
    Span4Mux_s3_h I__6847 (
            .O(N__30685),
            .I(N__30667));
    InMux I__6846 (
            .O(N__30684),
            .I(N__30662));
    InMux I__6845 (
            .O(N__30683),
            .I(N__30662));
    InMux I__6844 (
            .O(N__30680),
            .I(N__30659));
    InMux I__6843 (
            .O(N__30679),
            .I(N__30654));
    InMux I__6842 (
            .O(N__30678),
            .I(N__30654));
    InMux I__6841 (
            .O(N__30677),
            .I(N__30649));
    InMux I__6840 (
            .O(N__30676),
            .I(N__30649));
    Span4Mux_h I__6839 (
            .O(N__30673),
            .I(N__30646));
    LocalMux I__6838 (
            .O(N__30670),
            .I(N__30643));
    Sp12to4 I__6837 (
            .O(N__30667),
            .I(N__30638));
    LocalMux I__6836 (
            .O(N__30662),
            .I(N__30638));
    LocalMux I__6835 (
            .O(N__30659),
            .I(N__30631));
    LocalMux I__6834 (
            .O(N__30654),
            .I(N__30631));
    LocalMux I__6833 (
            .O(N__30649),
            .I(N__30631));
    Span4Mux_h I__6832 (
            .O(N__30646),
            .I(N__30628));
    Sp12to4 I__6831 (
            .O(N__30643),
            .I(N__30625));
    Span12Mux_s7_v I__6830 (
            .O(N__30638),
            .I(N__30620));
    Span12Mux_s3_h I__6829 (
            .O(N__30631),
            .I(N__30620));
    Odrv4 I__6828 (
            .O(N__30628),
            .I(\POWERLED.N_335 ));
    Odrv12 I__6827 (
            .O(N__30625),
            .I(\POWERLED.N_335 ));
    Odrv12 I__6826 (
            .O(N__30620),
            .I(\POWERLED.N_335 ));
    InMux I__6825 (
            .O(N__30613),
            .I(N__30607));
    InMux I__6824 (
            .O(N__30612),
            .I(N__30607));
    LocalMux I__6823 (
            .O(N__30607),
            .I(N_22_0));
    CascadeMux I__6822 (
            .O(N__30604),
            .I(N_22_0_cascade_));
    InMux I__6821 (
            .O(N__30601),
            .I(N__30597));
    CascadeMux I__6820 (
            .O(N__30600),
            .I(N__30593));
    LocalMux I__6819 (
            .O(N__30597),
            .I(N__30590));
    InMux I__6818 (
            .O(N__30596),
            .I(N__30585));
    InMux I__6817 (
            .O(N__30593),
            .I(N__30585));
    Span4Mux_s0_h I__6816 (
            .O(N__30590),
            .I(N__30580));
    LocalMux I__6815 (
            .O(N__30585),
            .I(N__30580));
    Odrv4 I__6814 (
            .O(N__30580),
            .I(N_2145_i));
    InMux I__6813 (
            .O(N__30577),
            .I(N__30574));
    LocalMux I__6812 (
            .O(N__30574),
            .I(g0_0_1));
    InMux I__6811 (
            .O(N__30571),
            .I(N__30565));
    InMux I__6810 (
            .O(N__30570),
            .I(N__30560));
    InMux I__6809 (
            .O(N__30569),
            .I(N__30560));
    InMux I__6808 (
            .O(N__30568),
            .I(N__30557));
    LocalMux I__6807 (
            .O(N__30565),
            .I(N__30552));
    LocalMux I__6806 (
            .O(N__30560),
            .I(N__30541));
    LocalMux I__6805 (
            .O(N__30557),
            .I(N__30541));
    InMux I__6804 (
            .O(N__30556),
            .I(N__30538));
    InMux I__6803 (
            .O(N__30555),
            .I(N__30535));
    Span4Mux_v I__6802 (
            .O(N__30552),
            .I(N__30529));
    InMux I__6801 (
            .O(N__30551),
            .I(N__30524));
    InMux I__6800 (
            .O(N__30550),
            .I(N__30515));
    InMux I__6799 (
            .O(N__30549),
            .I(N__30515));
    InMux I__6798 (
            .O(N__30548),
            .I(N__30515));
    InMux I__6797 (
            .O(N__30547),
            .I(N__30510));
    InMux I__6796 (
            .O(N__30546),
            .I(N__30510));
    Span4Mux_v I__6795 (
            .O(N__30541),
            .I(N__30505));
    LocalMux I__6794 (
            .O(N__30538),
            .I(N__30505));
    LocalMux I__6793 (
            .O(N__30535),
            .I(N__30502));
    InMux I__6792 (
            .O(N__30534),
            .I(N__30499));
    InMux I__6791 (
            .O(N__30533),
            .I(N__30494));
    InMux I__6790 (
            .O(N__30532),
            .I(N__30494));
    IoSpan4Mux I__6789 (
            .O(N__30529),
            .I(N__30491));
    InMux I__6788 (
            .O(N__30528),
            .I(N__30488));
    InMux I__6787 (
            .O(N__30527),
            .I(N__30485));
    LocalMux I__6786 (
            .O(N__30524),
            .I(N__30482));
    InMux I__6785 (
            .O(N__30523),
            .I(N__30479));
    InMux I__6784 (
            .O(N__30522),
            .I(N__30476));
    LocalMux I__6783 (
            .O(N__30515),
            .I(N__30470));
    LocalMux I__6782 (
            .O(N__30510),
            .I(N__30470));
    Span4Mux_h I__6781 (
            .O(N__30505),
            .I(N__30466));
    Span4Mux_v I__6780 (
            .O(N__30502),
            .I(N__30459));
    LocalMux I__6779 (
            .O(N__30499),
            .I(N__30459));
    LocalMux I__6778 (
            .O(N__30494),
            .I(N__30459));
    Span4Mux_s3_h I__6777 (
            .O(N__30491),
            .I(N__30452));
    LocalMux I__6776 (
            .O(N__30488),
            .I(N__30452));
    LocalMux I__6775 (
            .O(N__30485),
            .I(N__30452));
    Span4Mux_h I__6774 (
            .O(N__30482),
            .I(N__30444));
    LocalMux I__6773 (
            .O(N__30479),
            .I(N__30444));
    LocalMux I__6772 (
            .O(N__30476),
            .I(N__30444));
    InMux I__6771 (
            .O(N__30475),
            .I(N__30441));
    Span4Mux_v I__6770 (
            .O(N__30470),
            .I(N__30438));
    InMux I__6769 (
            .O(N__30469),
            .I(N__30435));
    Span4Mux_h I__6768 (
            .O(N__30466),
            .I(N__30430));
    Span4Mux_h I__6767 (
            .O(N__30459),
            .I(N__30430));
    Span4Mux_h I__6766 (
            .O(N__30452),
            .I(N__30427));
    InMux I__6765 (
            .O(N__30451),
            .I(N__30424));
    Span4Mux_h I__6764 (
            .O(N__30444),
            .I(N__30419));
    LocalMux I__6763 (
            .O(N__30441),
            .I(N__30419));
    Span4Mux_s3_v I__6762 (
            .O(N__30438),
            .I(N__30414));
    LocalMux I__6761 (
            .O(N__30435),
            .I(N__30414));
    Span4Mux_v I__6760 (
            .O(N__30430),
            .I(N__30411));
    Span4Mux_v I__6759 (
            .O(N__30427),
            .I(N__30408));
    LocalMux I__6758 (
            .O(N__30424),
            .I(N__30405));
    Span4Mux_v I__6757 (
            .O(N__30419),
            .I(N__30400));
    Span4Mux_h I__6756 (
            .O(N__30414),
            .I(N__30400));
    Odrv4 I__6755 (
            .O(N__30411),
            .I(slp_s4n));
    Odrv4 I__6754 (
            .O(N__30408),
            .I(slp_s4n));
    Odrv12 I__6753 (
            .O(N__30405),
            .I(slp_s4n));
    Odrv4 I__6752 (
            .O(N__30400),
            .I(slp_s4n));
    CascadeMux I__6751 (
            .O(N__30391),
            .I(N__30388));
    InMux I__6750 (
            .O(N__30388),
            .I(N__30377));
    CascadeMux I__6749 (
            .O(N__30387),
            .I(N__30368));
    CascadeMux I__6748 (
            .O(N__30386),
            .I(N__30362));
    CascadeMux I__6747 (
            .O(N__30385),
            .I(N__30359));
    CascadeMux I__6746 (
            .O(N__30384),
            .I(N__30355));
    InMux I__6745 (
            .O(N__30383),
            .I(N__30347));
    InMux I__6744 (
            .O(N__30382),
            .I(N__30347));
    InMux I__6743 (
            .O(N__30381),
            .I(N__30347));
    CascadeMux I__6742 (
            .O(N__30380),
            .I(N__30344));
    LocalMux I__6741 (
            .O(N__30377),
            .I(N__30341));
    InMux I__6740 (
            .O(N__30376),
            .I(N__30338));
    InMux I__6739 (
            .O(N__30375),
            .I(N__30333));
    InMux I__6738 (
            .O(N__30374),
            .I(N__30333));
    InMux I__6737 (
            .O(N__30373),
            .I(N__30328));
    InMux I__6736 (
            .O(N__30372),
            .I(N__30328));
    InMux I__6735 (
            .O(N__30371),
            .I(N__30325));
    InMux I__6734 (
            .O(N__30368),
            .I(N__30316));
    InMux I__6733 (
            .O(N__30367),
            .I(N__30316));
    InMux I__6732 (
            .O(N__30366),
            .I(N__30316));
    InMux I__6731 (
            .O(N__30365),
            .I(N__30316));
    InMux I__6730 (
            .O(N__30362),
            .I(N__30311));
    InMux I__6729 (
            .O(N__30359),
            .I(N__30311));
    InMux I__6728 (
            .O(N__30358),
            .I(N__30308));
    InMux I__6727 (
            .O(N__30355),
            .I(N__30305));
    InMux I__6726 (
            .O(N__30354),
            .I(N__30302));
    LocalMux I__6725 (
            .O(N__30347),
            .I(N__30299));
    InMux I__6724 (
            .O(N__30344),
            .I(N__30296));
    Span4Mux_s3_h I__6723 (
            .O(N__30341),
            .I(N__30292));
    LocalMux I__6722 (
            .O(N__30338),
            .I(N__30289));
    LocalMux I__6721 (
            .O(N__30333),
            .I(N__30284));
    LocalMux I__6720 (
            .O(N__30328),
            .I(N__30284));
    LocalMux I__6719 (
            .O(N__30325),
            .I(N__30277));
    LocalMux I__6718 (
            .O(N__30316),
            .I(N__30277));
    LocalMux I__6717 (
            .O(N__30311),
            .I(N__30277));
    LocalMux I__6716 (
            .O(N__30308),
            .I(N__30269));
    LocalMux I__6715 (
            .O(N__30305),
            .I(N__30269));
    LocalMux I__6714 (
            .O(N__30302),
            .I(N__30262));
    Span4Mux_h I__6713 (
            .O(N__30299),
            .I(N__30262));
    LocalMux I__6712 (
            .O(N__30296),
            .I(N__30262));
    InMux I__6711 (
            .O(N__30295),
            .I(N__30259));
    Span4Mux_h I__6710 (
            .O(N__30292),
            .I(N__30250));
    Span4Mux_h I__6709 (
            .O(N__30289),
            .I(N__30250));
    Span4Mux_v I__6708 (
            .O(N__30284),
            .I(N__30250));
    Span4Mux_v I__6707 (
            .O(N__30277),
            .I(N__30250));
    InMux I__6706 (
            .O(N__30276),
            .I(N__30245));
    InMux I__6705 (
            .O(N__30275),
            .I(N__30245));
    CascadeMux I__6704 (
            .O(N__30274),
            .I(N__30240));
    Span4Mux_v I__6703 (
            .O(N__30269),
            .I(N__30233));
    Span4Mux_v I__6702 (
            .O(N__30262),
            .I(N__30233));
    LocalMux I__6701 (
            .O(N__30259),
            .I(N__30233));
    Span4Mux_h I__6700 (
            .O(N__30250),
            .I(N__30228));
    LocalMux I__6699 (
            .O(N__30245),
            .I(N__30228));
    InMux I__6698 (
            .O(N__30244),
            .I(N__30225));
    InMux I__6697 (
            .O(N__30243),
            .I(N__30222));
    InMux I__6696 (
            .O(N__30240),
            .I(N__30219));
    Span4Mux_h I__6695 (
            .O(N__30233),
            .I(N__30214));
    IoSpan4Mux I__6694 (
            .O(N__30228),
            .I(N__30211));
    LocalMux I__6693 (
            .O(N__30225),
            .I(N__30206));
    LocalMux I__6692 (
            .O(N__30222),
            .I(N__30206));
    LocalMux I__6691 (
            .O(N__30219),
            .I(N__30203));
    InMux I__6690 (
            .O(N__30218),
            .I(N__30198));
    InMux I__6689 (
            .O(N__30217),
            .I(N__30198));
    IoSpan4Mux I__6688 (
            .O(N__30214),
            .I(N__30195));
    IoSpan4Mux I__6687 (
            .O(N__30211),
            .I(N__30192));
    Span12Mux_s10_h I__6686 (
            .O(N__30206),
            .I(N__30185));
    Span12Mux_s1_h I__6685 (
            .O(N__30203),
            .I(N__30185));
    LocalMux I__6684 (
            .O(N__30198),
            .I(N__30185));
    Odrv4 I__6683 (
            .O(N__30195),
            .I(slp_s3n));
    Odrv4 I__6682 (
            .O(N__30192),
            .I(slp_s3n));
    Odrv12 I__6681 (
            .O(N__30185),
            .I(slp_s3n));
    CascadeMux I__6680 (
            .O(N__30178),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_4_cascade_ ));
    InMux I__6679 (
            .O(N__30175),
            .I(N__30172));
    LocalMux I__6678 (
            .O(N__30172),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_4 ));
    CascadeMux I__6677 (
            .O(N__30169),
            .I(\POWERLED.o2_cascade_ ));
    InMux I__6676 (
            .O(N__30166),
            .I(N__30163));
    LocalMux I__6675 (
            .O(N__30163),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_10 ));
    CascadeMux I__6674 (
            .O(N__30160),
            .I(N__30154));
    InMux I__6673 (
            .O(N__30159),
            .I(N__30150));
    InMux I__6672 (
            .O(N__30158),
            .I(N__30140));
    InMux I__6671 (
            .O(N__30157),
            .I(N__30137));
    InMux I__6670 (
            .O(N__30154),
            .I(N__30134));
    InMux I__6669 (
            .O(N__30153),
            .I(N__30131));
    LocalMux I__6668 (
            .O(N__30150),
            .I(N__30128));
    InMux I__6667 (
            .O(N__30149),
            .I(N__30123));
    InMux I__6666 (
            .O(N__30148),
            .I(N__30123));
    CascadeMux I__6665 (
            .O(N__30147),
            .I(N__30120));
    CascadeMux I__6664 (
            .O(N__30146),
            .I(N__30110));
    CascadeMux I__6663 (
            .O(N__30145),
            .I(N__30105));
    InMux I__6662 (
            .O(N__30144),
            .I(N__30101));
    InMux I__6661 (
            .O(N__30143),
            .I(N__30098));
    LocalMux I__6660 (
            .O(N__30140),
            .I(N__30095));
    LocalMux I__6659 (
            .O(N__30137),
            .I(N__30092));
    LocalMux I__6658 (
            .O(N__30134),
            .I(N__30089));
    LocalMux I__6657 (
            .O(N__30131),
            .I(N__30082));
    Span4Mux_v I__6656 (
            .O(N__30128),
            .I(N__30082));
    LocalMux I__6655 (
            .O(N__30123),
            .I(N__30082));
    InMux I__6654 (
            .O(N__30120),
            .I(N__30077));
    InMux I__6653 (
            .O(N__30119),
            .I(N__30077));
    InMux I__6652 (
            .O(N__30118),
            .I(N__30074));
    InMux I__6651 (
            .O(N__30117),
            .I(N__30069));
    InMux I__6650 (
            .O(N__30116),
            .I(N__30069));
    InMux I__6649 (
            .O(N__30115),
            .I(N__30062));
    InMux I__6648 (
            .O(N__30114),
            .I(N__30062));
    InMux I__6647 (
            .O(N__30113),
            .I(N__30062));
    InMux I__6646 (
            .O(N__30110),
            .I(N__30057));
    InMux I__6645 (
            .O(N__30109),
            .I(N__30057));
    InMux I__6644 (
            .O(N__30108),
            .I(N__30050));
    InMux I__6643 (
            .O(N__30105),
            .I(N__30050));
    InMux I__6642 (
            .O(N__30104),
            .I(N__30050));
    LocalMux I__6641 (
            .O(N__30101),
            .I(N__30045));
    LocalMux I__6640 (
            .O(N__30098),
            .I(N__30045));
    Span4Mux_v I__6639 (
            .O(N__30095),
            .I(N__30038));
    Span4Mux_v I__6638 (
            .O(N__30092),
            .I(N__30038));
    Span4Mux_v I__6637 (
            .O(N__30089),
            .I(N__30038));
    Odrv4 I__6636 (
            .O(N__30082),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__6635 (
            .O(N__30077),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__6634 (
            .O(N__30074),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__6633 (
            .O(N__30069),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__6632 (
            .O(N__30062),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__6631 (
            .O(N__30057),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__6630 (
            .O(N__30050),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__6629 (
            .O(N__30045),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__6628 (
            .O(N__30038),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    CascadeMux I__6627 (
            .O(N__30019),
            .I(N__30014));
    CascadeMux I__6626 (
            .O(N__30018),
            .I(N__30010));
    CascadeMux I__6625 (
            .O(N__30017),
            .I(N__30007));
    InMux I__6624 (
            .O(N__30014),
            .I(N__30000));
    CascadeMux I__6623 (
            .O(N__30013),
            .I(N__29994));
    InMux I__6622 (
            .O(N__30010),
            .I(N__29990));
    InMux I__6621 (
            .O(N__30007),
            .I(N__29985));
    InMux I__6620 (
            .O(N__30006),
            .I(N__29985));
    CascadeMux I__6619 (
            .O(N__30005),
            .I(N__29982));
    InMux I__6618 (
            .O(N__30004),
            .I(N__29979));
    InMux I__6617 (
            .O(N__30003),
            .I(N__29975));
    LocalMux I__6616 (
            .O(N__30000),
            .I(N__29972));
    InMux I__6615 (
            .O(N__29999),
            .I(N__29968));
    InMux I__6614 (
            .O(N__29998),
            .I(N__29958));
    InMux I__6613 (
            .O(N__29997),
            .I(N__29958));
    InMux I__6612 (
            .O(N__29994),
            .I(N__29958));
    CascadeMux I__6611 (
            .O(N__29993),
            .I(N__29955));
    LocalMux I__6610 (
            .O(N__29990),
            .I(N__29949));
    LocalMux I__6609 (
            .O(N__29985),
            .I(N__29949));
    InMux I__6608 (
            .O(N__29982),
            .I(N__29946));
    LocalMux I__6607 (
            .O(N__29979),
            .I(N__29943));
    InMux I__6606 (
            .O(N__29978),
            .I(N__29940));
    LocalMux I__6605 (
            .O(N__29975),
            .I(N__29937));
    Span4Mux_v I__6604 (
            .O(N__29972),
            .I(N__29934));
    InMux I__6603 (
            .O(N__29971),
            .I(N__29931));
    LocalMux I__6602 (
            .O(N__29968),
            .I(N__29928));
    InMux I__6601 (
            .O(N__29967),
            .I(N__29921));
    InMux I__6600 (
            .O(N__29966),
            .I(N__29921));
    InMux I__6599 (
            .O(N__29965),
            .I(N__29921));
    LocalMux I__6598 (
            .O(N__29958),
            .I(N__29918));
    InMux I__6597 (
            .O(N__29955),
            .I(N__29913));
    InMux I__6596 (
            .O(N__29954),
            .I(N__29913));
    Span4Mux_v I__6595 (
            .O(N__29949),
            .I(N__29908));
    LocalMux I__6594 (
            .O(N__29946),
            .I(N__29908));
    Odrv12 I__6593 (
            .O(N__29943),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__6592 (
            .O(N__29940),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__6591 (
            .O(N__29937),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__6590 (
            .O(N__29934),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__6589 (
            .O(N__29931),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__6588 (
            .O(N__29928),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__6587 (
            .O(N__29921),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__6586 (
            .O(N__29918),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__6585 (
            .O(N__29913),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__6584 (
            .O(N__29908),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    CascadeMux I__6583 (
            .O(N__29887),
            .I(N__29876));
    CascadeMux I__6582 (
            .O(N__29886),
            .I(N__29873));
    CascadeMux I__6581 (
            .O(N__29885),
            .I(N__29865));
    CascadeMux I__6580 (
            .O(N__29884),
            .I(N__29860));
    CascadeMux I__6579 (
            .O(N__29883),
            .I(N__29857));
    InMux I__6578 (
            .O(N__29882),
            .I(N__29849));
    InMux I__6577 (
            .O(N__29881),
            .I(N__29849));
    InMux I__6576 (
            .O(N__29880),
            .I(N__29849));
    InMux I__6575 (
            .O(N__29879),
            .I(N__29846));
    InMux I__6574 (
            .O(N__29876),
            .I(N__29843));
    InMux I__6573 (
            .O(N__29873),
            .I(N__29838));
    InMux I__6572 (
            .O(N__29872),
            .I(N__29838));
    InMux I__6571 (
            .O(N__29871),
            .I(N__29835));
    InMux I__6570 (
            .O(N__29870),
            .I(N__29832));
    CascadeMux I__6569 (
            .O(N__29869),
            .I(N__29819));
    CascadeMux I__6568 (
            .O(N__29868),
            .I(N__29816));
    InMux I__6567 (
            .O(N__29865),
            .I(N__29812));
    InMux I__6566 (
            .O(N__29864),
            .I(N__29809));
    InMux I__6565 (
            .O(N__29863),
            .I(N__29802));
    InMux I__6564 (
            .O(N__29860),
            .I(N__29802));
    InMux I__6563 (
            .O(N__29857),
            .I(N__29802));
    InMux I__6562 (
            .O(N__29856),
            .I(N__29799));
    LocalMux I__6561 (
            .O(N__29849),
            .I(N__29796));
    LocalMux I__6560 (
            .O(N__29846),
            .I(N__29793));
    LocalMux I__6559 (
            .O(N__29843),
            .I(N__29789));
    LocalMux I__6558 (
            .O(N__29838),
            .I(N__29782));
    LocalMux I__6557 (
            .O(N__29835),
            .I(N__29782));
    LocalMux I__6556 (
            .O(N__29832),
            .I(N__29782));
    InMux I__6555 (
            .O(N__29831),
            .I(N__29775));
    InMux I__6554 (
            .O(N__29830),
            .I(N__29775));
    InMux I__6553 (
            .O(N__29829),
            .I(N__29775));
    InMux I__6552 (
            .O(N__29828),
            .I(N__29772));
    InMux I__6551 (
            .O(N__29827),
            .I(N__29767));
    InMux I__6550 (
            .O(N__29826),
            .I(N__29767));
    InMux I__6549 (
            .O(N__29825),
            .I(N__29760));
    InMux I__6548 (
            .O(N__29824),
            .I(N__29760));
    InMux I__6547 (
            .O(N__29823),
            .I(N__29760));
    InMux I__6546 (
            .O(N__29822),
            .I(N__29753));
    InMux I__6545 (
            .O(N__29819),
            .I(N__29753));
    InMux I__6544 (
            .O(N__29816),
            .I(N__29753));
    CascadeMux I__6543 (
            .O(N__29815),
            .I(N__29749));
    LocalMux I__6542 (
            .O(N__29812),
            .I(N__29745));
    LocalMux I__6541 (
            .O(N__29809),
            .I(N__29740));
    LocalMux I__6540 (
            .O(N__29802),
            .I(N__29740));
    LocalMux I__6539 (
            .O(N__29799),
            .I(N__29737));
    Span4Mux_s2_h I__6538 (
            .O(N__29796),
            .I(N__29734));
    Span4Mux_s2_h I__6537 (
            .O(N__29793),
            .I(N__29731));
    InMux I__6536 (
            .O(N__29792),
            .I(N__29728));
    Span4Mux_v I__6535 (
            .O(N__29789),
            .I(N__29723));
    Span4Mux_v I__6534 (
            .O(N__29782),
            .I(N__29723));
    LocalMux I__6533 (
            .O(N__29775),
            .I(N__29712));
    LocalMux I__6532 (
            .O(N__29772),
            .I(N__29712));
    LocalMux I__6531 (
            .O(N__29767),
            .I(N__29712));
    LocalMux I__6530 (
            .O(N__29760),
            .I(N__29712));
    LocalMux I__6529 (
            .O(N__29753),
            .I(N__29712));
    InMux I__6528 (
            .O(N__29752),
            .I(N__29705));
    InMux I__6527 (
            .O(N__29749),
            .I(N__29705));
    InMux I__6526 (
            .O(N__29748),
            .I(N__29705));
    Span4Mux_h I__6525 (
            .O(N__29745),
            .I(N__29700));
    Span4Mux_s2_h I__6524 (
            .O(N__29740),
            .I(N__29700));
    Odrv12 I__6523 (
            .O(N__29737),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__6522 (
            .O(N__29734),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__6521 (
            .O(N__29731),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__6520 (
            .O(N__29728),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__6519 (
            .O(N__29723),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv12 I__6518 (
            .O(N__29712),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__6517 (
            .O(N__29705),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__6516 (
            .O(N__29700),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    CascadeMux I__6515 (
            .O(N__29683),
            .I(N__29678));
    CascadeMux I__6514 (
            .O(N__29682),
            .I(N__29668));
    InMux I__6513 (
            .O(N__29681),
            .I(N__29662));
    InMux I__6512 (
            .O(N__29678),
            .I(N__29662));
    InMux I__6511 (
            .O(N__29677),
            .I(N__29652));
    InMux I__6510 (
            .O(N__29676),
            .I(N__29652));
    InMux I__6509 (
            .O(N__29675),
            .I(N__29652));
    CascadeMux I__6508 (
            .O(N__29674),
            .I(N__29649));
    InMux I__6507 (
            .O(N__29673),
            .I(N__29640));
    InMux I__6506 (
            .O(N__29672),
            .I(N__29640));
    InMux I__6505 (
            .O(N__29671),
            .I(N__29640));
    InMux I__6504 (
            .O(N__29668),
            .I(N__29636));
    CascadeMux I__6503 (
            .O(N__29667),
            .I(N__29632));
    LocalMux I__6502 (
            .O(N__29662),
            .I(N__29628));
    InMux I__6501 (
            .O(N__29661),
            .I(N__29623));
    InMux I__6500 (
            .O(N__29660),
            .I(N__29623));
    InMux I__6499 (
            .O(N__29659),
            .I(N__29620));
    LocalMux I__6498 (
            .O(N__29652),
            .I(N__29617));
    InMux I__6497 (
            .O(N__29649),
            .I(N__29597));
    InMux I__6496 (
            .O(N__29648),
            .I(N__29597));
    InMux I__6495 (
            .O(N__29647),
            .I(N__29597));
    LocalMux I__6494 (
            .O(N__29640),
            .I(N__29594));
    InMux I__6493 (
            .O(N__29639),
            .I(N__29591));
    LocalMux I__6492 (
            .O(N__29636),
            .I(N__29588));
    InMux I__6491 (
            .O(N__29635),
            .I(N__29583));
    InMux I__6490 (
            .O(N__29632),
            .I(N__29583));
    InMux I__6489 (
            .O(N__29631),
            .I(N__29580));
    Span4Mux_v I__6488 (
            .O(N__29628),
            .I(N__29571));
    LocalMux I__6487 (
            .O(N__29623),
            .I(N__29571));
    LocalMux I__6486 (
            .O(N__29620),
            .I(N__29571));
    Span4Mux_v I__6485 (
            .O(N__29617),
            .I(N__29571));
    InMux I__6484 (
            .O(N__29616),
            .I(N__29568));
    InMux I__6483 (
            .O(N__29615),
            .I(N__29561));
    InMux I__6482 (
            .O(N__29614),
            .I(N__29561));
    InMux I__6481 (
            .O(N__29613),
            .I(N__29561));
    InMux I__6480 (
            .O(N__29612),
            .I(N__29552));
    InMux I__6479 (
            .O(N__29611),
            .I(N__29552));
    InMux I__6478 (
            .O(N__29610),
            .I(N__29552));
    InMux I__6477 (
            .O(N__29609),
            .I(N__29552));
    InMux I__6476 (
            .O(N__29608),
            .I(N__29545));
    InMux I__6475 (
            .O(N__29607),
            .I(N__29545));
    InMux I__6474 (
            .O(N__29606),
            .I(N__29545));
    InMux I__6473 (
            .O(N__29605),
            .I(N__29540));
    InMux I__6472 (
            .O(N__29604),
            .I(N__29540));
    LocalMux I__6471 (
            .O(N__29597),
            .I(N__29537));
    Span4Mux_s1_h I__6470 (
            .O(N__29594),
            .I(N__29530));
    LocalMux I__6469 (
            .O(N__29591),
            .I(N__29530));
    Span4Mux_h I__6468 (
            .O(N__29588),
            .I(N__29530));
    LocalMux I__6467 (
            .O(N__29583),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__6466 (
            .O(N__29580),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__6465 (
            .O(N__29571),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__6464 (
            .O(N__29568),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__6463 (
            .O(N__29561),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__6462 (
            .O(N__29552),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__6461 (
            .O(N__29545),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__6460 (
            .O(N__29540),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv12 I__6459 (
            .O(N__29537),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__6458 (
            .O(N__29530),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    InMux I__6457 (
            .O(N__29509),
            .I(N__29503));
    InMux I__6456 (
            .O(N__29508),
            .I(N__29503));
    LocalMux I__6455 (
            .O(N__29503),
            .I(N__29499));
    CascadeMux I__6454 (
            .O(N__29502),
            .I(N__29496));
    Span4Mux_v I__6453 (
            .O(N__29499),
            .I(N__29493));
    InMux I__6452 (
            .O(N__29496),
            .I(N__29490));
    Odrv4 I__6451 (
            .O(N__29493),
            .I(\POWERLED.N_2191_i ));
    LocalMux I__6450 (
            .O(N__29490),
            .I(\POWERLED.N_2191_i ));
    CascadeMux I__6449 (
            .O(N__29485),
            .I(N__29480));
    InMux I__6448 (
            .O(N__29484),
            .I(N__29472));
    InMux I__6447 (
            .O(N__29483),
            .I(N__29469));
    InMux I__6446 (
            .O(N__29480),
            .I(N__29466));
    InMux I__6445 (
            .O(N__29479),
            .I(N__29460));
    InMux I__6444 (
            .O(N__29478),
            .I(N__29460));
    CascadeMux I__6443 (
            .O(N__29477),
            .I(N__29457));
    InMux I__6442 (
            .O(N__29476),
            .I(N__29454));
    InMux I__6441 (
            .O(N__29475),
            .I(N__29450));
    LocalMux I__6440 (
            .O(N__29472),
            .I(N__29445));
    LocalMux I__6439 (
            .O(N__29469),
            .I(N__29445));
    LocalMux I__6438 (
            .O(N__29466),
            .I(N__29442));
    InMux I__6437 (
            .O(N__29465),
            .I(N__29439));
    LocalMux I__6436 (
            .O(N__29460),
            .I(N__29434));
    InMux I__6435 (
            .O(N__29457),
            .I(N__29431));
    LocalMux I__6434 (
            .O(N__29454),
            .I(N__29428));
    InMux I__6433 (
            .O(N__29453),
            .I(N__29425));
    LocalMux I__6432 (
            .O(N__29450),
            .I(N__29420));
    Span4Mux_h I__6431 (
            .O(N__29445),
            .I(N__29420));
    Span4Mux_s1_h I__6430 (
            .O(N__29442),
            .I(N__29415));
    LocalMux I__6429 (
            .O(N__29439),
            .I(N__29415));
    InMux I__6428 (
            .O(N__29438),
            .I(N__29410));
    InMux I__6427 (
            .O(N__29437),
            .I(N__29410));
    Span4Mux_v I__6426 (
            .O(N__29434),
            .I(N__29405));
    LocalMux I__6425 (
            .O(N__29431),
            .I(N__29405));
    Span4Mux_s0_h I__6424 (
            .O(N__29428),
            .I(N__29402));
    LocalMux I__6423 (
            .O(N__29425),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv4 I__6422 (
            .O(N__29420),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv4 I__6421 (
            .O(N__29415),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__6420 (
            .O(N__29410),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv4 I__6419 (
            .O(N__29405),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv4 I__6418 (
            .O(N__29402),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    InMux I__6417 (
            .O(N__29389),
            .I(N__29385));
    CascadeMux I__6416 (
            .O(N__29388),
            .I(N__29382));
    LocalMux I__6415 (
            .O(N__29385),
            .I(N__29378));
    InMux I__6414 (
            .O(N__29382),
            .I(N__29372));
    InMux I__6413 (
            .O(N__29381),
            .I(N__29372));
    Span4Mux_v I__6412 (
            .O(N__29378),
            .I(N__29369));
    InMux I__6411 (
            .O(N__29377),
            .I(N__29366));
    LocalMux I__6410 (
            .O(N__29372),
            .I(N__29363));
    Span4Mux_h I__6409 (
            .O(N__29369),
            .I(N__29360));
    LocalMux I__6408 (
            .O(N__29366),
            .I(N__29357));
    Span4Mux_h I__6407 (
            .O(N__29363),
            .I(N__29354));
    Odrv4 I__6406 (
            .O(N__29360),
            .I(\POWERLED.N_2187_i ));
    Odrv12 I__6405 (
            .O(N__29357),
            .I(\POWERLED.N_2187_i ));
    Odrv4 I__6404 (
            .O(N__29354),
            .I(\POWERLED.N_2187_i ));
    CascadeMux I__6403 (
            .O(N__29347),
            .I(\POWERLED.un2_count_clk_17_0_0_a2_5_cascade_ ));
    InMux I__6402 (
            .O(N__29344),
            .I(N__29341));
    LocalMux I__6401 (
            .O(N__29341),
            .I(\POWERLED.un2_count_clk_17_0_0_a2_0 ));
    InMux I__6400 (
            .O(N__29338),
            .I(N__29335));
    LocalMux I__6399 (
            .O(N__29335),
            .I(N__29331));
    CascadeMux I__6398 (
            .O(N__29334),
            .I(N__29328));
    Span4Mux_h I__6397 (
            .O(N__29331),
            .I(N__29324));
    InMux I__6396 (
            .O(N__29328),
            .I(N__29321));
    InMux I__6395 (
            .O(N__29327),
            .I(N__29318));
    Span4Mux_h I__6394 (
            .O(N__29324),
            .I(N__29315));
    LocalMux I__6393 (
            .O(N__29321),
            .I(\POWERLED.N_501 ));
    LocalMux I__6392 (
            .O(N__29318),
            .I(\POWERLED.N_501 ));
    Odrv4 I__6391 (
            .O(N__29315),
            .I(\POWERLED.N_501 ));
    InMux I__6390 (
            .O(N__29308),
            .I(N__29299));
    InMux I__6389 (
            .O(N__29307),
            .I(N__29299));
    InMux I__6388 (
            .O(N__29306),
            .I(N__29289));
    CascadeMux I__6387 (
            .O(N__29305),
            .I(N__29286));
    CascadeMux I__6386 (
            .O(N__29304),
            .I(N__29282));
    LocalMux I__6385 (
            .O(N__29299),
            .I(N__29279));
    InMux I__6384 (
            .O(N__29298),
            .I(N__29274));
    InMux I__6383 (
            .O(N__29297),
            .I(N__29274));
    CascadeMux I__6382 (
            .O(N__29296),
            .I(N__29270));
    CascadeMux I__6381 (
            .O(N__29295),
            .I(N__29267));
    InMux I__6380 (
            .O(N__29294),
            .I(N__29262));
    InMux I__6379 (
            .O(N__29293),
            .I(N__29262));
    CascadeMux I__6378 (
            .O(N__29292),
            .I(N__29258));
    LocalMux I__6377 (
            .O(N__29289),
            .I(N__29253));
    InMux I__6376 (
            .O(N__29286),
            .I(N__29250));
    CascadeMux I__6375 (
            .O(N__29285),
            .I(N__29246));
    InMux I__6374 (
            .O(N__29282),
            .I(N__29242));
    Span4Mux_s0_h I__6373 (
            .O(N__29279),
            .I(N__29239));
    LocalMux I__6372 (
            .O(N__29274),
            .I(N__29236));
    InMux I__6371 (
            .O(N__29273),
            .I(N__29233));
    InMux I__6370 (
            .O(N__29270),
            .I(N__29228));
    InMux I__6369 (
            .O(N__29267),
            .I(N__29228));
    LocalMux I__6368 (
            .O(N__29262),
            .I(N__29225));
    CascadeMux I__6367 (
            .O(N__29261),
            .I(N__29221));
    InMux I__6366 (
            .O(N__29258),
            .I(N__29218));
    InMux I__6365 (
            .O(N__29257),
            .I(N__29215));
    InMux I__6364 (
            .O(N__29256),
            .I(N__29212));
    Span4Mux_v I__6363 (
            .O(N__29253),
            .I(N__29207));
    LocalMux I__6362 (
            .O(N__29250),
            .I(N__29207));
    InMux I__6361 (
            .O(N__29249),
            .I(N__29200));
    InMux I__6360 (
            .O(N__29246),
            .I(N__29200));
    InMux I__6359 (
            .O(N__29245),
            .I(N__29200));
    LocalMux I__6358 (
            .O(N__29242),
            .I(N__29195));
    Span4Mux_h I__6357 (
            .O(N__29239),
            .I(N__29195));
    Span4Mux_s3_h I__6356 (
            .O(N__29236),
            .I(N__29192));
    LocalMux I__6355 (
            .O(N__29233),
            .I(N__29187));
    LocalMux I__6354 (
            .O(N__29228),
            .I(N__29187));
    Span4Mux_s3_h I__6353 (
            .O(N__29225),
            .I(N__29184));
    InMux I__6352 (
            .O(N__29224),
            .I(N__29179));
    InMux I__6351 (
            .O(N__29221),
            .I(N__29179));
    LocalMux I__6350 (
            .O(N__29218),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__6349 (
            .O(N__29215),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__6348 (
            .O(N__29212),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__6347 (
            .O(N__29207),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__6346 (
            .O(N__29200),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__6345 (
            .O(N__29195),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__6344 (
            .O(N__29192),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv12 I__6343 (
            .O(N__29187),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__6342 (
            .O(N__29184),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__6341 (
            .O(N__29179),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    InMux I__6340 (
            .O(N__29158),
            .I(N__29146));
    InMux I__6339 (
            .O(N__29157),
            .I(N__29146));
    CascadeMux I__6338 (
            .O(N__29156),
            .I(N__29142));
    CascadeMux I__6337 (
            .O(N__29155),
            .I(N__29133));
    CascadeMux I__6336 (
            .O(N__29154),
            .I(N__29124));
    CascadeMux I__6335 (
            .O(N__29153),
            .I(N__29119));
    InMux I__6334 (
            .O(N__29152),
            .I(N__29114));
    InMux I__6333 (
            .O(N__29151),
            .I(N__29114));
    LocalMux I__6332 (
            .O(N__29146),
            .I(N__29111));
    InMux I__6331 (
            .O(N__29145),
            .I(N__29104));
    InMux I__6330 (
            .O(N__29142),
            .I(N__29104));
    InMux I__6329 (
            .O(N__29141),
            .I(N__29104));
    InMux I__6328 (
            .O(N__29140),
            .I(N__29093));
    InMux I__6327 (
            .O(N__29139),
            .I(N__29093));
    InMux I__6326 (
            .O(N__29138),
            .I(N__29093));
    InMux I__6325 (
            .O(N__29137),
            .I(N__29093));
    InMux I__6324 (
            .O(N__29136),
            .I(N__29090));
    InMux I__6323 (
            .O(N__29133),
            .I(N__29087));
    InMux I__6322 (
            .O(N__29132),
            .I(N__29080));
    InMux I__6321 (
            .O(N__29131),
            .I(N__29080));
    InMux I__6320 (
            .O(N__29130),
            .I(N__29080));
    InMux I__6319 (
            .O(N__29129),
            .I(N__29076));
    InMux I__6318 (
            .O(N__29128),
            .I(N__29071));
    InMux I__6317 (
            .O(N__29127),
            .I(N__29060));
    InMux I__6316 (
            .O(N__29124),
            .I(N__29060));
    InMux I__6315 (
            .O(N__29123),
            .I(N__29060));
    InMux I__6314 (
            .O(N__29122),
            .I(N__29060));
    InMux I__6313 (
            .O(N__29119),
            .I(N__29060));
    LocalMux I__6312 (
            .O(N__29114),
            .I(N__29055));
    Span4Mux_v I__6311 (
            .O(N__29111),
            .I(N__29055));
    LocalMux I__6310 (
            .O(N__29104),
            .I(N__29052));
    InMux I__6309 (
            .O(N__29103),
            .I(N__29049));
    InMux I__6308 (
            .O(N__29102),
            .I(N__29046));
    LocalMux I__6307 (
            .O(N__29093),
            .I(N__29043));
    LocalMux I__6306 (
            .O(N__29090),
            .I(N__29038));
    LocalMux I__6305 (
            .O(N__29087),
            .I(N__29038));
    LocalMux I__6304 (
            .O(N__29080),
            .I(N__29035));
    InMux I__6303 (
            .O(N__29079),
            .I(N__29032));
    LocalMux I__6302 (
            .O(N__29076),
            .I(N__29028));
    InMux I__6301 (
            .O(N__29075),
            .I(N__29022));
    InMux I__6300 (
            .O(N__29074),
            .I(N__29022));
    LocalMux I__6299 (
            .O(N__29071),
            .I(N__29017));
    LocalMux I__6298 (
            .O(N__29060),
            .I(N__29017));
    Span4Mux_v I__6297 (
            .O(N__29055),
            .I(N__29012));
    Span4Mux_v I__6296 (
            .O(N__29052),
            .I(N__29012));
    LocalMux I__6295 (
            .O(N__29049),
            .I(N__28999));
    LocalMux I__6294 (
            .O(N__29046),
            .I(N__28999));
    Span4Mux_v I__6293 (
            .O(N__29043),
            .I(N__28999));
    Span4Mux_v I__6292 (
            .O(N__29038),
            .I(N__28999));
    Span4Mux_s1_h I__6291 (
            .O(N__29035),
            .I(N__28999));
    LocalMux I__6290 (
            .O(N__29032),
            .I(N__28999));
    InMux I__6289 (
            .O(N__29031),
            .I(N__28996));
    Span4Mux_v I__6288 (
            .O(N__29028),
            .I(N__28993));
    InMux I__6287 (
            .O(N__29027),
            .I(N__28990));
    LocalMux I__6286 (
            .O(N__29022),
            .I(N__28985));
    Span4Mux_v I__6285 (
            .O(N__29017),
            .I(N__28985));
    Span4Mux_h I__6284 (
            .O(N__29012),
            .I(N__28982));
    Span4Mux_h I__6283 (
            .O(N__28999),
            .I(N__28979));
    LocalMux I__6282 (
            .O(N__28996),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__6281 (
            .O(N__28993),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__6280 (
            .O(N__28990),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__6279 (
            .O(N__28985),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__6278 (
            .O(N__28982),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__6277 (
            .O(N__28979),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    InMux I__6276 (
            .O(N__28966),
            .I(N__28959));
    InMux I__6275 (
            .O(N__28965),
            .I(N__28954));
    InMux I__6274 (
            .O(N__28964),
            .I(N__28954));
    InMux I__6273 (
            .O(N__28963),
            .I(N__28945));
    InMux I__6272 (
            .O(N__28962),
            .I(N__28945));
    LocalMux I__6271 (
            .O(N__28959),
            .I(N__28938));
    LocalMux I__6270 (
            .O(N__28954),
            .I(N__28938));
    InMux I__6269 (
            .O(N__28953),
            .I(N__28933));
    InMux I__6268 (
            .O(N__28952),
            .I(N__28933));
    InMux I__6267 (
            .O(N__28951),
            .I(N__28930));
    InMux I__6266 (
            .O(N__28950),
            .I(N__28927));
    LocalMux I__6265 (
            .O(N__28945),
            .I(N__28924));
    CascadeMux I__6264 (
            .O(N__28944),
            .I(N__28919));
    InMux I__6263 (
            .O(N__28943),
            .I(N__28916));
    Span4Mux_v I__6262 (
            .O(N__28938),
            .I(N__28913));
    LocalMux I__6261 (
            .O(N__28933),
            .I(N__28910));
    LocalMux I__6260 (
            .O(N__28930),
            .I(N__28902));
    LocalMux I__6259 (
            .O(N__28927),
            .I(N__28902));
    Span4Mux_v I__6258 (
            .O(N__28924),
            .I(N__28902));
    InMux I__6257 (
            .O(N__28923),
            .I(N__28895));
    InMux I__6256 (
            .O(N__28922),
            .I(N__28895));
    InMux I__6255 (
            .O(N__28919),
            .I(N__28895));
    LocalMux I__6254 (
            .O(N__28916),
            .I(N__28892));
    Span4Mux_v I__6253 (
            .O(N__28913),
            .I(N__28887));
    Span4Mux_v I__6252 (
            .O(N__28910),
            .I(N__28887));
    InMux I__6251 (
            .O(N__28909),
            .I(N__28884));
    Span4Mux_h I__6250 (
            .O(N__28902),
            .I(N__28881));
    LocalMux I__6249 (
            .O(N__28895),
            .I(N__28876));
    Span4Mux_h I__6248 (
            .O(N__28892),
            .I(N__28876));
    Span4Mux_h I__6247 (
            .O(N__28887),
            .I(N__28873));
    LocalMux I__6246 (
            .O(N__28884),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__6245 (
            .O(N__28881),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__6244 (
            .O(N__28876),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__6243 (
            .O(N__28873),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    CascadeMux I__6242 (
            .O(N__28864),
            .I(N__28852));
    InMux I__6241 (
            .O(N__28863),
            .I(N__28845));
    InMux I__6240 (
            .O(N__28862),
            .I(N__28845));
    InMux I__6239 (
            .O(N__28861),
            .I(N__28838));
    InMux I__6238 (
            .O(N__28860),
            .I(N__28838));
    CascadeMux I__6237 (
            .O(N__28859),
            .I(N__28835));
    InMux I__6236 (
            .O(N__28858),
            .I(N__28831));
    InMux I__6235 (
            .O(N__28857),
            .I(N__28826));
    InMux I__6234 (
            .O(N__28856),
            .I(N__28821));
    InMux I__6233 (
            .O(N__28855),
            .I(N__28821));
    InMux I__6232 (
            .O(N__28852),
            .I(N__28808));
    InMux I__6231 (
            .O(N__28851),
            .I(N__28808));
    InMux I__6230 (
            .O(N__28850),
            .I(N__28808));
    LocalMux I__6229 (
            .O(N__28845),
            .I(N__28805));
    InMux I__6228 (
            .O(N__28844),
            .I(N__28800));
    InMux I__6227 (
            .O(N__28843),
            .I(N__28800));
    LocalMux I__6226 (
            .O(N__28838),
            .I(N__28797));
    InMux I__6225 (
            .O(N__28835),
            .I(N__28794));
    InMux I__6224 (
            .O(N__28834),
            .I(N__28791));
    LocalMux I__6223 (
            .O(N__28831),
            .I(N__28788));
    CascadeMux I__6222 (
            .O(N__28830),
            .I(N__28785));
    CascadeMux I__6221 (
            .O(N__28829),
            .I(N__28781));
    LocalMux I__6220 (
            .O(N__28826),
            .I(N__28775));
    LocalMux I__6219 (
            .O(N__28821),
            .I(N__28775));
    InMux I__6218 (
            .O(N__28820),
            .I(N__28772));
    InMux I__6217 (
            .O(N__28819),
            .I(N__28769));
    InMux I__6216 (
            .O(N__28818),
            .I(N__28762));
    InMux I__6215 (
            .O(N__28817),
            .I(N__28762));
    InMux I__6214 (
            .O(N__28816),
            .I(N__28762));
    InMux I__6213 (
            .O(N__28815),
            .I(N__28753));
    LocalMux I__6212 (
            .O(N__28808),
            .I(N__28746));
    Span4Mux_s2_h I__6211 (
            .O(N__28805),
            .I(N__28746));
    LocalMux I__6210 (
            .O(N__28800),
            .I(N__28746));
    Span12Mux_s6_h I__6209 (
            .O(N__28797),
            .I(N__28743));
    LocalMux I__6208 (
            .O(N__28794),
            .I(N__28738));
    LocalMux I__6207 (
            .O(N__28791),
            .I(N__28738));
    Span4Mux_v I__6206 (
            .O(N__28788),
            .I(N__28735));
    InMux I__6205 (
            .O(N__28785),
            .I(N__28732));
    InMux I__6204 (
            .O(N__28784),
            .I(N__28729));
    InMux I__6203 (
            .O(N__28781),
            .I(N__28726));
    InMux I__6202 (
            .O(N__28780),
            .I(N__28723));
    Span4Mux_h I__6201 (
            .O(N__28775),
            .I(N__28720));
    LocalMux I__6200 (
            .O(N__28772),
            .I(N__28713));
    LocalMux I__6199 (
            .O(N__28769),
            .I(N__28713));
    LocalMux I__6198 (
            .O(N__28762),
            .I(N__28713));
    InMux I__6197 (
            .O(N__28761),
            .I(N__28706));
    InMux I__6196 (
            .O(N__28760),
            .I(N__28706));
    InMux I__6195 (
            .O(N__28759),
            .I(N__28706));
    InMux I__6194 (
            .O(N__28758),
            .I(N__28699));
    InMux I__6193 (
            .O(N__28757),
            .I(N__28699));
    InMux I__6192 (
            .O(N__28756),
            .I(N__28699));
    LocalMux I__6191 (
            .O(N__28753),
            .I(N__28694));
    Span4Mux_h I__6190 (
            .O(N__28746),
            .I(N__28694));
    Odrv12 I__6189 (
            .O(N__28743),
            .I(func_state_RNITGMHB_0_1));
    Odrv4 I__6188 (
            .O(N__28738),
            .I(func_state_RNITGMHB_0_1));
    Odrv4 I__6187 (
            .O(N__28735),
            .I(func_state_RNITGMHB_0_1));
    LocalMux I__6186 (
            .O(N__28732),
            .I(func_state_RNITGMHB_0_1));
    LocalMux I__6185 (
            .O(N__28729),
            .I(func_state_RNITGMHB_0_1));
    LocalMux I__6184 (
            .O(N__28726),
            .I(func_state_RNITGMHB_0_1));
    LocalMux I__6183 (
            .O(N__28723),
            .I(func_state_RNITGMHB_0_1));
    Odrv4 I__6182 (
            .O(N__28720),
            .I(func_state_RNITGMHB_0_1));
    Odrv12 I__6181 (
            .O(N__28713),
            .I(func_state_RNITGMHB_0_1));
    LocalMux I__6180 (
            .O(N__28706),
            .I(func_state_RNITGMHB_0_1));
    LocalMux I__6179 (
            .O(N__28699),
            .I(func_state_RNITGMHB_0_1));
    Odrv4 I__6178 (
            .O(N__28694),
            .I(func_state_RNITGMHB_0_1));
    CascadeMux I__6177 (
            .O(N__28669),
            .I(N__28665));
    InMux I__6176 (
            .O(N__28668),
            .I(N__28660));
    InMux I__6175 (
            .O(N__28665),
            .I(N__28660));
    LocalMux I__6174 (
            .O(N__28660),
            .I(\POWERLED.un2_count_clk_17_0_1 ));
    CascadeMux I__6173 (
            .O(N__28657),
            .I(\POWERLED.un2_count_clk_17_0_1_cascade_ ));
    CascadeMux I__6172 (
            .O(N__28654),
            .I(N__28650));
    InMux I__6171 (
            .O(N__28653),
            .I(N__28647));
    InMux I__6170 (
            .O(N__28650),
            .I(N__28644));
    LocalMux I__6169 (
            .O(N__28647),
            .I(N__28636));
    LocalMux I__6168 (
            .O(N__28644),
            .I(N__28633));
    InMux I__6167 (
            .O(N__28643),
            .I(N__28630));
    InMux I__6166 (
            .O(N__28642),
            .I(N__28627));
    InMux I__6165 (
            .O(N__28641),
            .I(N__28624));
    InMux I__6164 (
            .O(N__28640),
            .I(N__28621));
    InMux I__6163 (
            .O(N__28639),
            .I(N__28618));
    Span4Mux_s0_h I__6162 (
            .O(N__28636),
            .I(N__28615));
    Odrv4 I__6161 (
            .O(N__28633),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__6160 (
            .O(N__28630),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__6159 (
            .O(N__28627),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__6158 (
            .O(N__28624),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__6157 (
            .O(N__28621),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__6156 (
            .O(N__28618),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    Odrv4 I__6155 (
            .O(N__28615),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    InMux I__6154 (
            .O(N__28600),
            .I(N__28594));
    InMux I__6153 (
            .O(N__28599),
            .I(N__28591));
    InMux I__6152 (
            .O(N__28598),
            .I(N__28583));
    InMux I__6151 (
            .O(N__28597),
            .I(N__28580));
    LocalMux I__6150 (
            .O(N__28594),
            .I(N__28575));
    LocalMux I__6149 (
            .O(N__28591),
            .I(N__28575));
    InMux I__6148 (
            .O(N__28590),
            .I(N__28572));
    InMux I__6147 (
            .O(N__28589),
            .I(N__28569));
    InMux I__6146 (
            .O(N__28588),
            .I(N__28566));
    CascadeMux I__6145 (
            .O(N__28587),
            .I(N__28560));
    CascadeMux I__6144 (
            .O(N__28586),
            .I(N__28556));
    LocalMux I__6143 (
            .O(N__28583),
            .I(N__28546));
    LocalMux I__6142 (
            .O(N__28580),
            .I(N__28546));
    Span4Mux_s1_h I__6141 (
            .O(N__28575),
            .I(N__28546));
    LocalMux I__6140 (
            .O(N__28572),
            .I(N__28539));
    LocalMux I__6139 (
            .O(N__28569),
            .I(N__28539));
    LocalMux I__6138 (
            .O(N__28566),
            .I(N__28539));
    InMux I__6137 (
            .O(N__28565),
            .I(N__28534));
    InMux I__6136 (
            .O(N__28564),
            .I(N__28534));
    InMux I__6135 (
            .O(N__28563),
            .I(N__28529));
    InMux I__6134 (
            .O(N__28560),
            .I(N__28529));
    InMux I__6133 (
            .O(N__28559),
            .I(N__28524));
    InMux I__6132 (
            .O(N__28556),
            .I(N__28524));
    InMux I__6131 (
            .O(N__28555),
            .I(N__28521));
    InMux I__6130 (
            .O(N__28554),
            .I(N__28518));
    InMux I__6129 (
            .O(N__28553),
            .I(N__28515));
    Span4Mux_v I__6128 (
            .O(N__28546),
            .I(N__28512));
    Span12Mux_s4_h I__6127 (
            .O(N__28539),
            .I(N__28505));
    LocalMux I__6126 (
            .O(N__28534),
            .I(N__28505));
    LocalMux I__6125 (
            .O(N__28529),
            .I(N__28505));
    LocalMux I__6124 (
            .O(N__28524),
            .I(N__28502));
    LocalMux I__6123 (
            .O(N__28521),
            .I(POWERLED_func_state_0_sqmuxa));
    LocalMux I__6122 (
            .O(N__28518),
            .I(POWERLED_func_state_0_sqmuxa));
    LocalMux I__6121 (
            .O(N__28515),
            .I(POWERLED_func_state_0_sqmuxa));
    Odrv4 I__6120 (
            .O(N__28512),
            .I(POWERLED_func_state_0_sqmuxa));
    Odrv12 I__6119 (
            .O(N__28505),
            .I(POWERLED_func_state_0_sqmuxa));
    Odrv4 I__6118 (
            .O(N__28502),
            .I(POWERLED_func_state_0_sqmuxa));
    CascadeMux I__6117 (
            .O(N__28489),
            .I(\POWERLED.N_2191_i_cascade_ ));
    InMux I__6116 (
            .O(N__28486),
            .I(N__28476));
    InMux I__6115 (
            .O(N__28485),
            .I(N__28476));
    InMux I__6114 (
            .O(N__28484),
            .I(N__28473));
    CascadeMux I__6113 (
            .O(N__28483),
            .I(N__28470));
    InMux I__6112 (
            .O(N__28482),
            .I(N__28465));
    InMux I__6111 (
            .O(N__28481),
            .I(N__28462));
    LocalMux I__6110 (
            .O(N__28476),
            .I(N__28458));
    LocalMux I__6109 (
            .O(N__28473),
            .I(N__28454));
    InMux I__6108 (
            .O(N__28470),
            .I(N__28449));
    InMux I__6107 (
            .O(N__28469),
            .I(N__28449));
    InMux I__6106 (
            .O(N__28468),
            .I(N__28446));
    LocalMux I__6105 (
            .O(N__28465),
            .I(N__28443));
    LocalMux I__6104 (
            .O(N__28462),
            .I(N__28440));
    InMux I__6103 (
            .O(N__28461),
            .I(N__28437));
    Span4Mux_v I__6102 (
            .O(N__28458),
            .I(N__28432));
    InMux I__6101 (
            .O(N__28457),
            .I(N__28429));
    Span4Mux_v I__6100 (
            .O(N__28454),
            .I(N__28424));
    LocalMux I__6099 (
            .O(N__28449),
            .I(N__28424));
    LocalMux I__6098 (
            .O(N__28446),
            .I(N__28421));
    Span4Mux_s0_h I__6097 (
            .O(N__28443),
            .I(N__28414));
    Span4Mux_v I__6096 (
            .O(N__28440),
            .I(N__28414));
    LocalMux I__6095 (
            .O(N__28437),
            .I(N__28414));
    InMux I__6094 (
            .O(N__28436),
            .I(N__28411));
    InMux I__6093 (
            .O(N__28435),
            .I(N__28408));
    Span4Mux_v I__6092 (
            .O(N__28432),
            .I(N__28405));
    LocalMux I__6091 (
            .O(N__28429),
            .I(N__28400));
    Span4Mux_h I__6090 (
            .O(N__28424),
            .I(N__28400));
    Span4Mux_h I__6089 (
            .O(N__28421),
            .I(N__28395));
    Span4Mux_h I__6088 (
            .O(N__28414),
            .I(N__28395));
    LocalMux I__6087 (
            .O(N__28411),
            .I(\POWERLED.N_282_N ));
    LocalMux I__6086 (
            .O(N__28408),
            .I(\POWERLED.N_282_N ));
    Odrv4 I__6085 (
            .O(N__28405),
            .I(\POWERLED.N_282_N ));
    Odrv4 I__6084 (
            .O(N__28400),
            .I(\POWERLED.N_282_N ));
    Odrv4 I__6083 (
            .O(N__28395),
            .I(\POWERLED.N_282_N ));
    InMux I__6082 (
            .O(N__28384),
            .I(N__28378));
    InMux I__6081 (
            .O(N__28383),
            .I(N__28378));
    LocalMux I__6080 (
            .O(N__28378),
            .I(N__28375));
    Odrv12 I__6079 (
            .O(N__28375),
            .I(\POWERLED.dutycycle_eena_12 ));
    InMux I__6078 (
            .O(N__28372),
            .I(N__28369));
    LocalMux I__6077 (
            .O(N__28369),
            .I(\POWERLED.g0_i_i_a6_0_2 ));
    CascadeMux I__6076 (
            .O(N__28366),
            .I(N__28363));
    InMux I__6075 (
            .O(N__28363),
            .I(N__28360));
    LocalMux I__6074 (
            .O(N__28360),
            .I(\POWERLED.dutycycle_RNIZ0Z_4 ));
    CascadeMux I__6073 (
            .O(N__28357),
            .I(N__28352));
    InMux I__6072 (
            .O(N__28356),
            .I(N__28348));
    CascadeMux I__6071 (
            .O(N__28355),
            .I(N__28345));
    InMux I__6070 (
            .O(N__28352),
            .I(N__28340));
    InMux I__6069 (
            .O(N__28351),
            .I(N__28340));
    LocalMux I__6068 (
            .O(N__28348),
            .I(N__28337));
    InMux I__6067 (
            .O(N__28345),
            .I(N__28334));
    LocalMux I__6066 (
            .O(N__28340),
            .I(N__28331));
    Span4Mux_v I__6065 (
            .O(N__28337),
            .I(N__28325));
    LocalMux I__6064 (
            .O(N__28334),
            .I(N__28322));
    Span4Mux_h I__6063 (
            .O(N__28331),
            .I(N__28319));
    InMux I__6062 (
            .O(N__28330),
            .I(N__28312));
    InMux I__6061 (
            .O(N__28329),
            .I(N__28312));
    InMux I__6060 (
            .O(N__28328),
            .I(N__28312));
    Odrv4 I__6059 (
            .O(N__28325),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    Odrv4 I__6058 (
            .O(N__28322),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    Odrv4 I__6057 (
            .O(N__28319),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__6056 (
            .O(N__28312),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    CascadeMux I__6055 (
            .O(N__28303),
            .I(N__28300));
    InMux I__6054 (
            .O(N__28300),
            .I(N__28297));
    LocalMux I__6053 (
            .O(N__28297),
            .I(\POWERLED.g0_i_i_1 ));
    InMux I__6052 (
            .O(N__28294),
            .I(N__28291));
    LocalMux I__6051 (
            .O(N__28291),
            .I(\POWERLED.un1_dutycycle_53_axb_11_1 ));
    CascadeMux I__6050 (
            .O(N__28288),
            .I(N__28285));
    InMux I__6049 (
            .O(N__28285),
            .I(N__28282));
    LocalMux I__6048 (
            .O(N__28282),
            .I(N__28279));
    Span4Mux_h I__6047 (
            .O(N__28279),
            .I(N__28276));
    Span4Mux_h I__6046 (
            .O(N__28276),
            .I(N__28273));
    Odrv4 I__6045 (
            .O(N__28273),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_14 ));
    InMux I__6044 (
            .O(N__28270),
            .I(N__28263));
    InMux I__6043 (
            .O(N__28269),
            .I(N__28263));
    InMux I__6042 (
            .O(N__28268),
            .I(N__28260));
    LocalMux I__6041 (
            .O(N__28263),
            .I(N__28257));
    LocalMux I__6040 (
            .O(N__28260),
            .I(N__28254));
    Span4Mux_s2_h I__6039 (
            .O(N__28257),
            .I(N__28251));
    Span4Mux_v I__6038 (
            .O(N__28254),
            .I(N__28248));
    Span4Mux_v I__6037 (
            .O(N__28251),
            .I(N__28245));
    Odrv4 I__6036 (
            .O(N__28248),
            .I(\POWERLED.N_2293_i ));
    Odrv4 I__6035 (
            .O(N__28245),
            .I(\POWERLED.N_2293_i ));
    InMux I__6034 (
            .O(N__28240),
            .I(N__28237));
    LocalMux I__6033 (
            .O(N__28237),
            .I(\POWERLED.un1_dutycycle_53_4_1 ));
    CascadeMux I__6032 (
            .O(N__28234),
            .I(N__28231));
    InMux I__6031 (
            .O(N__28231),
            .I(N__28225));
    InMux I__6030 (
            .O(N__28230),
            .I(N__28225));
    LocalMux I__6029 (
            .O(N__28225),
            .I(N__28222));
    Span4Mux_v I__6028 (
            .O(N__28222),
            .I(N__28219));
    Odrv4 I__6027 (
            .O(N__28219),
            .I(\POWERLED.dutycycle_eena_10 ));
    InMux I__6026 (
            .O(N__28216),
            .I(N__28212));
    InMux I__6025 (
            .O(N__28215),
            .I(N__28209));
    LocalMux I__6024 (
            .O(N__28212),
            .I(N__28206));
    LocalMux I__6023 (
            .O(N__28209),
            .I(N__28202));
    Span4Mux_v I__6022 (
            .O(N__28206),
            .I(N__28199));
    InMux I__6021 (
            .O(N__28205),
            .I(N__28195));
    Span4Mux_v I__6020 (
            .O(N__28202),
            .I(N__28190));
    Span4Mux_h I__6019 (
            .O(N__28199),
            .I(N__28190));
    InMux I__6018 (
            .O(N__28198),
            .I(N__28187));
    LocalMux I__6017 (
            .O(N__28195),
            .I(\POWERLED.N_507 ));
    Odrv4 I__6016 (
            .O(N__28190),
            .I(\POWERLED.N_507 ));
    LocalMux I__6015 (
            .O(N__28187),
            .I(\POWERLED.N_507 ));
    CascadeMux I__6014 (
            .O(N__28180),
            .I(\POWERLED.N_84_f0_cascade_ ));
    CascadeMux I__6013 (
            .O(N__28177),
            .I(N__28171));
    IoInMux I__6012 (
            .O(N__28176),
            .I(N__28166));
    CascadeMux I__6011 (
            .O(N__28175),
            .I(N__28163));
    CascadeMux I__6010 (
            .O(N__28174),
            .I(N__28160));
    InMux I__6009 (
            .O(N__28171),
            .I(N__28156));
    CascadeMux I__6008 (
            .O(N__28170),
            .I(N__28152));
    CascadeMux I__6007 (
            .O(N__28169),
            .I(N__28144));
    LocalMux I__6006 (
            .O(N__28166),
            .I(N__28137));
    InMux I__6005 (
            .O(N__28163),
            .I(N__28130));
    InMux I__6004 (
            .O(N__28160),
            .I(N__28130));
    InMux I__6003 (
            .O(N__28159),
            .I(N__28130));
    LocalMux I__6002 (
            .O(N__28156),
            .I(N__28127));
    InMux I__6001 (
            .O(N__28155),
            .I(N__28118));
    InMux I__6000 (
            .O(N__28152),
            .I(N__28118));
    InMux I__5999 (
            .O(N__28151),
            .I(N__28118));
    InMux I__5998 (
            .O(N__28150),
            .I(N__28118));
    InMux I__5997 (
            .O(N__28149),
            .I(N__28115));
    CascadeMux I__5996 (
            .O(N__28148),
            .I(N__28112));
    CascadeMux I__5995 (
            .O(N__28147),
            .I(N__28108));
    InMux I__5994 (
            .O(N__28144),
            .I(N__28100));
    InMux I__5993 (
            .O(N__28143),
            .I(N__28100));
    InMux I__5992 (
            .O(N__28142),
            .I(N__28097));
    InMux I__5991 (
            .O(N__28141),
            .I(N__28092));
    InMux I__5990 (
            .O(N__28140),
            .I(N__28092));
    IoSpan4Mux I__5989 (
            .O(N__28137),
            .I(N__28088));
    LocalMux I__5988 (
            .O(N__28130),
            .I(N__28085));
    Span4Mux_v I__5987 (
            .O(N__28127),
            .I(N__28080));
    LocalMux I__5986 (
            .O(N__28118),
            .I(N__28080));
    LocalMux I__5985 (
            .O(N__28115),
            .I(N__28077));
    InMux I__5984 (
            .O(N__28112),
            .I(N__28072));
    InMux I__5983 (
            .O(N__28111),
            .I(N__28072));
    InMux I__5982 (
            .O(N__28108),
            .I(N__28069));
    CascadeMux I__5981 (
            .O(N__28107),
            .I(N__28064));
    CascadeMux I__5980 (
            .O(N__28106),
            .I(N__28061));
    CascadeMux I__5979 (
            .O(N__28105),
            .I(N__28058));
    LocalMux I__5978 (
            .O(N__28100),
            .I(N__28055));
    LocalMux I__5977 (
            .O(N__28097),
            .I(N__28052));
    LocalMux I__5976 (
            .O(N__28092),
            .I(N__28049));
    InMux I__5975 (
            .O(N__28091),
            .I(N__28046));
    Span4Mux_s1_h I__5974 (
            .O(N__28088),
            .I(N__28043));
    Span4Mux_v I__5973 (
            .O(N__28085),
            .I(N__28040));
    Span4Mux_v I__5972 (
            .O(N__28080),
            .I(N__28036));
    Span4Mux_s1_h I__5971 (
            .O(N__28077),
            .I(N__28031));
    LocalMux I__5970 (
            .O(N__28072),
            .I(N__28031));
    LocalMux I__5969 (
            .O(N__28069),
            .I(N__28022));
    InMux I__5968 (
            .O(N__28068),
            .I(N__28017));
    InMux I__5967 (
            .O(N__28067),
            .I(N__28017));
    InMux I__5966 (
            .O(N__28064),
            .I(N__28012));
    InMux I__5965 (
            .O(N__28061),
            .I(N__28012));
    InMux I__5964 (
            .O(N__28058),
            .I(N__28008));
    Span4Mux_h I__5963 (
            .O(N__28055),
            .I(N__28005));
    Span12Mux_s9_v I__5962 (
            .O(N__28052),
            .I(N__28002));
    Span4Mux_h I__5961 (
            .O(N__28049),
            .I(N__27997));
    LocalMux I__5960 (
            .O(N__28046),
            .I(N__27997));
    Span4Mux_h I__5959 (
            .O(N__28043),
            .I(N__27992));
    Span4Mux_v I__5958 (
            .O(N__28040),
            .I(N__27992));
    InMux I__5957 (
            .O(N__28039),
            .I(N__27989));
    Span4Mux_s1_h I__5956 (
            .O(N__28036),
            .I(N__27984));
    Span4Mux_v I__5955 (
            .O(N__28031),
            .I(N__27984));
    InMux I__5954 (
            .O(N__28030),
            .I(N__27981));
    InMux I__5953 (
            .O(N__28029),
            .I(N__27976));
    InMux I__5952 (
            .O(N__28028),
            .I(N__27976));
    InMux I__5951 (
            .O(N__28027),
            .I(N__27969));
    InMux I__5950 (
            .O(N__28026),
            .I(N__27969));
    InMux I__5949 (
            .O(N__28025),
            .I(N__27969));
    Span4Mux_v I__5948 (
            .O(N__28022),
            .I(N__27962));
    LocalMux I__5947 (
            .O(N__28017),
            .I(N__27962));
    LocalMux I__5946 (
            .O(N__28012),
            .I(N__27962));
    InMux I__5945 (
            .O(N__28011),
            .I(N__27959));
    LocalMux I__5944 (
            .O(N__28008),
            .I(G_156));
    Odrv4 I__5943 (
            .O(N__28005),
            .I(G_156));
    Odrv12 I__5942 (
            .O(N__28002),
            .I(G_156));
    Odrv4 I__5941 (
            .O(N__27997),
            .I(G_156));
    Odrv4 I__5940 (
            .O(N__27992),
            .I(G_156));
    LocalMux I__5939 (
            .O(N__27989),
            .I(G_156));
    Odrv4 I__5938 (
            .O(N__27984),
            .I(G_156));
    LocalMux I__5937 (
            .O(N__27981),
            .I(G_156));
    LocalMux I__5936 (
            .O(N__27976),
            .I(G_156));
    LocalMux I__5935 (
            .O(N__27969),
            .I(G_156));
    Odrv4 I__5934 (
            .O(N__27962),
            .I(G_156));
    LocalMux I__5933 (
            .O(N__27959),
            .I(G_156));
    InMux I__5932 (
            .O(N__27934),
            .I(N__27928));
    InMux I__5931 (
            .O(N__27933),
            .I(N__27928));
    LocalMux I__5930 (
            .O(N__27928),
            .I(\POWERLED.dutycycle_en_3 ));
    InMux I__5929 (
            .O(N__27925),
            .I(N__27922));
    LocalMux I__5928 (
            .O(N__27922),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_11 ));
    CascadeMux I__5927 (
            .O(N__27919),
            .I(\POWERLED.N_12_cascade_ ));
    CascadeMux I__5926 (
            .O(N__27916),
            .I(N__27909));
    CascadeMux I__5925 (
            .O(N__27915),
            .I(N__27906));
    InMux I__5924 (
            .O(N__27914),
            .I(N__27902));
    InMux I__5923 (
            .O(N__27913),
            .I(N__27897));
    InMux I__5922 (
            .O(N__27912),
            .I(N__27897));
    InMux I__5921 (
            .O(N__27909),
            .I(N__27892));
    InMux I__5920 (
            .O(N__27906),
            .I(N__27892));
    InMux I__5919 (
            .O(N__27905),
            .I(N__27889));
    LocalMux I__5918 (
            .O(N__27902),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_3 ));
    LocalMux I__5917 (
            .O(N__27897),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_3 ));
    LocalMux I__5916 (
            .O(N__27892),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_3 ));
    LocalMux I__5915 (
            .O(N__27889),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_3 ));
    InMux I__5914 (
            .O(N__27880),
            .I(N__27877));
    LocalMux I__5913 (
            .O(N__27877),
            .I(N__27874));
    Odrv12 I__5912 (
            .O(N__27874),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_4 ));
    InMux I__5911 (
            .O(N__27871),
            .I(N__27866));
    CascadeMux I__5910 (
            .O(N__27870),
            .I(N__27863));
    CascadeMux I__5909 (
            .O(N__27869),
            .I(N__27860));
    LocalMux I__5908 (
            .O(N__27866),
            .I(N__27857));
    InMux I__5907 (
            .O(N__27863),
            .I(N__27852));
    InMux I__5906 (
            .O(N__27860),
            .I(N__27852));
    Span4Mux_v I__5905 (
            .O(N__27857),
            .I(N__27847));
    LocalMux I__5904 (
            .O(N__27852),
            .I(N__27847));
    Odrv4 I__5903 (
            .O(N__27847),
            .I(\POWERLED.un1_dutycycle_53_25_0_tz ));
    InMux I__5902 (
            .O(N__27844),
            .I(N__27841));
    LocalMux I__5901 (
            .O(N__27841),
            .I(\POWERLED.N_6 ));
    SRMux I__5900 (
            .O(N__27838),
            .I(N__27835));
    LocalMux I__5899 (
            .O(N__27835),
            .I(N__27832));
    Span4Mux_v I__5898 (
            .O(N__27832),
            .I(N__27829));
    Odrv4 I__5897 (
            .O(N__27829),
            .I(\VPP_VDDQ.N_28_i ));
    InMux I__5896 (
            .O(N__27826),
            .I(N__27819));
    InMux I__5895 (
            .O(N__27825),
            .I(N__27819));
    InMux I__5894 (
            .O(N__27824),
            .I(N__27816));
    LocalMux I__5893 (
            .O(N__27819),
            .I(\VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0 ));
    LocalMux I__5892 (
            .O(N__27816),
            .I(\VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0 ));
    CascadeMux I__5891 (
            .O(N__27811),
            .I(N__27807));
    CascadeMux I__5890 (
            .O(N__27810),
            .I(N__27804));
    InMux I__5889 (
            .O(N__27807),
            .I(N__27799));
    InMux I__5888 (
            .O(N__27804),
            .I(N__27799));
    LocalMux I__5887 (
            .O(N__27799),
            .I(\VPP_VDDQ.delayed_vddq_okZ0 ));
    InMux I__5886 (
            .O(N__27796),
            .I(N__27790));
    InMux I__5885 (
            .O(N__27795),
            .I(N__27790));
    LocalMux I__5884 (
            .O(N__27790),
            .I(\VPP_VDDQ.delayed_vddq_ok_en ));
    InMux I__5883 (
            .O(N__27787),
            .I(N__27784));
    LocalMux I__5882 (
            .O(N__27784),
            .I(N__27781));
    Odrv12 I__5881 (
            .O(N__27781),
            .I(VPP_VDDQ_delayed_vddq_ok));
    CascadeMux I__5880 (
            .O(N__27778),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_9_cascade_ ));
    InMux I__5879 (
            .O(N__27775),
            .I(N__27772));
    LocalMux I__5878 (
            .O(N__27772),
            .I(N__27769));
    Odrv12 I__5877 (
            .O(N__27769),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_9 ));
    InMux I__5876 (
            .O(N__27766),
            .I(N__27763));
    LocalMux I__5875 (
            .O(N__27763),
            .I(\POWERLED.un1_dutycycle_53_4_a0_1 ));
    CascadeMux I__5874 (
            .O(N__27760),
            .I(\POWERLED.un1_dutycycle_53_4_a0_1_cascade_ ));
    InMux I__5873 (
            .O(N__27757),
            .I(N__27754));
    LocalMux I__5872 (
            .O(N__27754),
            .I(N__27751));
    Odrv4 I__5871 (
            .O(N__27751),
            .I(\POWERLED.un1_dutycycle_53_7_2 ));
    InMux I__5870 (
            .O(N__27748),
            .I(N__27745));
    LocalMux I__5869 (
            .O(N__27745),
            .I(\POWERLED.un1_dutycycle_53_8_1 ));
    CascadeMux I__5868 (
            .O(N__27742),
            .I(\POWERLED.un1_dutycycle_53_8_1_cascade_ ));
    InMux I__5867 (
            .O(N__27739),
            .I(N__27736));
    LocalMux I__5866 (
            .O(N__27736),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_9 ));
    InMux I__5865 (
            .O(N__27733),
            .I(N__27730));
    LocalMux I__5864 (
            .O(N__27730),
            .I(N__27727));
    Odrv12 I__5863 (
            .O(N__27727),
            .I(\POWERLED.dutycycle_RNIZ0Z_5 ));
    InMux I__5862 (
            .O(N__27724),
            .I(N__27721));
    LocalMux I__5861 (
            .O(N__27721),
            .I(\VPP_VDDQ.curr_state_2_0_0 ));
    CascadeMux I__5860 (
            .O(N__27718),
            .I(\VPP_VDDQ.N_190_cascade_ ));
    InMux I__5859 (
            .O(N__27715),
            .I(N__27712));
    LocalMux I__5858 (
            .O(N__27712),
            .I(N__27708));
    InMux I__5857 (
            .O(N__27711),
            .I(N__27705));
    Span4Mux_s3_v I__5856 (
            .O(N__27708),
            .I(N__27702));
    LocalMux I__5855 (
            .O(N__27705),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ));
    Odrv4 I__5854 (
            .O(N__27702),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ));
    CascadeMux I__5853 (
            .O(N__27697),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ));
    InMux I__5852 (
            .O(N__27694),
            .I(N__27691));
    LocalMux I__5851 (
            .O(N__27691),
            .I(N__27688));
    Span4Mux_s3_v I__5850 (
            .O(N__27688),
            .I(N__27685));
    Odrv4 I__5849 (
            .O(N__27685),
            .I(\VPP_VDDQ.count_2_0_3 ));
    CascadeMux I__5848 (
            .O(N__27682),
            .I(\VPP_VDDQ.count_2_1_3_cascade_ ));
    InMux I__5847 (
            .O(N__27679),
            .I(N__27675));
    InMux I__5846 (
            .O(N__27678),
            .I(N__27672));
    LocalMux I__5845 (
            .O(N__27675),
            .I(N__27667));
    LocalMux I__5844 (
            .O(N__27672),
            .I(N__27667));
    Span4Mux_h I__5843 (
            .O(N__27667),
            .I(N__27664));
    Odrv4 I__5842 (
            .O(N__27664),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    CascadeMux I__5841 (
            .O(N__27661),
            .I(\VPP_VDDQ.N_537_0_cascade_ ));
    CascadeMux I__5840 (
            .O(N__27658),
            .I(\VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0_cascade_ ));
    CascadeMux I__5839 (
            .O(N__27655),
            .I(N__27652));
    InMux I__5838 (
            .O(N__27652),
            .I(N__27649));
    LocalMux I__5837 (
            .O(N__27649),
            .I(\VPP_VDDQ.N_537_0 ));
    InMux I__5836 (
            .O(N__27646),
            .I(N__27642));
    InMux I__5835 (
            .O(N__27645),
            .I(N__27639));
    LocalMux I__5834 (
            .O(N__27642),
            .I(N__27636));
    LocalMux I__5833 (
            .O(N__27639),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    Odrv4 I__5832 (
            .O(N__27636),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    InMux I__5831 (
            .O(N__27631),
            .I(\RSMRST_PWRGD.un1_count_1_cry_9 ));
    InMux I__5830 (
            .O(N__27628),
            .I(N__27624));
    InMux I__5829 (
            .O(N__27627),
            .I(N__27621));
    LocalMux I__5828 (
            .O(N__27624),
            .I(N__27618));
    LocalMux I__5827 (
            .O(N__27621),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    Odrv4 I__5826 (
            .O(N__27618),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    InMux I__5825 (
            .O(N__27613),
            .I(\RSMRST_PWRGD.un1_count_1_cry_10 ));
    InMux I__5824 (
            .O(N__27610),
            .I(N__27606));
    InMux I__5823 (
            .O(N__27609),
            .I(N__27603));
    LocalMux I__5822 (
            .O(N__27606),
            .I(N__27600));
    LocalMux I__5821 (
            .O(N__27603),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    Odrv4 I__5820 (
            .O(N__27600),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    InMux I__5819 (
            .O(N__27595),
            .I(\RSMRST_PWRGD.un1_count_1_cry_11 ));
    InMux I__5818 (
            .O(N__27592),
            .I(N__27588));
    InMux I__5817 (
            .O(N__27591),
            .I(N__27585));
    LocalMux I__5816 (
            .O(N__27588),
            .I(N__27582));
    LocalMux I__5815 (
            .O(N__27585),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    Odrv4 I__5814 (
            .O(N__27582),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    InMux I__5813 (
            .O(N__27577),
            .I(\RSMRST_PWRGD.un1_count_1_cry_12 ));
    InMux I__5812 (
            .O(N__27574),
            .I(N__27513));
    InMux I__5811 (
            .O(N__27573),
            .I(N__27513));
    InMux I__5810 (
            .O(N__27572),
            .I(N__27513));
    InMux I__5809 (
            .O(N__27571),
            .I(N__27513));
    InMux I__5808 (
            .O(N__27570),
            .I(N__27504));
    InMux I__5807 (
            .O(N__27569),
            .I(N__27504));
    InMux I__5806 (
            .O(N__27568),
            .I(N__27504));
    InMux I__5805 (
            .O(N__27567),
            .I(N__27504));
    InMux I__5804 (
            .O(N__27566),
            .I(N__27495));
    InMux I__5803 (
            .O(N__27565),
            .I(N__27495));
    InMux I__5802 (
            .O(N__27564),
            .I(N__27495));
    InMux I__5801 (
            .O(N__27563),
            .I(N__27495));
    InMux I__5800 (
            .O(N__27562),
            .I(N__27486));
    InMux I__5799 (
            .O(N__27561),
            .I(N__27486));
    InMux I__5798 (
            .O(N__27560),
            .I(N__27486));
    InMux I__5797 (
            .O(N__27559),
            .I(N__27486));
    InMux I__5796 (
            .O(N__27558),
            .I(N__27479));
    InMux I__5795 (
            .O(N__27557),
            .I(N__27479));
    InMux I__5794 (
            .O(N__27556),
            .I(N__27479));
    InMux I__5793 (
            .O(N__27555),
            .I(N__27470));
    InMux I__5792 (
            .O(N__27554),
            .I(N__27470));
    InMux I__5791 (
            .O(N__27553),
            .I(N__27470));
    InMux I__5790 (
            .O(N__27552),
            .I(N__27470));
    InMux I__5789 (
            .O(N__27551),
            .I(N__27461));
    InMux I__5788 (
            .O(N__27550),
            .I(N__27461));
    InMux I__5787 (
            .O(N__27549),
            .I(N__27461));
    InMux I__5786 (
            .O(N__27548),
            .I(N__27461));
    InMux I__5785 (
            .O(N__27547),
            .I(N__27454));
    InMux I__5784 (
            .O(N__27546),
            .I(N__27454));
    InMux I__5783 (
            .O(N__27545),
            .I(N__27454));
    InMux I__5782 (
            .O(N__27544),
            .I(N__27445));
    InMux I__5781 (
            .O(N__27543),
            .I(N__27445));
    InMux I__5780 (
            .O(N__27542),
            .I(N__27445));
    InMux I__5779 (
            .O(N__27541),
            .I(N__27445));
    InMux I__5778 (
            .O(N__27540),
            .I(N__27436));
    InMux I__5777 (
            .O(N__27539),
            .I(N__27436));
    InMux I__5776 (
            .O(N__27538),
            .I(N__27436));
    InMux I__5775 (
            .O(N__27537),
            .I(N__27436));
    InMux I__5774 (
            .O(N__27536),
            .I(N__27427));
    InMux I__5773 (
            .O(N__27535),
            .I(N__27427));
    InMux I__5772 (
            .O(N__27534),
            .I(N__27427));
    InMux I__5771 (
            .O(N__27533),
            .I(N__27427));
    InMux I__5770 (
            .O(N__27532),
            .I(N__27420));
    InMux I__5769 (
            .O(N__27531),
            .I(N__27420));
    InMux I__5768 (
            .O(N__27530),
            .I(N__27420));
    InMux I__5767 (
            .O(N__27529),
            .I(N__27415));
    InMux I__5766 (
            .O(N__27528),
            .I(N__27415));
    InMux I__5765 (
            .O(N__27527),
            .I(N__27410));
    InMux I__5764 (
            .O(N__27526),
            .I(N__27410));
    InMux I__5763 (
            .O(N__27525),
            .I(N__27407));
    InMux I__5762 (
            .O(N__27524),
            .I(N__27402));
    InMux I__5761 (
            .O(N__27523),
            .I(N__27402));
    InMux I__5760 (
            .O(N__27522),
            .I(N__27399));
    LocalMux I__5759 (
            .O(N__27513),
            .I(N__27395));
    LocalMux I__5758 (
            .O(N__27504),
            .I(N__27391));
    LocalMux I__5757 (
            .O(N__27495),
            .I(N__27382));
    LocalMux I__5756 (
            .O(N__27486),
            .I(N__27377));
    LocalMux I__5755 (
            .O(N__27479),
            .I(N__27374));
    LocalMux I__5754 (
            .O(N__27470),
            .I(N__27371));
    LocalMux I__5753 (
            .O(N__27461),
            .I(N__27368));
    LocalMux I__5752 (
            .O(N__27454),
            .I(N__27365));
    LocalMux I__5751 (
            .O(N__27445),
            .I(N__27362));
    LocalMux I__5750 (
            .O(N__27436),
            .I(N__27359));
    LocalMux I__5749 (
            .O(N__27427),
            .I(N__27356));
    LocalMux I__5748 (
            .O(N__27420),
            .I(N__27353));
    LocalMux I__5747 (
            .O(N__27415),
            .I(N__27350));
    LocalMux I__5746 (
            .O(N__27410),
            .I(N__27347));
    LocalMux I__5745 (
            .O(N__27407),
            .I(N__27344));
    LocalMux I__5744 (
            .O(N__27402),
            .I(N__27341));
    LocalMux I__5743 (
            .O(N__27399),
            .I(N__27338));
    CEMux I__5742 (
            .O(N__27398),
            .I(N__27283));
    Glb2LocalMux I__5741 (
            .O(N__27395),
            .I(N__27283));
    CEMux I__5740 (
            .O(N__27394),
            .I(N__27283));
    Glb2LocalMux I__5739 (
            .O(N__27391),
            .I(N__27283));
    CEMux I__5738 (
            .O(N__27390),
            .I(N__27283));
    CEMux I__5737 (
            .O(N__27389),
            .I(N__27283));
    CEMux I__5736 (
            .O(N__27388),
            .I(N__27283));
    CEMux I__5735 (
            .O(N__27387),
            .I(N__27283));
    CEMux I__5734 (
            .O(N__27386),
            .I(N__27283));
    CEMux I__5733 (
            .O(N__27385),
            .I(N__27283));
    Glb2LocalMux I__5732 (
            .O(N__27382),
            .I(N__27283));
    CEMux I__5731 (
            .O(N__27381),
            .I(N__27283));
    CEMux I__5730 (
            .O(N__27380),
            .I(N__27283));
    Glb2LocalMux I__5729 (
            .O(N__27377),
            .I(N__27283));
    Glb2LocalMux I__5728 (
            .O(N__27374),
            .I(N__27283));
    Glb2LocalMux I__5727 (
            .O(N__27371),
            .I(N__27283));
    Glb2LocalMux I__5726 (
            .O(N__27368),
            .I(N__27283));
    Glb2LocalMux I__5725 (
            .O(N__27365),
            .I(N__27283));
    Glb2LocalMux I__5724 (
            .O(N__27362),
            .I(N__27283));
    Glb2LocalMux I__5723 (
            .O(N__27359),
            .I(N__27283));
    Glb2LocalMux I__5722 (
            .O(N__27356),
            .I(N__27283));
    Glb2LocalMux I__5721 (
            .O(N__27353),
            .I(N__27283));
    Glb2LocalMux I__5720 (
            .O(N__27350),
            .I(N__27283));
    Glb2LocalMux I__5719 (
            .O(N__27347),
            .I(N__27283));
    Glb2LocalMux I__5718 (
            .O(N__27344),
            .I(N__27283));
    Glb2LocalMux I__5717 (
            .O(N__27341),
            .I(N__27283));
    Glb2LocalMux I__5716 (
            .O(N__27338),
            .I(N__27283));
    GlobalMux I__5715 (
            .O(N__27283),
            .I(N__27280));
    gio2CtrlBuf I__5714 (
            .O(N__27280),
            .I(N_42_g));
    InMux I__5713 (
            .O(N__27277),
            .I(N__27273));
    InMux I__5712 (
            .O(N__27276),
            .I(N__27270));
    LocalMux I__5711 (
            .O(N__27273),
            .I(N__27267));
    LocalMux I__5710 (
            .O(N__27270),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    Odrv4 I__5709 (
            .O(N__27267),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    InMux I__5708 (
            .O(N__27262),
            .I(\RSMRST_PWRGD.un1_count_1_cry_13 ));
    InMux I__5707 (
            .O(N__27259),
            .I(N__27256));
    LocalMux I__5706 (
            .O(N__27256),
            .I(N__27251));
    IoInMux I__5705 (
            .O(N__27255),
            .I(N__27248));
    InMux I__5704 (
            .O(N__27254),
            .I(N__27245));
    Span4Mux_s3_h I__5703 (
            .O(N__27251),
            .I(N__27241));
    LocalMux I__5702 (
            .O(N__27248),
            .I(N__27238));
    LocalMux I__5701 (
            .O(N__27245),
            .I(N__27231));
    InMux I__5700 (
            .O(N__27244),
            .I(N__27228));
    Span4Mux_v I__5699 (
            .O(N__27241),
            .I(N__27223));
    Span4Mux_s3_h I__5698 (
            .O(N__27238),
            .I(N__27223));
    InMux I__5697 (
            .O(N__27237),
            .I(N__27220));
    InMux I__5696 (
            .O(N__27236),
            .I(N__27217));
    InMux I__5695 (
            .O(N__27235),
            .I(N__27214));
    InMux I__5694 (
            .O(N__27234),
            .I(N__27211));
    Span12Mux_s3_v I__5693 (
            .O(N__27231),
            .I(N__27208));
    LocalMux I__5692 (
            .O(N__27228),
            .I(N__27205));
    Span4Mux_v I__5691 (
            .O(N__27223),
            .I(N__27200));
    LocalMux I__5690 (
            .O(N__27220),
            .I(N__27200));
    LocalMux I__5689 (
            .O(N__27217),
            .I(N__27193));
    LocalMux I__5688 (
            .O(N__27214),
            .I(N__27193));
    LocalMux I__5687 (
            .O(N__27211),
            .I(N__27193));
    Span12Mux_v I__5686 (
            .O(N__27208),
            .I(N__27190));
    Span12Mux_s8_v I__5685 (
            .O(N__27205),
            .I(N__27187));
    Span4Mux_v I__5684 (
            .O(N__27200),
            .I(N__27184));
    Span4Mux_v I__5683 (
            .O(N__27193),
            .I(N__27181));
    Odrv12 I__5682 (
            .O(N__27190),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__5681 (
            .O(N__27187),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5680 (
            .O(N__27184),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5679 (
            .O(N__27181),
            .I(CONSTANT_ONE_NET));
    InMux I__5678 (
            .O(N__27172),
            .I(bfn_11_14_0_));
    CascadeMux I__5677 (
            .O(N__27169),
            .I(N__27166));
    InMux I__5676 (
            .O(N__27166),
            .I(N__27162));
    InMux I__5675 (
            .O(N__27165),
            .I(N__27159));
    LocalMux I__5674 (
            .O(N__27162),
            .I(N__27156));
    LocalMux I__5673 (
            .O(N__27159),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    Odrv12 I__5672 (
            .O(N__27156),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    CEMux I__5671 (
            .O(N__27151),
            .I(N__27148));
    LocalMux I__5670 (
            .O(N__27148),
            .I(N__27145));
    Span4Mux_h I__5669 (
            .O(N__27145),
            .I(N__27142));
    Odrv4 I__5668 (
            .O(N__27142),
            .I(\RSMRST_PWRGD.N_42_2 ));
    SRMux I__5667 (
            .O(N__27139),
            .I(N__27134));
    SRMux I__5666 (
            .O(N__27138),
            .I(N__27131));
    SRMux I__5665 (
            .O(N__27137),
            .I(N__27128));
    LocalMux I__5664 (
            .O(N__27134),
            .I(N__27124));
    LocalMux I__5663 (
            .O(N__27131),
            .I(N__27119));
    LocalMux I__5662 (
            .O(N__27128),
            .I(N__27119));
    InMux I__5661 (
            .O(N__27127),
            .I(N__27116));
    Span4Mux_v I__5660 (
            .O(N__27124),
            .I(N__27111));
    Span4Mux_v I__5659 (
            .O(N__27119),
            .I(N__27111));
    LocalMux I__5658 (
            .O(N__27116),
            .I(N__27108));
    Odrv4 I__5657 (
            .O(N__27111),
            .I(G_12));
    Odrv4 I__5656 (
            .O(N__27108),
            .I(G_12));
    InMux I__5655 (
            .O(N__27103),
            .I(N__27099));
    InMux I__5654 (
            .O(N__27102),
            .I(N__27096));
    LocalMux I__5653 (
            .O(N__27099),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    LocalMux I__5652 (
            .O(N__27096),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    InMux I__5651 (
            .O(N__27091),
            .I(\RSMRST_PWRGD.un1_count_1_cry_0 ));
    InMux I__5650 (
            .O(N__27088),
            .I(N__27084));
    InMux I__5649 (
            .O(N__27087),
            .I(N__27081));
    LocalMux I__5648 (
            .O(N__27084),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    LocalMux I__5647 (
            .O(N__27081),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    InMux I__5646 (
            .O(N__27076),
            .I(\RSMRST_PWRGD.un1_count_1_cry_1 ));
    CascadeMux I__5645 (
            .O(N__27073),
            .I(N__27070));
    InMux I__5644 (
            .O(N__27070),
            .I(N__27066));
    InMux I__5643 (
            .O(N__27069),
            .I(N__27063));
    LocalMux I__5642 (
            .O(N__27066),
            .I(N__27060));
    LocalMux I__5641 (
            .O(N__27063),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    Odrv4 I__5640 (
            .O(N__27060),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    InMux I__5639 (
            .O(N__27055),
            .I(\RSMRST_PWRGD.un1_count_1_cry_2 ));
    InMux I__5638 (
            .O(N__27052),
            .I(N__27048));
    InMux I__5637 (
            .O(N__27051),
            .I(N__27045));
    LocalMux I__5636 (
            .O(N__27048),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    LocalMux I__5635 (
            .O(N__27045),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    InMux I__5634 (
            .O(N__27040),
            .I(\RSMRST_PWRGD.un1_count_1_cry_3 ));
    InMux I__5633 (
            .O(N__27037),
            .I(N__27033));
    InMux I__5632 (
            .O(N__27036),
            .I(N__27030));
    LocalMux I__5631 (
            .O(N__27033),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    LocalMux I__5630 (
            .O(N__27030),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    InMux I__5629 (
            .O(N__27025),
            .I(\RSMRST_PWRGD.un1_count_1_cry_4 ));
    InMux I__5628 (
            .O(N__27022),
            .I(N__27018));
    InMux I__5627 (
            .O(N__27021),
            .I(N__27015));
    LocalMux I__5626 (
            .O(N__27018),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    LocalMux I__5625 (
            .O(N__27015),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    InMux I__5624 (
            .O(N__27010),
            .I(\RSMRST_PWRGD.un1_count_1_cry_5 ));
    InMux I__5623 (
            .O(N__27007),
            .I(N__27003));
    InMux I__5622 (
            .O(N__27006),
            .I(N__27000));
    LocalMux I__5621 (
            .O(N__27003),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    LocalMux I__5620 (
            .O(N__27000),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    InMux I__5619 (
            .O(N__26995),
            .I(\RSMRST_PWRGD.un1_count_1_cry_6 ));
    InMux I__5618 (
            .O(N__26992),
            .I(N__26988));
    InMux I__5617 (
            .O(N__26991),
            .I(N__26985));
    LocalMux I__5616 (
            .O(N__26988),
            .I(N__26982));
    LocalMux I__5615 (
            .O(N__26985),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    Odrv4 I__5614 (
            .O(N__26982),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    InMux I__5613 (
            .O(N__26977),
            .I(bfn_11_13_0_));
    CascadeMux I__5612 (
            .O(N__26974),
            .I(N__26971));
    InMux I__5611 (
            .O(N__26971),
            .I(N__26967));
    InMux I__5610 (
            .O(N__26970),
            .I(N__26964));
    LocalMux I__5609 (
            .O(N__26967),
            .I(N__26961));
    LocalMux I__5608 (
            .O(N__26964),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    Odrv4 I__5607 (
            .O(N__26961),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    InMux I__5606 (
            .O(N__26956),
            .I(\RSMRST_PWRGD.un1_count_1_cry_8 ));
    InMux I__5605 (
            .O(N__26953),
            .I(N__26950));
    LocalMux I__5604 (
            .O(N__26950),
            .I(N__26947));
    Span4Mux_h I__5603 (
            .O(N__26947),
            .I(N__26944));
    Odrv4 I__5602 (
            .O(N__26944),
            .I(\POWERLED.m69_0_o2_2 ));
    CascadeMux I__5601 (
            .O(N__26941),
            .I(N__26936));
    InMux I__5600 (
            .O(N__26940),
            .I(N__26933));
    InMux I__5599 (
            .O(N__26939),
            .I(N__26930));
    InMux I__5598 (
            .O(N__26936),
            .I(N__26927));
    LocalMux I__5597 (
            .O(N__26933),
            .I(N__26917));
    LocalMux I__5596 (
            .O(N__26930),
            .I(N__26917));
    LocalMux I__5595 (
            .O(N__26927),
            .I(N__26917));
    InMux I__5594 (
            .O(N__26926),
            .I(N__26914));
    InMux I__5593 (
            .O(N__26925),
            .I(N__26909));
    InMux I__5592 (
            .O(N__26924),
            .I(N__26909));
    Span4Mux_v I__5591 (
            .O(N__26917),
            .I(N__26904));
    LocalMux I__5590 (
            .O(N__26914),
            .I(N__26904));
    LocalMux I__5589 (
            .O(N__26909),
            .I(RSMRSTn_rep1));
    Odrv4 I__5588 (
            .O(N__26904),
            .I(RSMRSTn_rep1));
    InMux I__5587 (
            .O(N__26899),
            .I(N__26896));
    LocalMux I__5586 (
            .O(N__26896),
            .I(N__26893));
    Span4Mux_h I__5585 (
            .O(N__26893),
            .I(N__26890));
    Odrv4 I__5584 (
            .O(N__26890),
            .I(N_110_0));
    CascadeMux I__5583 (
            .O(N__26887),
            .I(\RSMRST_PWRGD.un4_count_9_cascade_ ));
    InMux I__5582 (
            .O(N__26884),
            .I(N__26878));
    InMux I__5581 (
            .O(N__26883),
            .I(N__26878));
    LocalMux I__5580 (
            .O(N__26878),
            .I(N__26875));
    Odrv4 I__5579 (
            .O(N__26875),
            .I(\RSMRST_PWRGD.N_1_i ));
    InMux I__5578 (
            .O(N__26872),
            .I(N__26869));
    LocalMux I__5577 (
            .O(N__26869),
            .I(\RSMRST_PWRGD.un4_count_8 ));
    InMux I__5576 (
            .O(N__26866),
            .I(N__26863));
    LocalMux I__5575 (
            .O(N__26863),
            .I(\RSMRST_PWRGD.un4_count_10 ));
    InMux I__5574 (
            .O(N__26860),
            .I(N__26857));
    LocalMux I__5573 (
            .O(N__26857),
            .I(\RSMRST_PWRGD.un4_count_11 ));
    CascadeMux I__5572 (
            .O(N__26854),
            .I(N__26850));
    InMux I__5571 (
            .O(N__26853),
            .I(N__26847));
    InMux I__5570 (
            .O(N__26850),
            .I(N__26844));
    LocalMux I__5569 (
            .O(N__26847),
            .I(N__26839));
    LocalMux I__5568 (
            .O(N__26844),
            .I(N__26839));
    Odrv4 I__5567 (
            .O(N__26839),
            .I(\RSMRST_PWRGD.N_445_i ));
    CascadeMux I__5566 (
            .O(N__26836),
            .I(N__26833));
    InMux I__5565 (
            .O(N__26833),
            .I(N__26829));
    InMux I__5564 (
            .O(N__26832),
            .I(N__26826));
    LocalMux I__5563 (
            .O(N__26829),
            .I(N__26823));
    LocalMux I__5562 (
            .O(N__26826),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    Odrv4 I__5561 (
            .O(N__26823),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    InMux I__5560 (
            .O(N__26818),
            .I(N__26815));
    LocalMux I__5559 (
            .O(N__26815),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_6 ));
    CascadeMux I__5558 (
            .O(N__26812),
            .I(\POWERLED.un1_dutycycle_172_m2s4_1_cascade_ ));
    InMux I__5557 (
            .O(N__26809),
            .I(N__26803));
    InMux I__5556 (
            .O(N__26808),
            .I(N__26803));
    LocalMux I__5555 (
            .O(N__26803),
            .I(N__26799));
    InMux I__5554 (
            .O(N__26802),
            .I(N__26796));
    Span4Mux_s2_h I__5553 (
            .O(N__26799),
            .I(N__26793));
    LocalMux I__5552 (
            .O(N__26796),
            .I(N__26790));
    Span4Mux_h I__5551 (
            .O(N__26793),
            .I(N__26787));
    Span4Mux_v I__5550 (
            .O(N__26790),
            .I(N__26784));
    Odrv4 I__5549 (
            .O(N__26787),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_1 ));
    Odrv4 I__5548 (
            .O(N__26784),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_1 ));
    InMux I__5547 (
            .O(N__26779),
            .I(N__26776));
    LocalMux I__5546 (
            .O(N__26776),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_3 ));
    InMux I__5545 (
            .O(N__26773),
            .I(N__26770));
    LocalMux I__5544 (
            .O(N__26770),
            .I(\POWERLED.N_414 ));
    CascadeMux I__5543 (
            .O(N__26767),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_3_cascade_ ));
    InMux I__5542 (
            .O(N__26764),
            .I(N__26761));
    LocalMux I__5541 (
            .O(N__26761),
            .I(N__26758));
    Odrv12 I__5540 (
            .O(N__26758),
            .I(\POWERLED.g0_i_1_1_0 ));
    InMux I__5539 (
            .O(N__26755),
            .I(N__26751));
    CascadeMux I__5538 (
            .O(N__26754),
            .I(N__26748));
    LocalMux I__5537 (
            .O(N__26751),
            .I(N__26745));
    InMux I__5536 (
            .O(N__26748),
            .I(N__26742));
    Span4Mux_s3_h I__5535 (
            .O(N__26745),
            .I(N__26739));
    LocalMux I__5534 (
            .O(N__26742),
            .I(N__26736));
    Odrv4 I__5533 (
            .O(N__26739),
            .I(\POWERLED.func_state_RNI56A8Z0Z_0 ));
    Odrv4 I__5532 (
            .O(N__26736),
            .I(\POWERLED.func_state_RNI56A8Z0Z_0 ));
    CascadeMux I__5531 (
            .O(N__26731),
            .I(N__26727));
    CascadeMux I__5530 (
            .O(N__26730),
            .I(N__26723));
    InMux I__5529 (
            .O(N__26727),
            .I(N__26720));
    InMux I__5528 (
            .O(N__26726),
            .I(N__26717));
    InMux I__5527 (
            .O(N__26723),
            .I(N__26714));
    LocalMux I__5526 (
            .O(N__26720),
            .I(N__26709));
    LocalMux I__5525 (
            .O(N__26717),
            .I(N__26709));
    LocalMux I__5524 (
            .O(N__26714),
            .I(N__26706));
    Span4Mux_s2_h I__5523 (
            .O(N__26709),
            .I(N__26703));
    Odrv12 I__5522 (
            .O(N__26706),
            .I(\POWERLED.N_239 ));
    Odrv4 I__5521 (
            .O(N__26703),
            .I(\POWERLED.N_239 ));
    InMux I__5520 (
            .O(N__26698),
            .I(N__26695));
    LocalMux I__5519 (
            .O(N__26695),
            .I(N__26692));
    Span4Mux_h I__5518 (
            .O(N__26692),
            .I(N__26689));
    Odrv4 I__5517 (
            .O(N__26689),
            .I(\POWERLED.N_462 ));
    InMux I__5516 (
            .O(N__26686),
            .I(N__26683));
    LocalMux I__5515 (
            .O(N__26683),
            .I(N__26680));
    Span4Mux_v I__5514 (
            .O(N__26680),
            .I(N__26676));
    InMux I__5513 (
            .O(N__26679),
            .I(N__26673));
    Odrv4 I__5512 (
            .O(N__26676),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_6 ));
    LocalMux I__5511 (
            .O(N__26673),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_6 ));
    CascadeMux I__5510 (
            .O(N__26668),
            .I(\POWERLED.un1_clk_100khz_52_and_i_0_m3_1_rn_1_cascade_ ));
    InMux I__5509 (
            .O(N__26665),
            .I(N__26662));
    LocalMux I__5508 (
            .O(N__26662),
            .I(N__26659));
    Span4Mux_h I__5507 (
            .O(N__26659),
            .I(N__26656));
    Odrv4 I__5506 (
            .O(N__26656),
            .I(POWERLED_un1_clk_100khz_52_and_i_0_m3_1));
    SRMux I__5505 (
            .O(N__26653),
            .I(N__26645));
    SRMux I__5504 (
            .O(N__26652),
            .I(N__26642));
    SRMux I__5503 (
            .O(N__26651),
            .I(N__26638));
    SRMux I__5502 (
            .O(N__26650),
            .I(N__26635));
    SRMux I__5501 (
            .O(N__26649),
            .I(N__26627));
    SRMux I__5500 (
            .O(N__26648),
            .I(N__26624));
    LocalMux I__5499 (
            .O(N__26645),
            .I(N__26621));
    LocalMux I__5498 (
            .O(N__26642),
            .I(N__26618));
    SRMux I__5497 (
            .O(N__26641),
            .I(N__26615));
    LocalMux I__5496 (
            .O(N__26638),
            .I(N__26612));
    LocalMux I__5495 (
            .O(N__26635),
            .I(N__26609));
    SRMux I__5494 (
            .O(N__26634),
            .I(N__26606));
    SRMux I__5493 (
            .O(N__26633),
            .I(N__26603));
    SRMux I__5492 (
            .O(N__26632),
            .I(N__26599));
    SRMux I__5491 (
            .O(N__26631),
            .I(N__26596));
    SRMux I__5490 (
            .O(N__26630),
            .I(N__26593));
    LocalMux I__5489 (
            .O(N__26627),
            .I(N__26590));
    LocalMux I__5488 (
            .O(N__26624),
            .I(N__26581));
    Span4Mux_v I__5487 (
            .O(N__26621),
            .I(N__26581));
    Span4Mux_h I__5486 (
            .O(N__26618),
            .I(N__26581));
    LocalMux I__5485 (
            .O(N__26615),
            .I(N__26581));
    Span4Mux_v I__5484 (
            .O(N__26612),
            .I(N__26578));
    Span4Mux_h I__5483 (
            .O(N__26609),
            .I(N__26573));
    LocalMux I__5482 (
            .O(N__26606),
            .I(N__26573));
    LocalMux I__5481 (
            .O(N__26603),
            .I(N__26570));
    SRMux I__5480 (
            .O(N__26602),
            .I(N__26567));
    LocalMux I__5479 (
            .O(N__26599),
            .I(N__26564));
    LocalMux I__5478 (
            .O(N__26596),
            .I(N__26561));
    LocalMux I__5477 (
            .O(N__26593),
            .I(N__26556));
    Span4Mux_v I__5476 (
            .O(N__26590),
            .I(N__26556));
    Span4Mux_v I__5475 (
            .O(N__26581),
            .I(N__26553));
    Span4Mux_h I__5474 (
            .O(N__26578),
            .I(N__26548));
    Span4Mux_v I__5473 (
            .O(N__26573),
            .I(N__26548));
    Span4Mux_v I__5472 (
            .O(N__26570),
            .I(N__26541));
    LocalMux I__5471 (
            .O(N__26567),
            .I(N__26541));
    Span4Mux_s2_v I__5470 (
            .O(N__26564),
            .I(N__26541));
    Span4Mux_v I__5469 (
            .O(N__26561),
            .I(N__26538));
    Span4Mux_h I__5468 (
            .O(N__26556),
            .I(N__26535));
    Span4Mux_v I__5467 (
            .O(N__26553),
            .I(N__26532));
    Span4Mux_h I__5466 (
            .O(N__26548),
            .I(N__26527));
    Span4Mux_v I__5465 (
            .O(N__26541),
            .I(N__26527));
    Odrv4 I__5464 (
            .O(N__26538),
            .I(\POWERLED.dutycycle_eena_5_0_s_tz_isoZ0 ));
    Odrv4 I__5463 (
            .O(N__26535),
            .I(\POWERLED.dutycycle_eena_5_0_s_tz_isoZ0 ));
    Odrv4 I__5462 (
            .O(N__26532),
            .I(\POWERLED.dutycycle_eena_5_0_s_tz_isoZ0 ));
    Odrv4 I__5461 (
            .O(N__26527),
            .I(\POWERLED.dutycycle_eena_5_0_s_tz_isoZ0 ));
    InMux I__5460 (
            .O(N__26518),
            .I(N__26515));
    LocalMux I__5459 (
            .O(N__26515),
            .I(\POWERLED.dutycycle_eena_4 ));
    InMux I__5458 (
            .O(N__26512),
            .I(N__26506));
    InMux I__5457 (
            .O(N__26511),
            .I(N__26506));
    LocalMux I__5456 (
            .O(N__26506),
            .I(\POWERLED.dutycycleZ1Z_10 ));
    CascadeMux I__5455 (
            .O(N__26503),
            .I(\POWERLED.dutycycle_eena_4_cascade_ ));
    InMux I__5454 (
            .O(N__26500),
            .I(N__26494));
    InMux I__5453 (
            .O(N__26499),
            .I(N__26494));
    LocalMux I__5452 (
            .O(N__26494),
            .I(N__26491));
    Odrv4 I__5451 (
            .O(N__26491),
            .I(\POWERLED.un1_dutycycle_94_cry_9_c_RNI4D3UZ0 ));
    CascadeMux I__5450 (
            .O(N__26488),
            .I(\POWERLED.dutycycleZ0Z_5_cascade_ ));
    InMux I__5449 (
            .O(N__26485),
            .I(N__26479));
    InMux I__5448 (
            .O(N__26484),
            .I(N__26479));
    LocalMux I__5447 (
            .O(N__26479),
            .I(\POWERLED.dutycycleZ1Z_12 ));
    CascadeMux I__5446 (
            .O(N__26476),
            .I(N__26473));
    InMux I__5445 (
            .O(N__26473),
            .I(N__26470));
    LocalMux I__5444 (
            .O(N__26470),
            .I(\POWERLED.dutycycle_eena_9 ));
    InMux I__5443 (
            .O(N__26467),
            .I(N__26463));
    InMux I__5442 (
            .O(N__26466),
            .I(N__26460));
    LocalMux I__5441 (
            .O(N__26463),
            .I(N__26457));
    LocalMux I__5440 (
            .O(N__26460),
            .I(N__26454));
    Odrv12 I__5439 (
            .O(N__26457),
            .I(\POWERLED.un1_dutycycle_94_cry_11_c_RNID2MBZ0Z1 ));
    Odrv4 I__5438 (
            .O(N__26454),
            .I(\POWERLED.un1_dutycycle_94_cry_11_c_RNID2MBZ0Z1 ));
    InMux I__5437 (
            .O(N__26449),
            .I(N__26446));
    LocalMux I__5436 (
            .O(N__26446),
            .I(\POWERLED.un1_dutycycle_53_7_3_0_1 ));
    CascadeMux I__5435 (
            .O(N__26443),
            .I(\POWERLED.dutycycleZ0Z_10_cascade_ ));
    InMux I__5434 (
            .O(N__26440),
            .I(N__26437));
    LocalMux I__5433 (
            .O(N__26437),
            .I(N__26434));
    Span4Mux_s1_h I__5432 (
            .O(N__26434),
            .I(N__26431));
    Odrv4 I__5431 (
            .O(N__26431),
            .I(\POWERLED.un1_dutycycle_53_7_3 ));
    CascadeMux I__5430 (
            .O(N__26428),
            .I(N__26422));
    InMux I__5429 (
            .O(N__26427),
            .I(N__26416));
    InMux I__5428 (
            .O(N__26426),
            .I(N__26411));
    InMux I__5427 (
            .O(N__26425),
            .I(N__26406));
    InMux I__5426 (
            .O(N__26422),
            .I(N__26406));
    InMux I__5425 (
            .O(N__26421),
            .I(N__26403));
    CascadeMux I__5424 (
            .O(N__26420),
            .I(N__26400));
    CascadeMux I__5423 (
            .O(N__26419),
            .I(N__26397));
    LocalMux I__5422 (
            .O(N__26416),
            .I(N__26393));
    InMux I__5421 (
            .O(N__26415),
            .I(N__26390));
    InMux I__5420 (
            .O(N__26414),
            .I(N__26387));
    LocalMux I__5419 (
            .O(N__26411),
            .I(N__26382));
    LocalMux I__5418 (
            .O(N__26406),
            .I(N__26382));
    LocalMux I__5417 (
            .O(N__26403),
            .I(N__26379));
    InMux I__5416 (
            .O(N__26400),
            .I(N__26376));
    InMux I__5415 (
            .O(N__26397),
            .I(N__26373));
    InMux I__5414 (
            .O(N__26396),
            .I(N__26370));
    Span4Mux_s3_h I__5413 (
            .O(N__26393),
            .I(N__26363));
    LocalMux I__5412 (
            .O(N__26390),
            .I(N__26363));
    LocalMux I__5411 (
            .O(N__26387),
            .I(N__26363));
    Sp12to4 I__5410 (
            .O(N__26382),
            .I(N__26360));
    Span4Mux_h I__5409 (
            .O(N__26379),
            .I(N__26355));
    LocalMux I__5408 (
            .O(N__26376),
            .I(N__26355));
    LocalMux I__5407 (
            .O(N__26373),
            .I(dutycycle_RNINBHJ5_0_2));
    LocalMux I__5406 (
            .O(N__26370),
            .I(dutycycle_RNINBHJ5_0_2));
    Odrv4 I__5405 (
            .O(N__26363),
            .I(dutycycle_RNINBHJ5_0_2));
    Odrv12 I__5404 (
            .O(N__26360),
            .I(dutycycle_RNINBHJ5_0_2));
    Odrv4 I__5403 (
            .O(N__26355),
            .I(dutycycle_RNINBHJ5_0_2));
    InMux I__5402 (
            .O(N__26344),
            .I(N__26340));
    InMux I__5401 (
            .O(N__26343),
            .I(N__26337));
    LocalMux I__5400 (
            .O(N__26340),
            .I(N__26334));
    LocalMux I__5399 (
            .O(N__26337),
            .I(N__26331));
    Span4Mux_v I__5398 (
            .O(N__26334),
            .I(N__26328));
    Span4Mux_v I__5397 (
            .O(N__26331),
            .I(N__26325));
    Span4Mux_h I__5396 (
            .O(N__26328),
            .I(N__26322));
    Odrv4 I__5395 (
            .O(N__26325),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_1 ));
    Odrv4 I__5394 (
            .O(N__26322),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_1 ));
    CascadeMux I__5393 (
            .O(N__26317),
            .I(\POWERLED.un1_dutycycle_172_m2s4_1_1_cascade_ ));
    CascadeMux I__5392 (
            .O(N__26314),
            .I(\POWERLED.un1_dutycycle_53_13_a1_1_cascade_ ));
    InMux I__5391 (
            .O(N__26311),
            .I(N__26307));
    InMux I__5390 (
            .O(N__26310),
            .I(N__26304));
    LocalMux I__5389 (
            .O(N__26307),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__5388 (
            .O(N__26304),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    CascadeMux I__5387 (
            .O(N__26299),
            .I(N__26295));
    InMux I__5386 (
            .O(N__26298),
            .I(N__26292));
    InMux I__5385 (
            .O(N__26295),
            .I(N__26289));
    LocalMux I__5384 (
            .O(N__26292),
            .I(N__26284));
    LocalMux I__5383 (
            .O(N__26289),
            .I(N__26284));
    Span4Mux_s2_h I__5382 (
            .O(N__26284),
            .I(N__26281));
    Odrv4 I__5381 (
            .O(N__26281),
            .I(\POWERLED.un1_dutycycle_94_cry_10_c_RNIC0LBZ0Z1 ));
    InMux I__5380 (
            .O(N__26278),
            .I(N__26272));
    InMux I__5379 (
            .O(N__26277),
            .I(N__26272));
    LocalMux I__5378 (
            .O(N__26272),
            .I(\POWERLED.dutycycle_eena_7 ));
    CascadeMux I__5377 (
            .O(N__26269),
            .I(\POWERLED.dutycycleZ0Z_7_cascade_ ));
    InMux I__5376 (
            .O(N__26266),
            .I(N__26263));
    LocalMux I__5375 (
            .O(N__26263),
            .I(\POWERLED.un1_dutycycle_53_46_a3_1 ));
    CascadeMux I__5374 (
            .O(N__26260),
            .I(\POWERLED.un1_dutycycle_53_46_a3_1_cascade_ ));
    InMux I__5373 (
            .O(N__26257),
            .I(N__26254));
    LocalMux I__5372 (
            .O(N__26254),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_7 ));
    InMux I__5371 (
            .O(N__26251),
            .I(N__26248));
    LocalMux I__5370 (
            .O(N__26248),
            .I(\POWERLED.un1_dutycycle_53_46_a3_d ));
    CascadeMux I__5369 (
            .O(N__26245),
            .I(\POWERLED.dutycycle_eena_9_cascade_ ));
    InMux I__5368 (
            .O(N__26242),
            .I(N__26236));
    InMux I__5367 (
            .O(N__26241),
            .I(N__26236));
    LocalMux I__5366 (
            .O(N__26236),
            .I(\POWERLED.dutycycleZ1Z_8 ));
    CascadeMux I__5365 (
            .O(N__26233),
            .I(N__26229));
    InMux I__5364 (
            .O(N__26232),
            .I(N__26224));
    InMux I__5363 (
            .O(N__26229),
            .I(N__26224));
    LocalMux I__5362 (
            .O(N__26224),
            .I(N__26221));
    Span4Mux_s2_h I__5361 (
            .O(N__26221),
            .I(N__26218));
    Odrv4 I__5360 (
            .O(N__26218),
            .I(\POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ));
    CascadeMux I__5359 (
            .O(N__26215),
            .I(\POWERLED.dutycycleZ0Z_1_cascade_ ));
    CascadeMux I__5358 (
            .O(N__26212),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_11_cascade_ ));
    InMux I__5357 (
            .O(N__26209),
            .I(N__26203));
    InMux I__5356 (
            .O(N__26208),
            .I(N__26203));
    LocalMux I__5355 (
            .O(N__26203),
            .I(N__26200));
    Odrv4 I__5354 (
            .O(N__26200),
            .I(\POWERLED.un1_dutycycle_53_57_a0_1_1 ));
    CascadeMux I__5353 (
            .O(N__26197),
            .I(\POWERLED.un1_dutycycle_53_2_0_cascade_ ));
    InMux I__5352 (
            .O(N__26194),
            .I(N__26191));
    LocalMux I__5351 (
            .O(N__26191),
            .I(\POWERLED.dutycycle_RNI_10Z0Z_10 ));
    InMux I__5350 (
            .O(N__26188),
            .I(N__26185));
    LocalMux I__5349 (
            .O(N__26185),
            .I(N__26182));
    Span4Mux_h I__5348 (
            .O(N__26182),
            .I(N__26179));
    Odrv4 I__5347 (
            .O(N__26179),
            .I(\POWERLED.dutycycle_RNI_11Z0Z_10 ));
    InMux I__5346 (
            .O(N__26176),
            .I(N__26173));
    LocalMux I__5345 (
            .O(N__26173),
            .I(N__26169));
    InMux I__5344 (
            .O(N__26172),
            .I(N__26166));
    Span12Mux_s7_v I__5343 (
            .O(N__26169),
            .I(N__26163));
    LocalMux I__5342 (
            .O(N__26166),
            .I(N__26160));
    Odrv12 I__5341 (
            .O(N__26163),
            .I(\POWERLED.un1_dutycycle_94_cry_13_c_RNIF6OBZ0Z1 ));
    Odrv12 I__5340 (
            .O(N__26160),
            .I(\POWERLED.un1_dutycycle_94_cry_13_c_RNIF6OBZ0Z1 ));
    InMux I__5339 (
            .O(N__26155),
            .I(N__26152));
    LocalMux I__5338 (
            .O(N__26152),
            .I(N__26149));
    Span4Mux_s2_h I__5337 (
            .O(N__26149),
            .I(N__26145));
    InMux I__5336 (
            .O(N__26148),
            .I(N__26142));
    Odrv4 I__5335 (
            .O(N__26145),
            .I(\POWERLED.dutycycle_eena_11 ));
    LocalMux I__5334 (
            .O(N__26142),
            .I(\POWERLED.dutycycle_eena_11 ));
    InMux I__5333 (
            .O(N__26137),
            .I(N__26134));
    LocalMux I__5332 (
            .O(N__26134),
            .I(N__26130));
    InMux I__5331 (
            .O(N__26133),
            .I(N__26127));
    Span4Mux_h I__5330 (
            .O(N__26130),
            .I(N__26124));
    LocalMux I__5329 (
            .O(N__26127),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    Odrv4 I__5328 (
            .O(N__26124),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    CascadeMux I__5327 (
            .O(N__26119),
            .I(\POWERLED.un1_dutycycle_53_8_a3_1_0_cascade_ ));
    CascadeMux I__5326 (
            .O(N__26116),
            .I(N__26111));
    InMux I__5325 (
            .O(N__26115),
            .I(N__26107));
    InMux I__5324 (
            .O(N__26114),
            .I(N__26102));
    InMux I__5323 (
            .O(N__26111),
            .I(N__26102));
    InMux I__5322 (
            .O(N__26110),
            .I(N__26099));
    LocalMux I__5321 (
            .O(N__26107),
            .I(N__26094));
    LocalMux I__5320 (
            .O(N__26102),
            .I(N__26091));
    LocalMux I__5319 (
            .O(N__26099),
            .I(N__26087));
    InMux I__5318 (
            .O(N__26098),
            .I(N__26084));
    InMux I__5317 (
            .O(N__26097),
            .I(N__26081));
    Span4Mux_v I__5316 (
            .O(N__26094),
            .I(N__26076));
    Span4Mux_h I__5315 (
            .O(N__26091),
            .I(N__26076));
    InMux I__5314 (
            .O(N__26090),
            .I(N__26073));
    Span4Mux_h I__5313 (
            .O(N__26087),
            .I(N__26068));
    LocalMux I__5312 (
            .O(N__26084),
            .I(N__26068));
    LocalMux I__5311 (
            .O(N__26081),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__5310 (
            .O(N__26076),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__5309 (
            .O(N__26073),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__5308 (
            .O(N__26068),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    CascadeMux I__5307 (
            .O(N__26059),
            .I(\POWERLED.un1_dutycycle_53_7_4_cascade_ ));
    CascadeMux I__5306 (
            .O(N__26056),
            .I(N__26053));
    InMux I__5305 (
            .O(N__26053),
            .I(N__26050));
    LocalMux I__5304 (
            .O(N__26050),
            .I(N__26047));
    Span4Mux_h I__5303 (
            .O(N__26047),
            .I(N__26044));
    Odrv4 I__5302 (
            .O(N__26044),
            .I(\POWERLED.dutycycle_RNIZ0Z_13 ));
    InMux I__5301 (
            .O(N__26041),
            .I(N__26038));
    LocalMux I__5300 (
            .O(N__26038),
            .I(\POWERLED.un1_N_5_mux ));
    CascadeMux I__5299 (
            .O(N__26035),
            .I(\POWERLED.un1_dutycycle_53_8_6_tz_sx_cascade_ ));
    InMux I__5298 (
            .O(N__26032),
            .I(N__26029));
    LocalMux I__5297 (
            .O(N__26029),
            .I(\POWERLED.un1_dutycycle_53_8_2_0_tz ));
    InMux I__5296 (
            .O(N__26026),
            .I(N__26023));
    LocalMux I__5295 (
            .O(N__26023),
            .I(N__26020));
    Odrv12 I__5294 (
            .O(N__26020),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_10 ));
    InMux I__5293 (
            .O(N__26017),
            .I(N__26011));
    InMux I__5292 (
            .O(N__26016),
            .I(N__26011));
    LocalMux I__5291 (
            .O(N__26011),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_9 ));
    InMux I__5290 (
            .O(N__26008),
            .I(N__26004));
    InMux I__5289 (
            .O(N__26007),
            .I(N__26001));
    LocalMux I__5288 (
            .O(N__26004),
            .I(N__25998));
    LocalMux I__5287 (
            .O(N__26001),
            .I(N__25995));
    Span4Mux_v I__5286 (
            .O(N__25998),
            .I(N__25992));
    Odrv12 I__5285 (
            .O(N__25995),
            .I(\POWERLED.mult1_un61_sum ));
    Odrv4 I__5284 (
            .O(N__25992),
            .I(\POWERLED.mult1_un61_sum ));
    InMux I__5283 (
            .O(N__25987),
            .I(N__25984));
    LocalMux I__5282 (
            .O(N__25984),
            .I(N__25981));
    Span4Mux_h I__5281 (
            .O(N__25981),
            .I(N__25978));
    Odrv4 I__5280 (
            .O(N__25978),
            .I(\POWERLED.mult1_un54_sum_i ));
    CascadeMux I__5279 (
            .O(N__25975),
            .I(N__25972));
    InMux I__5278 (
            .O(N__25972),
            .I(N__25969));
    LocalMux I__5277 (
            .O(N__25969),
            .I(\POWERLED.mult1_un61_sum_cry_3_s ));
    InMux I__5276 (
            .O(N__25966),
            .I(\POWERLED.mult1_un61_sum_cry_2 ));
    CascadeMux I__5275 (
            .O(N__25963),
            .I(N__25960));
    InMux I__5274 (
            .O(N__25960),
            .I(N__25957));
    LocalMux I__5273 (
            .O(N__25957),
            .I(N__25954));
    Span4Mux_s1_h I__5272 (
            .O(N__25954),
            .I(N__25951));
    Odrv4 I__5271 (
            .O(N__25951),
            .I(\POWERLED.mult1_un54_sum_cry_3_s ));
    InMux I__5270 (
            .O(N__25948),
            .I(N__25945));
    LocalMux I__5269 (
            .O(N__25945),
            .I(\POWERLED.mult1_un61_sum_cry_4_s ));
    InMux I__5268 (
            .O(N__25942),
            .I(\POWERLED.mult1_un61_sum_cry_3 ));
    InMux I__5267 (
            .O(N__25939),
            .I(N__25936));
    LocalMux I__5266 (
            .O(N__25936),
            .I(N__25933));
    Odrv4 I__5265 (
            .O(N__25933),
            .I(\POWERLED.mult1_un54_sum_cry_4_s ));
    CascadeMux I__5264 (
            .O(N__25930),
            .I(N__25927));
    InMux I__5263 (
            .O(N__25927),
            .I(N__25924));
    LocalMux I__5262 (
            .O(N__25924),
            .I(\POWERLED.mult1_un61_sum_cry_5_s ));
    InMux I__5261 (
            .O(N__25921),
            .I(\POWERLED.mult1_un61_sum_cry_4 ));
    CascadeMux I__5260 (
            .O(N__25918),
            .I(N__25914));
    InMux I__5259 (
            .O(N__25917),
            .I(N__25908));
    InMux I__5258 (
            .O(N__25914),
            .I(N__25908));
    InMux I__5257 (
            .O(N__25913),
            .I(N__25905));
    LocalMux I__5256 (
            .O(N__25908),
            .I(N__25901));
    LocalMux I__5255 (
            .O(N__25905),
            .I(N__25898));
    InMux I__5254 (
            .O(N__25904),
            .I(N__25895));
    Span4Mux_s2_h I__5253 (
            .O(N__25901),
            .I(N__25892));
    Span4Mux_s2_h I__5252 (
            .O(N__25898),
            .I(N__25889));
    LocalMux I__5251 (
            .O(N__25895),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    Odrv4 I__5250 (
            .O(N__25892),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    Odrv4 I__5249 (
            .O(N__25889),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    CascadeMux I__5248 (
            .O(N__25882),
            .I(N__25879));
    InMux I__5247 (
            .O(N__25879),
            .I(N__25876));
    LocalMux I__5246 (
            .O(N__25876),
            .I(N__25873));
    Odrv4 I__5245 (
            .O(N__25873),
            .I(\POWERLED.mult1_un54_sum_cry_5_s ));
    InMux I__5244 (
            .O(N__25870),
            .I(N__25867));
    LocalMux I__5243 (
            .O(N__25867),
            .I(\POWERLED.mult1_un61_sum_cry_6_s ));
    InMux I__5242 (
            .O(N__25864),
            .I(\POWERLED.mult1_un61_sum_cry_5 ));
    InMux I__5241 (
            .O(N__25861),
            .I(N__25858));
    LocalMux I__5240 (
            .O(N__25858),
            .I(N__25855));
    Odrv4 I__5239 (
            .O(N__25855),
            .I(\POWERLED.mult1_un54_sum_cry_6_s ));
    CascadeMux I__5238 (
            .O(N__25852),
            .I(N__25848));
    CascadeMux I__5237 (
            .O(N__25851),
            .I(N__25844));
    InMux I__5236 (
            .O(N__25848),
            .I(N__25837));
    InMux I__5235 (
            .O(N__25847),
            .I(N__25837));
    InMux I__5234 (
            .O(N__25844),
            .I(N__25837));
    LocalMux I__5233 (
            .O(N__25837),
            .I(\POWERLED.mult1_un54_sum_i_8 ));
    CascadeMux I__5232 (
            .O(N__25834),
            .I(N__25831));
    InMux I__5231 (
            .O(N__25831),
            .I(N__25828));
    LocalMux I__5230 (
            .O(N__25828),
            .I(\POWERLED.mult1_un68_sum_axb_8 ));
    InMux I__5229 (
            .O(N__25825),
            .I(\POWERLED.mult1_un61_sum_cry_6 ));
    CascadeMux I__5228 (
            .O(N__25822),
            .I(N__25819));
    InMux I__5227 (
            .O(N__25819),
            .I(N__25816));
    LocalMux I__5226 (
            .O(N__25816),
            .I(N__25813));
    Odrv4 I__5225 (
            .O(N__25813),
            .I(\POWERLED.mult1_un61_sum_axb_8 ));
    InMux I__5224 (
            .O(N__25810),
            .I(\POWERLED.mult1_un61_sum_cry_7 ));
    InMux I__5223 (
            .O(N__25807),
            .I(N__25804));
    LocalMux I__5222 (
            .O(N__25804),
            .I(N__25800));
    CascadeMux I__5221 (
            .O(N__25803),
            .I(N__25796));
    Span4Mux_h I__5220 (
            .O(N__25800),
            .I(N__25792));
    InMux I__5219 (
            .O(N__25799),
            .I(N__25787));
    InMux I__5218 (
            .O(N__25796),
            .I(N__25787));
    InMux I__5217 (
            .O(N__25795),
            .I(N__25784));
    Odrv4 I__5216 (
            .O(N__25792),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__5215 (
            .O(N__25787),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__5214 (
            .O(N__25784),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    CascadeMux I__5213 (
            .O(N__25777),
            .I(\POWERLED.mult1_un61_sum_s_8_cascade_ ));
    CascadeMux I__5212 (
            .O(N__25774),
            .I(N__25770));
    CascadeMux I__5211 (
            .O(N__25773),
            .I(N__25766));
    InMux I__5210 (
            .O(N__25770),
            .I(N__25759));
    InMux I__5209 (
            .O(N__25769),
            .I(N__25759));
    InMux I__5208 (
            .O(N__25766),
            .I(N__25759));
    LocalMux I__5207 (
            .O(N__25759),
            .I(\POWERLED.mult1_un61_sum_i_0_8 ));
    CascadeMux I__5206 (
            .O(N__25756),
            .I(N__25753));
    InMux I__5205 (
            .O(N__25753),
            .I(N__25750));
    LocalMux I__5204 (
            .O(N__25750),
            .I(N__25746));
    InMux I__5203 (
            .O(N__25749),
            .I(N__25743));
    Odrv4 I__5202 (
            .O(N__25746),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ));
    LocalMux I__5201 (
            .O(N__25743),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ));
    InMux I__5200 (
            .O(N__25738),
            .I(N__25735));
    LocalMux I__5199 (
            .O(N__25735),
            .I(N__25732));
    Span4Mux_h I__5198 (
            .O(N__25732),
            .I(N__25729));
    Odrv4 I__5197 (
            .O(N__25729),
            .I(\VPP_VDDQ.count_2_0_14 ));
    InMux I__5196 (
            .O(N__25726),
            .I(N__25722));
    InMux I__5195 (
            .O(N__25725),
            .I(N__25719));
    LocalMux I__5194 (
            .O(N__25722),
            .I(N__25716));
    LocalMux I__5193 (
            .O(N__25719),
            .I(N__25713));
    Span4Mux_h I__5192 (
            .O(N__25716),
            .I(N__25710));
    Odrv12 I__5191 (
            .O(N__25713),
            .I(\POWERLED.mult1_un68_sum ));
    Odrv4 I__5190 (
            .O(N__25710),
            .I(\POWERLED.mult1_un68_sum ));
    InMux I__5189 (
            .O(N__25705),
            .I(N__25702));
    LocalMux I__5188 (
            .O(N__25702),
            .I(N__25699));
    Span4Mux_s2_h I__5187 (
            .O(N__25699),
            .I(N__25696));
    Odrv4 I__5186 (
            .O(N__25696),
            .I(\POWERLED.mult1_un61_sum_i ));
    CascadeMux I__5185 (
            .O(N__25693),
            .I(N__25690));
    InMux I__5184 (
            .O(N__25690),
            .I(N__25687));
    LocalMux I__5183 (
            .O(N__25687),
            .I(N__25684));
    Odrv4 I__5182 (
            .O(N__25684),
            .I(\POWERLED.mult1_un68_sum_cry_3_s ));
    InMux I__5181 (
            .O(N__25681),
            .I(\POWERLED.mult1_un68_sum_cry_2 ));
    InMux I__5180 (
            .O(N__25678),
            .I(N__25675));
    LocalMux I__5179 (
            .O(N__25675),
            .I(N__25672));
    Odrv4 I__5178 (
            .O(N__25672),
            .I(\POWERLED.mult1_un68_sum_cry_4_s ));
    InMux I__5177 (
            .O(N__25669),
            .I(\POWERLED.mult1_un68_sum_cry_3 ));
    CascadeMux I__5176 (
            .O(N__25666),
            .I(N__25663));
    InMux I__5175 (
            .O(N__25663),
            .I(N__25660));
    LocalMux I__5174 (
            .O(N__25660),
            .I(N__25657));
    Odrv4 I__5173 (
            .O(N__25657),
            .I(\POWERLED.mult1_un68_sum_cry_5_s ));
    InMux I__5172 (
            .O(N__25654),
            .I(\POWERLED.mult1_un68_sum_cry_4 ));
    InMux I__5171 (
            .O(N__25651),
            .I(N__25648));
    LocalMux I__5170 (
            .O(N__25648),
            .I(N__25645));
    Odrv4 I__5169 (
            .O(N__25645),
            .I(\POWERLED.mult1_un68_sum_cry_6_s ));
    InMux I__5168 (
            .O(N__25642),
            .I(\POWERLED.mult1_un68_sum_cry_5 ));
    InMux I__5167 (
            .O(N__25639),
            .I(N__25636));
    LocalMux I__5166 (
            .O(N__25636),
            .I(N__25633));
    Odrv4 I__5165 (
            .O(N__25633),
            .I(\POWERLED.mult1_un75_sum_axb_8 ));
    InMux I__5164 (
            .O(N__25630),
            .I(\POWERLED.mult1_un68_sum_cry_6 ));
    InMux I__5163 (
            .O(N__25627),
            .I(\POWERLED.mult1_un68_sum_cry_7 ));
    CascadeMux I__5162 (
            .O(N__25624),
            .I(N__25619));
    InMux I__5161 (
            .O(N__25623),
            .I(N__25615));
    InMux I__5160 (
            .O(N__25622),
            .I(N__25609));
    InMux I__5159 (
            .O(N__25619),
            .I(N__25609));
    InMux I__5158 (
            .O(N__25618),
            .I(N__25606));
    LocalMux I__5157 (
            .O(N__25615),
            .I(N__25603));
    InMux I__5156 (
            .O(N__25614),
            .I(N__25600));
    LocalMux I__5155 (
            .O(N__25609),
            .I(N__25597));
    LocalMux I__5154 (
            .O(N__25606),
            .I(N__25594));
    Span4Mux_h I__5153 (
            .O(N__25603),
            .I(N__25585));
    LocalMux I__5152 (
            .O(N__25600),
            .I(N__25585));
    Span4Mux_s1_v I__5151 (
            .O(N__25597),
            .I(N__25585));
    Span4Mux_s1_v I__5150 (
            .O(N__25594),
            .I(N__25585));
    Odrv4 I__5149 (
            .O(N__25585),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    InMux I__5148 (
            .O(N__25582),
            .I(N__25576));
    InMux I__5147 (
            .O(N__25581),
            .I(N__25576));
    LocalMux I__5146 (
            .O(N__25576),
            .I(\VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ));
    InMux I__5145 (
            .O(N__25573),
            .I(N__25570));
    LocalMux I__5144 (
            .O(N__25570),
            .I(\VPP_VDDQ.count_2_0_10 ));
    CascadeMux I__5143 (
            .O(N__25567),
            .I(\VPP_VDDQ.count_2_1_10_cascade_ ));
    CascadeMux I__5142 (
            .O(N__25564),
            .I(\VPP_VDDQ.count_2_1_12_cascade_ ));
    InMux I__5141 (
            .O(N__25561),
            .I(N__25555));
    InMux I__5140 (
            .O(N__25560),
            .I(N__25555));
    LocalMux I__5139 (
            .O(N__25555),
            .I(N__25552));
    Odrv4 I__5138 (
            .O(N__25552),
            .I(\VPP_VDDQ.count_2Z0Z_12 ));
    InMux I__5137 (
            .O(N__25549),
            .I(N__25543));
    InMux I__5136 (
            .O(N__25548),
            .I(N__25543));
    LocalMux I__5135 (
            .O(N__25543),
            .I(N__25540));
    Odrv4 I__5134 (
            .O(N__25540),
            .I(\VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0 ));
    InMux I__5133 (
            .O(N__25537),
            .I(N__25534));
    LocalMux I__5132 (
            .O(N__25534),
            .I(\VPP_VDDQ.count_2_0_12 ));
    CascadeMux I__5131 (
            .O(N__25531),
            .I(\VPP_VDDQ.count_2_1_13_cascade_ ));
    InMux I__5130 (
            .O(N__25528),
            .I(N__25522));
    InMux I__5129 (
            .O(N__25527),
            .I(N__25522));
    LocalMux I__5128 (
            .O(N__25522),
            .I(N__25519));
    Odrv4 I__5127 (
            .O(N__25519),
            .I(\VPP_VDDQ.count_2Z0Z_13 ));
    InMux I__5126 (
            .O(N__25516),
            .I(N__25510));
    InMux I__5125 (
            .O(N__25515),
            .I(N__25510));
    LocalMux I__5124 (
            .O(N__25510),
            .I(N__25507));
    Odrv4 I__5123 (
            .O(N__25507),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ));
    InMux I__5122 (
            .O(N__25504),
            .I(N__25501));
    LocalMux I__5121 (
            .O(N__25501),
            .I(\VPP_VDDQ.count_2_0_13 ));
    InMux I__5120 (
            .O(N__25498),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12 ));
    InMux I__5119 (
            .O(N__25495),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13 ));
    InMux I__5118 (
            .O(N__25492),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14 ));
    InMux I__5117 (
            .O(N__25489),
            .I(N__25483));
    InMux I__5116 (
            .O(N__25488),
            .I(N__25483));
    LocalMux I__5115 (
            .O(N__25483),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ));
    InMux I__5114 (
            .O(N__25480),
            .I(N__25474));
    InMux I__5113 (
            .O(N__25479),
            .I(N__25474));
    LocalMux I__5112 (
            .O(N__25474),
            .I(\VPP_VDDQ.count_2Z0Z_15 ));
    CascadeMux I__5111 (
            .O(N__25471),
            .I(N__25468));
    InMux I__5110 (
            .O(N__25468),
            .I(N__25464));
    InMux I__5109 (
            .O(N__25467),
            .I(N__25461));
    LocalMux I__5108 (
            .O(N__25464),
            .I(\VPP_VDDQ.count_2Z0Z_14 ));
    LocalMux I__5107 (
            .O(N__25461),
            .I(\VPP_VDDQ.count_2Z0Z_14 ));
    InMux I__5106 (
            .O(N__25456),
            .I(N__25450));
    InMux I__5105 (
            .O(N__25455),
            .I(N__25450));
    LocalMux I__5104 (
            .O(N__25450),
            .I(N__25447));
    Odrv4 I__5103 (
            .O(N__25447),
            .I(\VPP_VDDQ.count_2_1_6 ));
    CascadeMux I__5102 (
            .O(N__25444),
            .I(N__25440));
    InMux I__5101 (
            .O(N__25443),
            .I(N__25435));
    InMux I__5100 (
            .O(N__25440),
            .I(N__25435));
    LocalMux I__5099 (
            .O(N__25435),
            .I(N__25432));
    Odrv4 I__5098 (
            .O(N__25432),
            .I(\VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661 ));
    InMux I__5097 (
            .O(N__25429),
            .I(N__25423));
    InMux I__5096 (
            .O(N__25428),
            .I(N__25423));
    LocalMux I__5095 (
            .O(N__25423),
            .I(N__25420));
    Odrv12 I__5094 (
            .O(N__25420),
            .I(\VPP_VDDQ.count_2Z0Z_6 ));
    CascadeMux I__5093 (
            .O(N__25417),
            .I(\VPP_VDDQ.count_2_1_9_cascade_ ));
    CascadeMux I__5092 (
            .O(N__25414),
            .I(N__25410));
    CascadeMux I__5091 (
            .O(N__25413),
            .I(N__25407));
    InMux I__5090 (
            .O(N__25410),
            .I(N__25402));
    InMux I__5089 (
            .O(N__25407),
            .I(N__25402));
    LocalMux I__5088 (
            .O(N__25402),
            .I(\VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ));
    InMux I__5087 (
            .O(N__25399),
            .I(N__25396));
    LocalMux I__5086 (
            .O(N__25396),
            .I(\VPP_VDDQ.count_2_0_9 ));
    InMux I__5085 (
            .O(N__25393),
            .I(N__25389));
    InMux I__5084 (
            .O(N__25392),
            .I(N__25386));
    LocalMux I__5083 (
            .O(N__25389),
            .I(\VPP_VDDQ.count_2Z0Z_5 ));
    LocalMux I__5082 (
            .O(N__25386),
            .I(\VPP_VDDQ.count_2Z0Z_5 ));
    CascadeMux I__5081 (
            .O(N__25381),
            .I(N__25377));
    InMux I__5080 (
            .O(N__25380),
            .I(N__25372));
    InMux I__5079 (
            .O(N__25377),
            .I(N__25372));
    LocalMux I__5078 (
            .O(N__25372),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7 ));
    InMux I__5077 (
            .O(N__25369),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4 ));
    InMux I__5076 (
            .O(N__25366),
            .I(N__25363));
    LocalMux I__5075 (
            .O(N__25363),
            .I(\VPP_VDDQ.un1_count_2_1_axb_6 ));
    InMux I__5074 (
            .O(N__25360),
            .I(\VPP_VDDQ.un1_count_2_1_cry_5 ));
    InMux I__5073 (
            .O(N__25357),
            .I(\VPP_VDDQ.un1_count_2_1_cry_6 ));
    InMux I__5072 (
            .O(N__25354),
            .I(N__25350));
    InMux I__5071 (
            .O(N__25353),
            .I(N__25347));
    LocalMux I__5070 (
            .O(N__25350),
            .I(N__25344));
    LocalMux I__5069 (
            .O(N__25347),
            .I(N__25341));
    Span4Mux_v I__5068 (
            .O(N__25344),
            .I(N__25336));
    Span4Mux_v I__5067 (
            .O(N__25341),
            .I(N__25336));
    Span4Mux_v I__5066 (
            .O(N__25336),
            .I(N__25333));
    Odrv4 I__5065 (
            .O(N__25333),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    InMux I__5064 (
            .O(N__25330),
            .I(N__25324));
    InMux I__5063 (
            .O(N__25329),
            .I(N__25324));
    LocalMux I__5062 (
            .O(N__25324),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7 ));
    InMux I__5061 (
            .O(N__25321),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7 ));
    InMux I__5060 (
            .O(N__25318),
            .I(bfn_9_14_0_));
    InMux I__5059 (
            .O(N__25315),
            .I(\VPP_VDDQ.un1_count_2_1_cry_9 ));
    InMux I__5058 (
            .O(N__25312),
            .I(\VPP_VDDQ.un1_count_2_1_cry_10 ));
    InMux I__5057 (
            .O(N__25309),
            .I(\VPP_VDDQ.un1_count_2_1_cry_11 ));
    IoInMux I__5056 (
            .O(N__25306),
            .I(N__25303));
    LocalMux I__5055 (
            .O(N__25303),
            .I(N__25300));
    IoSpan4Mux I__5054 (
            .O(N__25300),
            .I(N__25297));
    IoSpan4Mux I__5053 (
            .O(N__25297),
            .I(N__25294));
    Span4Mux_s3_h I__5052 (
            .O(N__25294),
            .I(N__25290));
    InMux I__5051 (
            .O(N__25293),
            .I(N__25287));
    Sp12to4 I__5050 (
            .O(N__25290),
            .I(N__25282));
    LocalMux I__5049 (
            .O(N__25287),
            .I(N__25282));
    Odrv12 I__5048 (
            .O(N__25282),
            .I(v1p8a_ok));
    InMux I__5047 (
            .O(N__25279),
            .I(N__25276));
    LocalMux I__5046 (
            .O(N__25276),
            .I(N__25273));
    Span4Mux_v I__5045 (
            .O(N__25273),
            .I(N__25270));
    Span4Mux_h I__5044 (
            .O(N__25270),
            .I(N__25267));
    Span4Mux_h I__5043 (
            .O(N__25267),
            .I(N__25264));
    Span4Mux_v I__5042 (
            .O(N__25264),
            .I(N__25261));
    Odrv4 I__5041 (
            .O(N__25261),
            .I(v5a_ok));
    CascadeMux I__5040 (
            .O(N__25258),
            .I(N_171_cascade_));
    InMux I__5039 (
            .O(N__25255),
            .I(N__25252));
    LocalMux I__5038 (
            .O(N__25252),
            .I(N__25249));
    Span4Mux_v I__5037 (
            .O(N__25249),
            .I(N__25246));
    Span4Mux_v I__5036 (
            .O(N__25246),
            .I(N__25243));
    Odrv4 I__5035 (
            .O(N__25243),
            .I(vr_ready_vccinaux));
    InMux I__5034 (
            .O(N__25240),
            .I(N__25224));
    InMux I__5033 (
            .O(N__25239),
            .I(N__25224));
    InMux I__5032 (
            .O(N__25238),
            .I(N__25224));
    InMux I__5031 (
            .O(N__25237),
            .I(N__25224));
    InMux I__5030 (
            .O(N__25236),
            .I(N__25224));
    InMux I__5029 (
            .O(N__25235),
            .I(N__25221));
    LocalMux I__5028 (
            .O(N__25224),
            .I(N_283));
    LocalMux I__5027 (
            .O(N__25221),
            .I(N_283));
    InMux I__5026 (
            .O(N__25216),
            .I(N__25199));
    InMux I__5025 (
            .O(N__25215),
            .I(N__25199));
    InMux I__5024 (
            .O(N__25214),
            .I(N__25199));
    InMux I__5023 (
            .O(N__25213),
            .I(N__25199));
    InMux I__5022 (
            .O(N__25212),
            .I(N__25199));
    InMux I__5021 (
            .O(N__25211),
            .I(N__25194));
    InMux I__5020 (
            .O(N__25210),
            .I(N__25194));
    LocalMux I__5019 (
            .O(N__25199),
            .I(RSMRST_PWRGD_curr_state_0));
    LocalMux I__5018 (
            .O(N__25194),
            .I(RSMRST_PWRGD_curr_state_0));
    CascadeMux I__5017 (
            .O(N__25189),
            .I(N_283_cascade_));
    CascadeMux I__5016 (
            .O(N__25186),
            .I(N__25181));
    InMux I__5015 (
            .O(N__25185),
            .I(N__25172));
    InMux I__5014 (
            .O(N__25184),
            .I(N__25172));
    InMux I__5013 (
            .O(N__25181),
            .I(N__25165));
    InMux I__5012 (
            .O(N__25180),
            .I(N__25165));
    InMux I__5011 (
            .O(N__25179),
            .I(N__25165));
    InMux I__5010 (
            .O(N__25178),
            .I(N__25160));
    InMux I__5009 (
            .O(N__25177),
            .I(N__25160));
    LocalMux I__5008 (
            .O(N__25172),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__5007 (
            .O(N__25165),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__5006 (
            .O(N__25160),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    IoInMux I__5005 (
            .O(N__25153),
            .I(N__25150));
    LocalMux I__5004 (
            .O(N__25150),
            .I(N__25147));
    IoSpan4Mux I__5003 (
            .O(N__25147),
            .I(N__25140));
    InMux I__5002 (
            .O(N__25146),
            .I(N__25137));
    CascadeMux I__5001 (
            .O(N__25145),
            .I(N__25133));
    InMux I__5000 (
            .O(N__25144),
            .I(N__25129));
    InMux I__4999 (
            .O(N__25143),
            .I(N__25126));
    Span4Mux_s2_v I__4998 (
            .O(N__25140),
            .I(N__25119));
    LocalMux I__4997 (
            .O(N__25137),
            .I(N__25119));
    InMux I__4996 (
            .O(N__25136),
            .I(N__25112));
    InMux I__4995 (
            .O(N__25133),
            .I(N__25112));
    InMux I__4994 (
            .O(N__25132),
            .I(N__25112));
    LocalMux I__4993 (
            .O(N__25129),
            .I(N__25109));
    LocalMux I__4992 (
            .O(N__25126),
            .I(N__25106));
    InMux I__4991 (
            .O(N__25125),
            .I(N__25103));
    InMux I__4990 (
            .O(N__25124),
            .I(N__25100));
    Span4Mux_v I__4989 (
            .O(N__25119),
            .I(N__25096));
    LocalMux I__4988 (
            .O(N__25112),
            .I(N__25093));
    Span4Mux_h I__4987 (
            .O(N__25109),
            .I(N__25086));
    Span4Mux_v I__4986 (
            .O(N__25106),
            .I(N__25086));
    LocalMux I__4985 (
            .O(N__25103),
            .I(N__25086));
    LocalMux I__4984 (
            .O(N__25100),
            .I(N__25083));
    InMux I__4983 (
            .O(N__25099),
            .I(N__25080));
    Span4Mux_h I__4982 (
            .O(N__25096),
            .I(N__25073));
    Span4Mux_v I__4981 (
            .O(N__25093),
            .I(N__25073));
    Span4Mux_h I__4980 (
            .O(N__25086),
            .I(N__25073));
    Odrv4 I__4979 (
            .O(N__25083),
            .I(rsmrstn));
    LocalMux I__4978 (
            .O(N__25080),
            .I(rsmrstn));
    Odrv4 I__4977 (
            .O(N__25073),
            .I(rsmrstn));
    InMux I__4976 (
            .O(N__25066),
            .I(N__25063));
    LocalMux I__4975 (
            .O(N__25063),
            .I(\VPP_VDDQ.un9_clk_100khz_9 ));
    CascadeMux I__4974 (
            .O(N__25060),
            .I(\VPP_VDDQ.un9_clk_100khz_0_cascade_ ));
    InMux I__4973 (
            .O(N__25057),
            .I(N__25054));
    LocalMux I__4972 (
            .O(N__25054),
            .I(\VPP_VDDQ.count_2Z0Z_2 ));
    CascadeMux I__4971 (
            .O(N__25051),
            .I(N__25047));
    InMux I__4970 (
            .O(N__25050),
            .I(N__25042));
    InMux I__4969 (
            .O(N__25047),
            .I(N__25042));
    LocalMux I__4968 (
            .O(N__25042),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087 ));
    InMux I__4967 (
            .O(N__25039),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1 ));
    InMux I__4966 (
            .O(N__25036),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2 ));
    InMux I__4965 (
            .O(N__25033),
            .I(N__25029));
    InMux I__4964 (
            .O(N__25032),
            .I(N__25026));
    LocalMux I__4963 (
            .O(N__25029),
            .I(\VPP_VDDQ.count_2Z0Z_4 ));
    LocalMux I__4962 (
            .O(N__25026),
            .I(\VPP_VDDQ.count_2Z0Z_4 ));
    InMux I__4961 (
            .O(N__25021),
            .I(N__25015));
    InMux I__4960 (
            .O(N__25020),
            .I(N__25015));
    LocalMux I__4959 (
            .O(N__25015),
            .I(\VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7 ));
    InMux I__4958 (
            .O(N__25012),
            .I(\VPP_VDDQ.un1_count_2_1_cry_3 ));
    IoInMux I__4957 (
            .O(N__25009),
            .I(N__25005));
    InMux I__4956 (
            .O(N__25008),
            .I(N__25001));
    LocalMux I__4955 (
            .O(N__25005),
            .I(N__24996));
    IoInMux I__4954 (
            .O(N__25004),
            .I(N__24992));
    LocalMux I__4953 (
            .O(N__25001),
            .I(N__24989));
    InMux I__4952 (
            .O(N__25000),
            .I(N__24986));
    InMux I__4951 (
            .O(N__24999),
            .I(N__24983));
    Span4Mux_s0_h I__4950 (
            .O(N__24996),
            .I(N__24980));
    InMux I__4949 (
            .O(N__24995),
            .I(N__24977));
    LocalMux I__4948 (
            .O(N__24992),
            .I(N__24973));
    Span4Mux_v I__4947 (
            .O(N__24989),
            .I(N__24970));
    LocalMux I__4946 (
            .O(N__24986),
            .I(N__24967));
    LocalMux I__4945 (
            .O(N__24983),
            .I(N__24963));
    Span4Mux_h I__4944 (
            .O(N__24980),
            .I(N__24958));
    LocalMux I__4943 (
            .O(N__24977),
            .I(N__24958));
    InMux I__4942 (
            .O(N__24976),
            .I(N__24955));
    Span4Mux_s2_h I__4941 (
            .O(N__24973),
            .I(N__24946));
    Span4Mux_v I__4940 (
            .O(N__24970),
            .I(N__24946));
    Span4Mux_v I__4939 (
            .O(N__24967),
            .I(N__24946));
    InMux I__4938 (
            .O(N__24966),
            .I(N__24943));
    Span4Mux_h I__4937 (
            .O(N__24963),
            .I(N__24936));
    Span4Mux_v I__4936 (
            .O(N__24958),
            .I(N__24936));
    LocalMux I__4935 (
            .O(N__24955),
            .I(N__24936));
    InMux I__4934 (
            .O(N__24954),
            .I(N__24931));
    InMux I__4933 (
            .O(N__24953),
            .I(N__24928));
    Span4Mux_h I__4932 (
            .O(N__24946),
            .I(N__24925));
    LocalMux I__4931 (
            .O(N__24943),
            .I(N__24922));
    Span4Mux_h I__4930 (
            .O(N__24936),
            .I(N__24919));
    InMux I__4929 (
            .O(N__24935),
            .I(N__24914));
    InMux I__4928 (
            .O(N__24934),
            .I(N__24914));
    LocalMux I__4927 (
            .O(N__24931),
            .I(v5s_enn));
    LocalMux I__4926 (
            .O(N__24928),
            .I(v5s_enn));
    Odrv4 I__4925 (
            .O(N__24925),
            .I(v5s_enn));
    Odrv4 I__4924 (
            .O(N__24922),
            .I(v5s_enn));
    Odrv4 I__4923 (
            .O(N__24919),
            .I(v5s_enn));
    LocalMux I__4922 (
            .O(N__24914),
            .I(v5s_enn));
    CascadeMux I__4921 (
            .O(N__24901),
            .I(\VCCIN_PWRGD.un10_outputZ0Z_3_cascade_ ));
    IoInMux I__4920 (
            .O(N__24898),
            .I(N__24895));
    LocalMux I__4919 (
            .O(N__24895),
            .I(N__24892));
    Span4Mux_s3_v I__4918 (
            .O(N__24892),
            .I(N__24889));
    Odrv4 I__4917 (
            .O(N__24889),
            .I(vccin_en));
    InMux I__4916 (
            .O(N__24886),
            .I(N__24883));
    LocalMux I__4915 (
            .O(N__24883),
            .I(N_323));
    CascadeMux I__4914 (
            .O(N__24880),
            .I(N_323_cascade_));
    IoInMux I__4913 (
            .O(N__24877),
            .I(N__24874));
    LocalMux I__4912 (
            .O(N__24874),
            .I(N__24871));
    Span4Mux_s3_h I__4911 (
            .O(N__24871),
            .I(N__24867));
    InMux I__4910 (
            .O(N__24870),
            .I(N__24864));
    Span4Mux_h I__4909 (
            .O(N__24867),
            .I(N__24861));
    LocalMux I__4908 (
            .O(N__24864),
            .I(N__24857));
    Sp12to4 I__4907 (
            .O(N__24861),
            .I(N__24854));
    InMux I__4906 (
            .O(N__24860),
            .I(N__24851));
    Span4Mux_v I__4905 (
            .O(N__24857),
            .I(N__24848));
    Span12Mux_v I__4904 (
            .O(N__24854),
            .I(N__24843));
    LocalMux I__4903 (
            .O(N__24851),
            .I(N__24843));
    Odrv4 I__4902 (
            .O(N__24848),
            .I(v33a_ok));
    Odrv12 I__4901 (
            .O(N__24843),
            .I(v33a_ok));
    InMux I__4900 (
            .O(N__24838),
            .I(N__24834));
    InMux I__4899 (
            .O(N__24837),
            .I(N__24831));
    LocalMux I__4898 (
            .O(N__24834),
            .I(N__24828));
    LocalMux I__4897 (
            .O(N__24831),
            .I(N__24825));
    Odrv12 I__4896 (
            .O(N__24828),
            .I(slp_susn));
    Odrv4 I__4895 (
            .O(N__24825),
            .I(slp_susn));
    InMux I__4894 (
            .O(N__24820),
            .I(N__24817));
    LocalMux I__4893 (
            .O(N__24817),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_6 ));
    InMux I__4892 (
            .O(N__24814),
            .I(N__24809));
    InMux I__4891 (
            .O(N__24813),
            .I(N__24802));
    InMux I__4890 (
            .O(N__24812),
            .I(N__24802));
    LocalMux I__4889 (
            .O(N__24809),
            .I(N__24799));
    CascadeMux I__4888 (
            .O(N__24808),
            .I(N__24794));
    CascadeMux I__4887 (
            .O(N__24807),
            .I(N__24791));
    LocalMux I__4886 (
            .O(N__24802),
            .I(N__24788));
    Span4Mux_v I__4885 (
            .O(N__24799),
            .I(N__24785));
    InMux I__4884 (
            .O(N__24798),
            .I(N__24780));
    InMux I__4883 (
            .O(N__24797),
            .I(N__24780));
    InMux I__4882 (
            .O(N__24794),
            .I(N__24777));
    InMux I__4881 (
            .O(N__24791),
            .I(N__24774));
    Span4Mux_h I__4880 (
            .O(N__24788),
            .I(N__24771));
    Span4Mux_h I__4879 (
            .O(N__24785),
            .I(N__24766));
    LocalMux I__4878 (
            .O(N__24780),
            .I(N__24766));
    LocalMux I__4877 (
            .O(N__24777),
            .I(\POWERLED.N_258 ));
    LocalMux I__4876 (
            .O(N__24774),
            .I(\POWERLED.N_258 ));
    Odrv4 I__4875 (
            .O(N__24771),
            .I(\POWERLED.N_258 ));
    Odrv4 I__4874 (
            .O(N__24766),
            .I(\POWERLED.N_258 ));
    InMux I__4873 (
            .O(N__24757),
            .I(N__24754));
    LocalMux I__4872 (
            .O(N__24754),
            .I(N__24750));
    InMux I__4871 (
            .O(N__24753),
            .I(N__24747));
    Odrv4 I__4870 (
            .O(N__24750),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_5 ));
    LocalMux I__4869 (
            .O(N__24747),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_5 ));
    InMux I__4868 (
            .O(N__24742),
            .I(N__24736));
    InMux I__4867 (
            .O(N__24741),
            .I(N__24733));
    InMux I__4866 (
            .O(N__24740),
            .I(N__24728));
    InMux I__4865 (
            .O(N__24739),
            .I(N__24728));
    LocalMux I__4864 (
            .O(N__24736),
            .I(N__24725));
    LocalMux I__4863 (
            .O(N__24733),
            .I(N__24718));
    LocalMux I__4862 (
            .O(N__24728),
            .I(N__24718));
    Span4Mux_v I__4861 (
            .O(N__24725),
            .I(N__24715));
    InMux I__4860 (
            .O(N__24724),
            .I(N__24710));
    InMux I__4859 (
            .O(N__24723),
            .I(N__24710));
    Span4Mux_h I__4858 (
            .O(N__24718),
            .I(N__24707));
    Odrv4 I__4857 (
            .O(N__24715),
            .I(\POWERLED.N_505 ));
    LocalMux I__4856 (
            .O(N__24710),
            .I(\POWERLED.N_505 ));
    Odrv4 I__4855 (
            .O(N__24707),
            .I(\POWERLED.N_505 ));
    CascadeMux I__4854 (
            .O(N__24700),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_5_cascade_ ));
    InMux I__4853 (
            .O(N__24697),
            .I(N__24694));
    LocalMux I__4852 (
            .O(N__24694),
            .I(\POWERLED.dutycycle_RNI2O4A1Z0Z_6 ));
    CascadeMux I__4851 (
            .O(N__24691),
            .I(\POWERLED.func_state_RNIOGRS_0Z0Z_1_cascade_ ));
    InMux I__4850 (
            .O(N__24688),
            .I(N__24685));
    LocalMux I__4849 (
            .O(N__24685),
            .I(N__24680));
    InMux I__4848 (
            .O(N__24684),
            .I(N__24677));
    InMux I__4847 (
            .O(N__24683),
            .I(N__24674));
    Span4Mux_h I__4846 (
            .O(N__24680),
            .I(N__24669));
    LocalMux I__4845 (
            .O(N__24677),
            .I(N__24669));
    LocalMux I__4844 (
            .O(N__24674),
            .I(N__24666));
    Span4Mux_h I__4843 (
            .O(N__24669),
            .I(N__24663));
    Odrv12 I__4842 (
            .O(N__24666),
            .I(\POWERLED.N_487 ));
    Odrv4 I__4841 (
            .O(N__24663),
            .I(\POWERLED.N_487 ));
    CascadeMux I__4840 (
            .O(N__24658),
            .I(\POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ));
    InMux I__4839 (
            .O(N__24655),
            .I(N__24648));
    InMux I__4838 (
            .O(N__24654),
            .I(N__24648));
    InMux I__4837 (
            .O(N__24653),
            .I(N__24645));
    LocalMux I__4836 (
            .O(N__24648),
            .I(N__24642));
    LocalMux I__4835 (
            .O(N__24645),
            .I(\POWERLED.N_379_N ));
    Odrv4 I__4834 (
            .O(N__24642),
            .I(\POWERLED.N_379_N ));
    InMux I__4833 (
            .O(N__24637),
            .I(N__24634));
    LocalMux I__4832 (
            .O(N__24634),
            .I(G_22_i_a2_1));
    InMux I__4831 (
            .O(N__24631),
            .I(N__24628));
    LocalMux I__4830 (
            .O(N__24628),
            .I(N__24623));
    InMux I__4829 (
            .O(N__24627),
            .I(N__24618));
    InMux I__4828 (
            .O(N__24626),
            .I(N__24618));
    Span4Mux_h I__4827 (
            .O(N__24623),
            .I(N__24615));
    LocalMux I__4826 (
            .O(N__24618),
            .I(SUSWARN_N_fast));
    Odrv4 I__4825 (
            .O(N__24615),
            .I(SUSWARN_N_fast));
    InMux I__4824 (
            .O(N__24610),
            .I(N__24604));
    InMux I__4823 (
            .O(N__24609),
            .I(N__24604));
    LocalMux I__4822 (
            .O(N__24604),
            .I(\POWERLED.N_564 ));
    InMux I__4821 (
            .O(N__24601),
            .I(N__24598));
    LocalMux I__4820 (
            .O(N__24598),
            .I(N__24595));
    Span4Mux_v I__4819 (
            .O(N__24595),
            .I(N__24592));
    Span4Mux_v I__4818 (
            .O(N__24592),
            .I(N__24589));
    Odrv4 I__4817 (
            .O(N__24589),
            .I(v5s_ok));
    InMux I__4816 (
            .O(N__24586),
            .I(N__24583));
    LocalMux I__4815 (
            .O(N__24583),
            .I(N__24580));
    Sp12to4 I__4814 (
            .O(N__24580),
            .I(N__24577));
    Span12Mux_v I__4813 (
            .O(N__24577),
            .I(N__24574));
    Odrv12 I__4812 (
            .O(N__24574),
            .I(vccst_cpu_ok));
    CascadeMux I__4811 (
            .O(N__24571),
            .I(N__24568));
    InMux I__4810 (
            .O(N__24568),
            .I(N__24565));
    LocalMux I__4809 (
            .O(N__24565),
            .I(N__24562));
    Span4Mux_v I__4808 (
            .O(N__24562),
            .I(N__24559));
    Odrv4 I__4807 (
            .O(N__24559),
            .I(v33s_ok));
    IoInMux I__4806 (
            .O(N__24556),
            .I(N__24552));
    InMux I__4805 (
            .O(N__24555),
            .I(N__24549));
    LocalMux I__4804 (
            .O(N__24552),
            .I(N__24546));
    LocalMux I__4803 (
            .O(N__24549),
            .I(N__24543));
    IoSpan4Mux I__4802 (
            .O(N__24546),
            .I(N__24540));
    Span12Mux_v I__4801 (
            .O(N__24543),
            .I(N__24537));
    Span4Mux_s1_h I__4800 (
            .O(N__24540),
            .I(N__24534));
    Odrv12 I__4799 (
            .O(N__24537),
            .I(dsw_pwrok));
    Odrv4 I__4798 (
            .O(N__24534),
            .I(dsw_pwrok));
    InMux I__4797 (
            .O(N__24529),
            .I(\POWERLED.un1_dutycycle_94_cry_11 ));
    CascadeMux I__4796 (
            .O(N__24526),
            .I(N__24522));
    InMux I__4795 (
            .O(N__24525),
            .I(N__24517));
    InMux I__4794 (
            .O(N__24522),
            .I(N__24517));
    LocalMux I__4793 (
            .O(N__24517),
            .I(N__24514));
    Odrv4 I__4792 (
            .O(N__24514),
            .I(\POWERLED.un1_dutycycle_94_cry_12_c_RNIE4NBZ0Z1 ));
    InMux I__4791 (
            .O(N__24511),
            .I(\POWERLED.un1_dutycycle_94_cry_12 ));
    CascadeMux I__4790 (
            .O(N__24508),
            .I(N__24503));
    CascadeMux I__4789 (
            .O(N__24507),
            .I(N__24496));
    InMux I__4788 (
            .O(N__24506),
            .I(N__24489));
    InMux I__4787 (
            .O(N__24503),
            .I(N__24476));
    InMux I__4786 (
            .O(N__24502),
            .I(N__24476));
    InMux I__4785 (
            .O(N__24501),
            .I(N__24476));
    InMux I__4784 (
            .O(N__24500),
            .I(N__24476));
    InMux I__4783 (
            .O(N__24499),
            .I(N__24476));
    InMux I__4782 (
            .O(N__24496),
            .I(N__24476));
    CascadeMux I__4781 (
            .O(N__24495),
            .I(N__24473));
    CascadeMux I__4780 (
            .O(N__24494),
            .I(N__24469));
    CascadeMux I__4779 (
            .O(N__24493),
            .I(N__24465));
    CascadeMux I__4778 (
            .O(N__24492),
            .I(N__24461));
    LocalMux I__4777 (
            .O(N__24489),
            .I(N__24456));
    LocalMux I__4776 (
            .O(N__24476),
            .I(N__24456));
    InMux I__4775 (
            .O(N__24473),
            .I(N__24451));
    InMux I__4774 (
            .O(N__24472),
            .I(N__24451));
    InMux I__4773 (
            .O(N__24469),
            .I(N__24440));
    InMux I__4772 (
            .O(N__24468),
            .I(N__24440));
    InMux I__4771 (
            .O(N__24465),
            .I(N__24440));
    InMux I__4770 (
            .O(N__24464),
            .I(N__24440));
    InMux I__4769 (
            .O(N__24461),
            .I(N__24440));
    Span4Mux_h I__4768 (
            .O(N__24456),
            .I(N__24437));
    LocalMux I__4767 (
            .O(N__24451),
            .I(N__24432));
    LocalMux I__4766 (
            .O(N__24440),
            .I(N__24432));
    Odrv4 I__4765 (
            .O(N__24437),
            .I(\POWERLED.N_341_i ));
    Odrv12 I__4764 (
            .O(N__24432),
            .I(\POWERLED.N_341_i ));
    InMux I__4763 (
            .O(N__24427),
            .I(\POWERLED.un1_dutycycle_94_cry_13 ));
    InMux I__4762 (
            .O(N__24424),
            .I(\POWERLED.un1_dutycycle_94_cry_14 ));
    InMux I__4761 (
            .O(N__24421),
            .I(N__24415));
    InMux I__4760 (
            .O(N__24420),
            .I(N__24415));
    LocalMux I__4759 (
            .O(N__24415),
            .I(\POWERLED.un1_dutycycle_94_cry_14_c_RNIG8PBZ0Z1 ));
    InMux I__4758 (
            .O(N__24412),
            .I(N__24409));
    LocalMux I__4757 (
            .O(N__24409),
            .I(N__24406));
    Span4Mux_h I__4756 (
            .O(N__24406),
            .I(N__24402));
    InMux I__4755 (
            .O(N__24405),
            .I(N__24399));
    Span4Mux_v I__4754 (
            .O(N__24402),
            .I(N__24396));
    LocalMux I__4753 (
            .O(N__24399),
            .I(N__24393));
    Odrv4 I__4752 (
            .O(N__24396),
            .I(\POWERLED.N_292 ));
    Odrv4 I__4751 (
            .O(N__24393),
            .I(\POWERLED.N_292 ));
    CascadeMux I__4750 (
            .O(N__24388),
            .I(\POWERLED.dutycycle_1_0_iv_i_a3_0_2_cascade_ ));
    InMux I__4749 (
            .O(N__24385),
            .I(N__24382));
    LocalMux I__4748 (
            .O(N__24382),
            .I(N__24379));
    Odrv4 I__4747 (
            .O(N__24379),
            .I(\POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ));
    InMux I__4746 (
            .O(N__24376),
            .I(N__24370));
    InMux I__4745 (
            .O(N__24375),
            .I(N__24370));
    LocalMux I__4744 (
            .O(N__24370),
            .I(\POWERLED.N_145 ));
    InMux I__4743 (
            .O(N__24367),
            .I(N__24364));
    LocalMux I__4742 (
            .O(N__24364),
            .I(N__24361));
    Span4Mux_v I__4741 (
            .O(N__24361),
            .I(N__24358));
    Odrv4 I__4740 (
            .O(N__24358),
            .I(m57_i_o2_3));
    CascadeMux I__4739 (
            .O(N__24355),
            .I(N__24352));
    InMux I__4738 (
            .O(N__24352),
            .I(N__24349));
    LocalMux I__4737 (
            .O(N__24349),
            .I(N__24346));
    Odrv4 I__4736 (
            .O(N__24346),
            .I(\POWERLED.un1_dutycycle_94_cry_5_c_RNIZ0 ));
    InMux I__4735 (
            .O(N__24343),
            .I(N__24340));
    LocalMux I__4734 (
            .O(N__24340),
            .I(N__24337));
    Span12Mux_s8_h I__4733 (
            .O(N__24337),
            .I(N__24333));
    InMux I__4732 (
            .O(N__24336),
            .I(N__24330));
    Odrv12 I__4731 (
            .O(N__24333),
            .I(\POWERLED.un1_dutycycle_94_cry_5_c_RNIEVTSZ0Z3 ));
    LocalMux I__4730 (
            .O(N__24330),
            .I(\POWERLED.un1_dutycycle_94_cry_5_c_RNIEVTSZ0Z3 ));
    InMux I__4729 (
            .O(N__24325),
            .I(N__24322));
    LocalMux I__4728 (
            .O(N__24322),
            .I(N__24319));
    Odrv4 I__4727 (
            .O(N__24319),
            .I(\POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ));
    InMux I__4726 (
            .O(N__24316),
            .I(N__24310));
    InMux I__4725 (
            .O(N__24315),
            .I(N__24310));
    LocalMux I__4724 (
            .O(N__24310),
            .I(\POWERLED.dutycycle_set_1 ));
    InMux I__4723 (
            .O(N__24307),
            .I(N__24301));
    InMux I__4722 (
            .O(N__24306),
            .I(N__24301));
    LocalMux I__4721 (
            .O(N__24301),
            .I(N__24298));
    Span4Mux_h I__4720 (
            .O(N__24298),
            .I(N__24295));
    Span4Mux_v I__4719 (
            .O(N__24295),
            .I(N__24292));
    Odrv4 I__4718 (
            .O(N__24292),
            .I(\POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ));
    InMux I__4717 (
            .O(N__24289),
            .I(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ));
    InMux I__4716 (
            .O(N__24286),
            .I(N__24280));
    InMux I__4715 (
            .O(N__24285),
            .I(N__24280));
    LocalMux I__4714 (
            .O(N__24280),
            .I(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ));
    InMux I__4713 (
            .O(N__24277),
            .I(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ));
    InMux I__4712 (
            .O(N__24274),
            .I(\POWERLED.un1_dutycycle_94_cry_4 ));
    InMux I__4711 (
            .O(N__24271),
            .I(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ));
    InMux I__4710 (
            .O(N__24268),
            .I(N__24265));
    LocalMux I__4709 (
            .O(N__24265),
            .I(N__24261));
    InMux I__4708 (
            .O(N__24264),
            .I(N__24258));
    Span4Mux_s2_v I__4707 (
            .O(N__24261),
            .I(N__24255));
    LocalMux I__4706 (
            .O(N__24258),
            .I(N__24252));
    Span4Mux_v I__4705 (
            .O(N__24255),
            .I(N__24249));
    Span4Mux_h I__4704 (
            .O(N__24252),
            .I(N__24246));
    Odrv4 I__4703 (
            .O(N__24249),
            .I(\POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ));
    Odrv4 I__4702 (
            .O(N__24246),
            .I(\POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ));
    InMux I__4701 (
            .O(N__24241),
            .I(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ));
    InMux I__4700 (
            .O(N__24238),
            .I(bfn_9_8_0_));
    InMux I__4699 (
            .O(N__24235),
            .I(N__24229));
    InMux I__4698 (
            .O(N__24234),
            .I(N__24229));
    LocalMux I__4697 (
            .O(N__24229),
            .I(N__24226));
    Odrv4 I__4696 (
            .O(N__24226),
            .I(\POWERLED.un1_dutycycle_94_cry_8_c_RNI3B2UZ0 ));
    InMux I__4695 (
            .O(N__24223),
            .I(\POWERLED.un1_dutycycle_94_cry_8 ));
    InMux I__4694 (
            .O(N__24220),
            .I(\POWERLED.un1_dutycycle_94_cry_9 ));
    InMux I__4693 (
            .O(N__24217),
            .I(\POWERLED.un1_dutycycle_94_cry_10 ));
    CascadeMux I__4692 (
            .O(N__24214),
            .I(\POWERLED.dutycycleZ0Z_9_cascade_ ));
    CascadeMux I__4691 (
            .O(N__24211),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_13_cascade_ ));
    CascadeMux I__4690 (
            .O(N__24208),
            .I(N__24205));
    InMux I__4689 (
            .O(N__24205),
            .I(N__24202));
    LocalMux I__4688 (
            .O(N__24202),
            .I(N__24199));
    Span4Mux_h I__4687 (
            .O(N__24199),
            .I(N__24196));
    Odrv4 I__4686 (
            .O(N__24196),
            .I(\POWERLED.dutycycle_RNIZ0Z_14 ));
    InMux I__4685 (
            .O(N__24193),
            .I(N__24190));
    LocalMux I__4684 (
            .O(N__24190),
            .I(\POWERLED.un1_dutycycle_53_12_0 ));
    InMux I__4683 (
            .O(N__24187),
            .I(N__24184));
    LocalMux I__4682 (
            .O(N__24184),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_13 ));
    CascadeMux I__4681 (
            .O(N__24181),
            .I(N__24178));
    InMux I__4680 (
            .O(N__24178),
            .I(N__24175));
    LocalMux I__4679 (
            .O(N__24175),
            .I(N__24172));
    Odrv4 I__4678 (
            .O(N__24172),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_14 ));
    InMux I__4677 (
            .O(N__24169),
            .I(N__24166));
    LocalMux I__4676 (
            .O(N__24166),
            .I(N__24163));
    Odrv4 I__4675 (
            .O(N__24163),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_7 ));
    CascadeMux I__4674 (
            .O(N__24160),
            .I(\POWERLED.un1_dutycycle_53_57_a0_d_cascade_ ));
    InMux I__4673 (
            .O(N__24157),
            .I(N__24154));
    LocalMux I__4672 (
            .O(N__24154),
            .I(N__24151));
    Odrv4 I__4671 (
            .O(N__24151),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_13 ));
    InMux I__4670 (
            .O(N__24148),
            .I(N__24145));
    LocalMux I__4669 (
            .O(N__24145),
            .I(\POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ));
    InMux I__4668 (
            .O(N__24142),
            .I(\POWERLED.un1_dutycycle_94_cry_0 ));
    InMux I__4667 (
            .O(N__24139),
            .I(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ));
    CascadeMux I__4666 (
            .O(N__24136),
            .I(\POWERLED.dutycycleZ0Z_13_cascade_ ));
    CascadeMux I__4665 (
            .O(N__24133),
            .I(\POWERLED.N_2293_i_cascade_ ));
    InMux I__4664 (
            .O(N__24130),
            .I(N__24127));
    LocalMux I__4663 (
            .O(N__24127),
            .I(\POWERLED.dutycycle_eena_2 ));
    InMux I__4662 (
            .O(N__24124),
            .I(N__24118));
    InMux I__4661 (
            .O(N__24123),
            .I(N__24118));
    LocalMux I__4660 (
            .O(N__24118),
            .I(\POWERLED.dutycycleZ1Z_9 ));
    CascadeMux I__4659 (
            .O(N__24115),
            .I(\POWERLED.dutycycle_eena_2_cascade_ ));
    CascadeMux I__4658 (
            .O(N__24112),
            .I(\POWERLED.dutycycleZ0Z_2_cascade_ ));
    InMux I__4657 (
            .O(N__24109),
            .I(N__24103));
    InMux I__4656 (
            .O(N__24108),
            .I(N__24103));
    LocalMux I__4655 (
            .O(N__24103),
            .I(\POWERLED.dutycycleZ1Z_13 ));
    CascadeMux I__4654 (
            .O(N__24100),
            .I(N__24096));
    InMux I__4653 (
            .O(N__24099),
            .I(N__24093));
    InMux I__4652 (
            .O(N__24096),
            .I(N__24090));
    LocalMux I__4651 (
            .O(N__24093),
            .I(\POWERLED.un1_dutycycle_53_7_a0_0 ));
    LocalMux I__4650 (
            .O(N__24090),
            .I(\POWERLED.un1_dutycycle_53_7_a0_0 ));
    CascadeMux I__4649 (
            .O(N__24085),
            .I(N__24081));
    InMux I__4648 (
            .O(N__24084),
            .I(N__24078));
    InMux I__4647 (
            .O(N__24081),
            .I(N__24075));
    LocalMux I__4646 (
            .O(N__24078),
            .I(N__24072));
    LocalMux I__4645 (
            .O(N__24075),
            .I(N__24069));
    Span4Mux_s3_v I__4644 (
            .O(N__24072),
            .I(N__24064));
    Span4Mux_h I__4643 (
            .O(N__24069),
            .I(N__24064));
    Odrv4 I__4642 (
            .O(N__24064),
            .I(\POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434 ));
    CascadeMux I__4641 (
            .O(N__24061),
            .I(N__24058));
    InMux I__4640 (
            .O(N__24058),
            .I(N__24055));
    LocalMux I__4639 (
            .O(N__24055),
            .I(\POWERLED.un1_dutycycle_53_i_29 ));
    InMux I__4638 (
            .O(N__24052),
            .I(\POWERLED.mult1_un47_sum_cry_2 ));
    CascadeMux I__4637 (
            .O(N__24049),
            .I(N__24046));
    InMux I__4636 (
            .O(N__24046),
            .I(N__24043));
    LocalMux I__4635 (
            .O(N__24043),
            .I(\POWERLED.mult1_un47_sum_axb_4 ));
    CascadeMux I__4634 (
            .O(N__24040),
            .I(N__24037));
    InMux I__4633 (
            .O(N__24037),
            .I(N__24034));
    LocalMux I__4632 (
            .O(N__24034),
            .I(\POWERLED.mult1_un47_sum_cry_4_s ));
    InMux I__4631 (
            .O(N__24031),
            .I(\POWERLED.mult1_un47_sum_cry_3 ));
    CascadeMux I__4630 (
            .O(N__24028),
            .I(N__24025));
    InMux I__4629 (
            .O(N__24025),
            .I(N__24022));
    LocalMux I__4628 (
            .O(N__24022),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_4 ));
    CascadeMux I__4627 (
            .O(N__24019),
            .I(N__24016));
    InMux I__4626 (
            .O(N__24016),
            .I(N__24013));
    LocalMux I__4625 (
            .O(N__24013),
            .I(\POWERLED.mult1_un47_sum_cry_5_s ));
    InMux I__4624 (
            .O(N__24010),
            .I(\POWERLED.mult1_un47_sum_cry_4 ));
    CascadeMux I__4623 (
            .O(N__24007),
            .I(N__24004));
    InMux I__4622 (
            .O(N__24004),
            .I(N__24001));
    LocalMux I__4621 (
            .O(N__24001),
            .I(N__23998));
    Span4Mux_h I__4620 (
            .O(N__23998),
            .I(N__23995));
    Odrv4 I__4619 (
            .O(N__23995),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_5 ));
    InMux I__4618 (
            .O(N__23992),
            .I(N__23985));
    InMux I__4617 (
            .O(N__23991),
            .I(N__23985));
    InMux I__4616 (
            .O(N__23990),
            .I(N__23982));
    LocalMux I__4615 (
            .O(N__23985),
            .I(\POWERLED.mult1_un47_sum_cry_6_s ));
    LocalMux I__4614 (
            .O(N__23982),
            .I(\POWERLED.mult1_un47_sum_cry_6_s ));
    InMux I__4613 (
            .O(N__23977),
            .I(\POWERLED.mult1_un47_sum_cry_5 ));
    CascadeMux I__4612 (
            .O(N__23974),
            .I(N__23971));
    InMux I__4611 (
            .O(N__23971),
            .I(N__23968));
    LocalMux I__4610 (
            .O(N__23968),
            .I(\POWERLED.mult1_un54_sum_cry_7_THRU_CO ));
    InMux I__4609 (
            .O(N__23965),
            .I(\POWERLED.mult1_un47_sum_cry_6 ));
    InMux I__4608 (
            .O(N__23962),
            .I(N__23959));
    LocalMux I__4607 (
            .O(N__23959),
            .I(N__23956));
    Odrv12 I__4606 (
            .O(N__23956),
            .I(\POWERLED.mult1_un61_sum_i_8 ));
    CascadeMux I__4605 (
            .O(N__23953),
            .I(N__23950));
    InMux I__4604 (
            .O(N__23950),
            .I(N__23945));
    InMux I__4603 (
            .O(N__23949),
            .I(N__23942));
    InMux I__4602 (
            .O(N__23948),
            .I(N__23939));
    LocalMux I__4601 (
            .O(N__23945),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__4600 (
            .O(N__23942),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__4599 (
            .O(N__23939),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    InMux I__4598 (
            .O(N__23932),
            .I(N__23929));
    LocalMux I__4597 (
            .O(N__23929),
            .I(\POWERLED.mult1_un47_sum_l_fx_3 ));
    CascadeMux I__4596 (
            .O(N__23926),
            .I(\POWERLED.mult1_un75_sum_s_8_cascade_ ));
    CascadeMux I__4595 (
            .O(N__23923),
            .I(N__23919));
    CascadeMux I__4594 (
            .O(N__23922),
            .I(N__23915));
    InMux I__4593 (
            .O(N__23919),
            .I(N__23908));
    InMux I__4592 (
            .O(N__23918),
            .I(N__23908));
    InMux I__4591 (
            .O(N__23915),
            .I(N__23908));
    LocalMux I__4590 (
            .O(N__23908),
            .I(\POWERLED.mult1_un75_sum_i_0_8 ));
    InMux I__4589 (
            .O(N__23905),
            .I(N__23901));
    InMux I__4588 (
            .O(N__23904),
            .I(N__23898));
    LocalMux I__4587 (
            .O(N__23901),
            .I(N__23895));
    LocalMux I__4586 (
            .O(N__23898),
            .I(N__23892));
    Span4Mux_v I__4585 (
            .O(N__23895),
            .I(N__23889));
    Odrv12 I__4584 (
            .O(N__23892),
            .I(\POWERLED.mult1_un54_sum ));
    Odrv4 I__4583 (
            .O(N__23889),
            .I(\POWERLED.mult1_un54_sum ));
    CascadeMux I__4582 (
            .O(N__23884),
            .I(N__23881));
    InMux I__4581 (
            .O(N__23881),
            .I(N__23878));
    LocalMux I__4580 (
            .O(N__23878),
            .I(N__23875));
    Odrv4 I__4579 (
            .O(N__23875),
            .I(\POWERLED.un1_dutycycle_53_i_28 ));
    InMux I__4578 (
            .O(N__23872),
            .I(\POWERLED.mult1_un54_sum_cry_2 ));
    InMux I__4577 (
            .O(N__23869),
            .I(\POWERLED.mult1_un54_sum_cry_3 ));
    InMux I__4576 (
            .O(N__23866),
            .I(\POWERLED.mult1_un54_sum_cry_4 ));
    InMux I__4575 (
            .O(N__23863),
            .I(\POWERLED.mult1_un54_sum_cry_5 ));
    InMux I__4574 (
            .O(N__23860),
            .I(\POWERLED.mult1_un54_sum_cry_6 ));
    InMux I__4573 (
            .O(N__23857),
            .I(\POWERLED.mult1_un54_sum_cry_7 ));
    CascadeMux I__4572 (
            .O(N__23854),
            .I(N__23851));
    InMux I__4571 (
            .O(N__23851),
            .I(N__23848));
    LocalMux I__4570 (
            .O(N__23848),
            .I(\POWERLED.mult1_un47_sum_l_fx_6 ));
    InMux I__4569 (
            .O(N__23845),
            .I(N__23842));
    LocalMux I__4568 (
            .O(N__23842),
            .I(N__23838));
    CascadeMux I__4567 (
            .O(N__23841),
            .I(N__23834));
    Span4Mux_h I__4566 (
            .O(N__23838),
            .I(N__23829));
    InMux I__4565 (
            .O(N__23837),
            .I(N__23824));
    InMux I__4564 (
            .O(N__23834),
            .I(N__23824));
    InMux I__4563 (
            .O(N__23833),
            .I(N__23821));
    InMux I__4562 (
            .O(N__23832),
            .I(N__23818));
    Odrv4 I__4561 (
            .O(N__23829),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__4560 (
            .O(N__23824),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__4559 (
            .O(N__23821),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__4558 (
            .O(N__23818),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    InMux I__4557 (
            .O(N__23809),
            .I(N__23805));
    InMux I__4556 (
            .O(N__23808),
            .I(N__23802));
    LocalMux I__4555 (
            .O(N__23805),
            .I(N__23797));
    LocalMux I__4554 (
            .O(N__23802),
            .I(N__23797));
    Span4Mux_h I__4553 (
            .O(N__23797),
            .I(N__23794));
    Odrv4 I__4552 (
            .O(N__23794),
            .I(\POWERLED.mult1_un75_sum ));
    InMux I__4551 (
            .O(N__23791),
            .I(N__23788));
    LocalMux I__4550 (
            .O(N__23788),
            .I(N__23785));
    Span4Mux_s1_v I__4549 (
            .O(N__23785),
            .I(N__23782));
    Odrv4 I__4548 (
            .O(N__23782),
            .I(\POWERLED.mult1_un68_sum_i ));
    CascadeMux I__4547 (
            .O(N__23779),
            .I(N__23776));
    InMux I__4546 (
            .O(N__23776),
            .I(N__23773));
    LocalMux I__4545 (
            .O(N__23773),
            .I(\POWERLED.mult1_un75_sum_cry_3_s ));
    InMux I__4544 (
            .O(N__23770),
            .I(\POWERLED.mult1_un75_sum_cry_2 ));
    InMux I__4543 (
            .O(N__23767),
            .I(N__23764));
    LocalMux I__4542 (
            .O(N__23764),
            .I(\POWERLED.mult1_un75_sum_cry_4_s ));
    InMux I__4541 (
            .O(N__23761),
            .I(\POWERLED.mult1_un75_sum_cry_3 ));
    CascadeMux I__4540 (
            .O(N__23758),
            .I(N__23755));
    InMux I__4539 (
            .O(N__23755),
            .I(N__23752));
    LocalMux I__4538 (
            .O(N__23752),
            .I(\POWERLED.mult1_un75_sum_cry_5_s ));
    InMux I__4537 (
            .O(N__23749),
            .I(\POWERLED.mult1_un75_sum_cry_4 ));
    InMux I__4536 (
            .O(N__23746),
            .I(N__23743));
    LocalMux I__4535 (
            .O(N__23743),
            .I(\POWERLED.mult1_un75_sum_cry_6_s ));
    InMux I__4534 (
            .O(N__23740),
            .I(\POWERLED.mult1_un75_sum_cry_5 ));
    CascadeMux I__4533 (
            .O(N__23737),
            .I(N__23733));
    CascadeMux I__4532 (
            .O(N__23736),
            .I(N__23729));
    InMux I__4531 (
            .O(N__23733),
            .I(N__23722));
    InMux I__4530 (
            .O(N__23732),
            .I(N__23722));
    InMux I__4529 (
            .O(N__23729),
            .I(N__23722));
    LocalMux I__4528 (
            .O(N__23722),
            .I(\POWERLED.mult1_un68_sum_i_0_8 ));
    CascadeMux I__4527 (
            .O(N__23719),
            .I(N__23716));
    InMux I__4526 (
            .O(N__23716),
            .I(N__23713));
    LocalMux I__4525 (
            .O(N__23713),
            .I(\POWERLED.mult1_un82_sum_axb_8 ));
    InMux I__4524 (
            .O(N__23710),
            .I(\POWERLED.mult1_un75_sum_cry_6 ));
    InMux I__4523 (
            .O(N__23707),
            .I(\POWERLED.mult1_un75_sum_cry_7 ));
    InMux I__4522 (
            .O(N__23704),
            .I(N__23700));
    CascadeMux I__4521 (
            .O(N__23703),
            .I(N__23696));
    LocalMux I__4520 (
            .O(N__23700),
            .I(N__23692));
    InMux I__4519 (
            .O(N__23699),
            .I(N__23687));
    InMux I__4518 (
            .O(N__23696),
            .I(N__23687));
    InMux I__4517 (
            .O(N__23695),
            .I(N__23684));
    Odrv4 I__4516 (
            .O(N__23692),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__4515 (
            .O(N__23687),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__4514 (
            .O(N__23684),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    InMux I__4513 (
            .O(N__23677),
            .I(N__23673));
    InMux I__4512 (
            .O(N__23676),
            .I(N__23670));
    LocalMux I__4511 (
            .O(N__23673),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    LocalMux I__4510 (
            .O(N__23670),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    InMux I__4509 (
            .O(N__23665),
            .I(N__23661));
    InMux I__4508 (
            .O(N__23664),
            .I(N__23658));
    LocalMux I__4507 (
            .O(N__23661),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    LocalMux I__4506 (
            .O(N__23658),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    CascadeMux I__4505 (
            .O(N__23653),
            .I(N__23649));
    InMux I__4504 (
            .O(N__23652),
            .I(N__23646));
    InMux I__4503 (
            .O(N__23649),
            .I(N__23643));
    LocalMux I__4502 (
            .O(N__23646),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    LocalMux I__4501 (
            .O(N__23643),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    InMux I__4500 (
            .O(N__23638),
            .I(N__23634));
    InMux I__4499 (
            .O(N__23637),
            .I(N__23631));
    LocalMux I__4498 (
            .O(N__23634),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    LocalMux I__4497 (
            .O(N__23631),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    InMux I__4496 (
            .O(N__23626),
            .I(N__23623));
    LocalMux I__4495 (
            .O(N__23623),
            .I(\VPP_VDDQ.un6_count_8 ));
    IoInMux I__4494 (
            .O(N__23620),
            .I(N__23617));
    LocalMux I__4493 (
            .O(N__23617),
            .I(N__23614));
    Span4Mux_s3_h I__4492 (
            .O(N__23614),
            .I(N__23611));
    Span4Mux_h I__4491 (
            .O(N__23611),
            .I(N__23608));
    Odrv4 I__4490 (
            .O(N__23608),
            .I(v1p8a_en));
    InMux I__4489 (
            .O(N__23605),
            .I(N__23602));
    LocalMux I__4488 (
            .O(N__23602),
            .I(N__23598));
    InMux I__4487 (
            .O(N__23601),
            .I(N__23595));
    Span4Mux_s1_v I__4486 (
            .O(N__23598),
            .I(N__23592));
    LocalMux I__4485 (
            .O(N__23595),
            .I(N__23589));
    Span4Mux_v I__4484 (
            .O(N__23592),
            .I(N__23586));
    Odrv12 I__4483 (
            .O(N__23589),
            .I(\POWERLED.mult1_un82_sum ));
    Odrv4 I__4482 (
            .O(N__23586),
            .I(\POWERLED.mult1_un82_sum ));
    InMux I__4481 (
            .O(N__23581),
            .I(N__23578));
    LocalMux I__4480 (
            .O(N__23578),
            .I(N__23575));
    Span4Mux_s1_v I__4479 (
            .O(N__23575),
            .I(N__23572));
    Odrv4 I__4478 (
            .O(N__23572),
            .I(\POWERLED.mult1_un75_sum_i ));
    CascadeMux I__4477 (
            .O(N__23569),
            .I(N__23566));
    InMux I__4476 (
            .O(N__23566),
            .I(N__23563));
    LocalMux I__4475 (
            .O(N__23563),
            .I(\POWERLED.mult1_un82_sum_cry_3_s ));
    InMux I__4474 (
            .O(N__23560),
            .I(\POWERLED.mult1_un82_sum_cry_2_c ));
    InMux I__4473 (
            .O(N__23557),
            .I(N__23554));
    LocalMux I__4472 (
            .O(N__23554),
            .I(\POWERLED.mult1_un82_sum_cry_4_s ));
    InMux I__4471 (
            .O(N__23551),
            .I(\POWERLED.mult1_un82_sum_cry_3_c ));
    CascadeMux I__4470 (
            .O(N__23548),
            .I(N__23545));
    InMux I__4469 (
            .O(N__23545),
            .I(N__23542));
    LocalMux I__4468 (
            .O(N__23542),
            .I(\POWERLED.mult1_un82_sum_cry_5_s ));
    InMux I__4467 (
            .O(N__23539),
            .I(\POWERLED.mult1_un82_sum_cry_4_c ));
    InMux I__4466 (
            .O(N__23536),
            .I(N__23533));
    LocalMux I__4465 (
            .O(N__23533),
            .I(\POWERLED.mult1_un82_sum_cry_6_s ));
    InMux I__4464 (
            .O(N__23530),
            .I(\POWERLED.mult1_un82_sum_cry_5_c ));
    CascadeMux I__4463 (
            .O(N__23527),
            .I(N__23524));
    InMux I__4462 (
            .O(N__23524),
            .I(N__23521));
    LocalMux I__4461 (
            .O(N__23521),
            .I(\POWERLED.mult1_un89_sum_axb_8 ));
    InMux I__4460 (
            .O(N__23518),
            .I(\POWERLED.mult1_un82_sum_cry_6_c ));
    InMux I__4459 (
            .O(N__23515),
            .I(\POWERLED.mult1_un82_sum_cry_7 ));
    InMux I__4458 (
            .O(N__23512),
            .I(N__23508));
    InMux I__4457 (
            .O(N__23511),
            .I(N__23505));
    LocalMux I__4456 (
            .O(N__23508),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    LocalMux I__4455 (
            .O(N__23505),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    InMux I__4454 (
            .O(N__23500),
            .I(N__23496));
    InMux I__4453 (
            .O(N__23499),
            .I(N__23493));
    LocalMux I__4452 (
            .O(N__23496),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    LocalMux I__4451 (
            .O(N__23493),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    CascadeMux I__4450 (
            .O(N__23488),
            .I(N__23484));
    InMux I__4449 (
            .O(N__23487),
            .I(N__23481));
    InMux I__4448 (
            .O(N__23484),
            .I(N__23478));
    LocalMux I__4447 (
            .O(N__23481),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    LocalMux I__4446 (
            .O(N__23478),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    InMux I__4445 (
            .O(N__23473),
            .I(N__23469));
    InMux I__4444 (
            .O(N__23472),
            .I(N__23466));
    LocalMux I__4443 (
            .O(N__23469),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    LocalMux I__4442 (
            .O(N__23466),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    InMux I__4441 (
            .O(N__23461),
            .I(N__23447));
    InMux I__4440 (
            .O(N__23460),
            .I(N__23447));
    InMux I__4439 (
            .O(N__23459),
            .I(N__23447));
    InMux I__4438 (
            .O(N__23458),
            .I(N__23447));
    InMux I__4437 (
            .O(N__23457),
            .I(N__23442));
    InMux I__4436 (
            .O(N__23456),
            .I(N__23442));
    LocalMux I__4435 (
            .O(N__23447),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    LocalMux I__4434 (
            .O(N__23442),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    InMux I__4433 (
            .O(N__23437),
            .I(N__23434));
    LocalMux I__4432 (
            .O(N__23434),
            .I(N_325));
    InMux I__4431 (
            .O(N__23431),
            .I(N__23425));
    InMux I__4430 (
            .O(N__23430),
            .I(N__23425));
    LocalMux I__4429 (
            .O(N__23425),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    InMux I__4428 (
            .O(N__23422),
            .I(N__23412));
    InMux I__4427 (
            .O(N__23421),
            .I(N__23412));
    InMux I__4426 (
            .O(N__23420),
            .I(N__23403));
    InMux I__4425 (
            .O(N__23419),
            .I(N__23403));
    InMux I__4424 (
            .O(N__23418),
            .I(N__23403));
    InMux I__4423 (
            .O(N__23417),
            .I(N__23403));
    LocalMux I__4422 (
            .O(N__23412),
            .I(VPP_VDDQ_curr_state_0));
    LocalMux I__4421 (
            .O(N__23403),
            .I(VPP_VDDQ_curr_state_0));
    CascadeMux I__4420 (
            .O(N__23398),
            .I(N_325_cascade_));
    CascadeMux I__4419 (
            .O(N__23395),
            .I(N__23392));
    InMux I__4418 (
            .O(N__23392),
            .I(N__23389));
    LocalMux I__4417 (
            .O(N__23389),
            .I(\VPP_VDDQ.delayed_vddq_pwrgd_0 ));
    InMux I__4416 (
            .O(N__23386),
            .I(N__23381));
    InMux I__4415 (
            .O(N__23385),
            .I(N__23378));
    InMux I__4414 (
            .O(N__23384),
            .I(N__23375));
    LocalMux I__4413 (
            .O(N__23381),
            .I(N__23371));
    LocalMux I__4412 (
            .O(N__23378),
            .I(N__23365));
    LocalMux I__4411 (
            .O(N__23375),
            .I(N__23362));
    InMux I__4410 (
            .O(N__23374),
            .I(N__23359));
    Span4Mux_h I__4409 (
            .O(N__23371),
            .I(N__23356));
    InMux I__4408 (
            .O(N__23370),
            .I(N__23353));
    InMux I__4407 (
            .O(N__23369),
            .I(N__23348));
    InMux I__4406 (
            .O(N__23368),
            .I(N__23348));
    Span4Mux_h I__4405 (
            .O(N__23365),
            .I(N__23345));
    Span4Mux_v I__4404 (
            .O(N__23362),
            .I(N__23340));
    LocalMux I__4403 (
            .O(N__23359),
            .I(N__23340));
    Span4Mux_v I__4402 (
            .O(N__23356),
            .I(N__23335));
    LocalMux I__4401 (
            .O(N__23353),
            .I(N__23332));
    LocalMux I__4400 (
            .O(N__23348),
            .I(N__23325));
    Span4Mux_v I__4399 (
            .O(N__23345),
            .I(N__23325));
    Span4Mux_h I__4398 (
            .O(N__23340),
            .I(N__23325));
    InMux I__4397 (
            .O(N__23339),
            .I(N__23322));
    InMux I__4396 (
            .O(N__23338),
            .I(N__23319));
    Odrv4 I__4395 (
            .O(N__23335),
            .I(VCCST_EN_i_0));
    Odrv4 I__4394 (
            .O(N__23332),
            .I(VCCST_EN_i_0));
    Odrv4 I__4393 (
            .O(N__23325),
            .I(VCCST_EN_i_0));
    LocalMux I__4392 (
            .O(N__23322),
            .I(VCCST_EN_i_0));
    LocalMux I__4391 (
            .O(N__23319),
            .I(VCCST_EN_i_0));
    InMux I__4390 (
            .O(N__23308),
            .I(N__23297));
    InMux I__4389 (
            .O(N__23307),
            .I(N__23297));
    InMux I__4388 (
            .O(N__23306),
            .I(N__23297));
    InMux I__4387 (
            .O(N__23305),
            .I(N__23292));
    InMux I__4386 (
            .O(N__23304),
            .I(N__23292));
    LocalMux I__4385 (
            .O(N__23297),
            .I(N__23289));
    LocalMux I__4384 (
            .O(N__23292),
            .I(\VPP_VDDQ.N_541 ));
    Odrv4 I__4383 (
            .O(N__23289),
            .I(\VPP_VDDQ.N_541 ));
    InMux I__4382 (
            .O(N__23284),
            .I(N__23280));
    InMux I__4381 (
            .O(N__23283),
            .I(N__23277));
    LocalMux I__4380 (
            .O(N__23280),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    LocalMux I__4379 (
            .O(N__23277),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    InMux I__4378 (
            .O(N__23272),
            .I(N__23268));
    InMux I__4377 (
            .O(N__23271),
            .I(N__23265));
    LocalMux I__4376 (
            .O(N__23268),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    LocalMux I__4375 (
            .O(N__23265),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    CascadeMux I__4374 (
            .O(N__23260),
            .I(N__23256));
    InMux I__4373 (
            .O(N__23259),
            .I(N__23253));
    InMux I__4372 (
            .O(N__23256),
            .I(N__23250));
    LocalMux I__4371 (
            .O(N__23253),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    LocalMux I__4370 (
            .O(N__23250),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    InMux I__4369 (
            .O(N__23245),
            .I(N__23241));
    InMux I__4368 (
            .O(N__23244),
            .I(N__23238));
    LocalMux I__4367 (
            .O(N__23241),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    LocalMux I__4366 (
            .O(N__23238),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    InMux I__4365 (
            .O(N__23233),
            .I(N__23230));
    LocalMux I__4364 (
            .O(N__23230),
            .I(N__23227));
    Odrv4 I__4363 (
            .O(N__23227),
            .I(\VPP_VDDQ.un6_count_10 ));
    CascadeMux I__4362 (
            .O(N__23224),
            .I(\VPP_VDDQ.un6_count_9_cascade_ ));
    CascadeMux I__4361 (
            .O(N__23221),
            .I(N__23218));
    InMux I__4360 (
            .O(N__23218),
            .I(N__23212));
    InMux I__4359 (
            .O(N__23217),
            .I(N__23212));
    LocalMux I__4358 (
            .O(N__23212),
            .I(N__23209));
    Odrv4 I__4357 (
            .O(N__23209),
            .I(\VPP_VDDQ.un6_count ));
    InMux I__4356 (
            .O(N__23206),
            .I(N__23202));
    InMux I__4355 (
            .O(N__23205),
            .I(N__23199));
    LocalMux I__4354 (
            .O(N__23202),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    LocalMux I__4353 (
            .O(N__23199),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    InMux I__4352 (
            .O(N__23194),
            .I(N__23190));
    InMux I__4351 (
            .O(N__23193),
            .I(N__23187));
    LocalMux I__4350 (
            .O(N__23190),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    LocalMux I__4349 (
            .O(N__23187),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    CascadeMux I__4348 (
            .O(N__23182),
            .I(N__23178));
    InMux I__4347 (
            .O(N__23181),
            .I(N__23175));
    InMux I__4346 (
            .O(N__23178),
            .I(N__23172));
    LocalMux I__4345 (
            .O(N__23175),
            .I(N__23167));
    LocalMux I__4344 (
            .O(N__23172),
            .I(N__23167));
    Odrv4 I__4343 (
            .O(N__23167),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    InMux I__4342 (
            .O(N__23164),
            .I(N__23160));
    InMux I__4341 (
            .O(N__23163),
            .I(N__23157));
    LocalMux I__4340 (
            .O(N__23160),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    LocalMux I__4339 (
            .O(N__23157),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    InMux I__4338 (
            .O(N__23152),
            .I(N__23149));
    LocalMux I__4337 (
            .O(N__23149),
            .I(\VPP_VDDQ.un6_count_11 ));
    CascadeMux I__4336 (
            .O(N__23146),
            .I(\VPP_VDDQ.count_2Z0Z_2_cascade_ ));
    CascadeMux I__4335 (
            .O(N__23143),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_ ));
    InMux I__4334 (
            .O(N__23140),
            .I(N__23137));
    LocalMux I__4333 (
            .O(N__23137),
            .I(\VPP_VDDQ.count_2_0_15 ));
    InMux I__4332 (
            .O(N__23134),
            .I(N__23131));
    LocalMux I__4331 (
            .O(N__23131),
            .I(\VPP_VDDQ.N_551 ));
    IoInMux I__4330 (
            .O(N__23128),
            .I(N__23125));
    LocalMux I__4329 (
            .O(N__23125),
            .I(N__23122));
    IoSpan4Mux I__4328 (
            .O(N__23122),
            .I(N__23119));
    Span4Mux_s1_h I__4327 (
            .O(N__23119),
            .I(N__23116));
    Odrv4 I__4326 (
            .O(N__23116),
            .I(vpp_en));
    CascadeMux I__4325 (
            .O(N__23113),
            .I(\VPP_VDDQ.count_2_1_14_cascade_ ));
    InMux I__4324 (
            .O(N__23110),
            .I(N__23107));
    LocalMux I__4323 (
            .O(N__23107),
            .I(\VPP_VDDQ.count_2_0_4 ));
    InMux I__4322 (
            .O(N__23104),
            .I(N__23101));
    LocalMux I__4321 (
            .O(N__23101),
            .I(\VPP_VDDQ.count_2_0_5 ));
    CascadeMux I__4320 (
            .O(N__23098),
            .I(\VPP_VDDQ.count_2_1_5_cascade_ ));
    CascadeMux I__4319 (
            .O(N__23095),
            .I(N__23092));
    InMux I__4318 (
            .O(N__23092),
            .I(N__23089));
    LocalMux I__4317 (
            .O(N__23089),
            .I(N__23086));
    Span12Mux_s5_v I__4316 (
            .O(N__23086),
            .I(N__23083));
    Odrv12 I__4315 (
            .O(N__23083),
            .I(\VPP_VDDQ.count_2_0_8 ));
    InMux I__4314 (
            .O(N__23080),
            .I(N__23077));
    LocalMux I__4313 (
            .O(N__23077),
            .I(N__23074));
    Span12Mux_s6_v I__4312 (
            .O(N__23074),
            .I(N__23071));
    Odrv12 I__4311 (
            .O(N__23071),
            .I(\VPP_VDDQ.count_2_1_8 ));
    InMux I__4310 (
            .O(N__23068),
            .I(N__23065));
    LocalMux I__4309 (
            .O(N__23065),
            .I(\VPP_VDDQ.count_2_0_2 ));
    CascadeMux I__4308 (
            .O(N__23062),
            .I(\VPP_VDDQ.count_2_1_2_cascade_ ));
    InMux I__4307 (
            .O(N__23059),
            .I(N__23052));
    InMux I__4306 (
            .O(N__23058),
            .I(N__23052));
    InMux I__4305 (
            .O(N__23057),
            .I(N__23049));
    LocalMux I__4304 (
            .O(N__23052),
            .I(N__23046));
    LocalMux I__4303 (
            .O(N__23049),
            .I(\POWERLED.func_state_RNI_0Z0Z_0 ));
    Odrv4 I__4302 (
            .O(N__23046),
            .I(\POWERLED.func_state_RNI_0Z0Z_0 ));
    CascadeMux I__4301 (
            .O(N__23041),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_5_cascade_ ));
    InMux I__4300 (
            .O(N__23038),
            .I(N__23035));
    LocalMux I__4299 (
            .O(N__23035),
            .I(N__23032));
    Span4Mux_h I__4298 (
            .O(N__23032),
            .I(N__23028));
    InMux I__4297 (
            .O(N__23031),
            .I(N__23025));
    Odrv4 I__4296 (
            .O(N__23028),
            .I(\POWERLED.func_state_RNI_5Z0Z_0 ));
    LocalMux I__4295 (
            .O(N__23025),
            .I(\POWERLED.func_state_RNI_5Z0Z_0 ));
    InMux I__4294 (
            .O(N__23020),
            .I(N__23012));
    InMux I__4293 (
            .O(N__23019),
            .I(N__23005));
    InMux I__4292 (
            .O(N__23018),
            .I(N__23005));
    InMux I__4291 (
            .O(N__23017),
            .I(N__23005));
    InMux I__4290 (
            .O(N__23016),
            .I(N__23000));
    InMux I__4289 (
            .O(N__23015),
            .I(N__23000));
    LocalMux I__4288 (
            .O(N__23012),
            .I(SUSWARN_N_rep1));
    LocalMux I__4287 (
            .O(N__23005),
            .I(SUSWARN_N_rep1));
    LocalMux I__4286 (
            .O(N__23000),
            .I(SUSWARN_N_rep1));
    CascadeMux I__4285 (
            .O(N__22993),
            .I(\POWERLED.dutycycle_eena_5_0_s_tzZ0Z_1_cascade_ ));
    CascadeMux I__4284 (
            .O(N__22990),
            .I(N__22984));
    InMux I__4283 (
            .O(N__22989),
            .I(N__22980));
    CascadeMux I__4282 (
            .O(N__22988),
            .I(N__22977));
    CascadeMux I__4281 (
            .O(N__22987),
            .I(N__22974));
    InMux I__4280 (
            .O(N__22984),
            .I(N__22969));
    InMux I__4279 (
            .O(N__22983),
            .I(N__22969));
    LocalMux I__4278 (
            .O(N__22980),
            .I(N__22966));
    InMux I__4277 (
            .O(N__22977),
            .I(N__22961));
    InMux I__4276 (
            .O(N__22974),
            .I(N__22961));
    LocalMux I__4275 (
            .O(N__22969),
            .I(N__22957));
    Span4Mux_v I__4274 (
            .O(N__22966),
            .I(N__22952));
    LocalMux I__4273 (
            .O(N__22961),
            .I(N__22952));
    InMux I__4272 (
            .O(N__22960),
            .I(N__22949));
    Span4Mux_v I__4271 (
            .O(N__22957),
            .I(N__22944));
    Span4Mux_h I__4270 (
            .O(N__22952),
            .I(N__22944));
    LocalMux I__4269 (
            .O(N__22949),
            .I(\POWERLED.N_443 ));
    Odrv4 I__4268 (
            .O(N__22944),
            .I(\POWERLED.N_443 ));
    CascadeMux I__4267 (
            .O(N__22939),
            .I(POWERLED_func_state_0_sqmuxa_cascade_));
    CascadeMux I__4266 (
            .O(N__22936),
            .I(N__22933));
    InMux I__4265 (
            .O(N__22933),
            .I(N__22930));
    LocalMux I__4264 (
            .O(N__22930),
            .I(N__22927));
    Odrv4 I__4263 (
            .O(N__22927),
            .I(N_14));
    CascadeMux I__4262 (
            .O(N__22924),
            .I(\VPP_VDDQ.count_2_1_4_cascade_ ));
    InMux I__4261 (
            .O(N__22921),
            .I(N__22918));
    LocalMux I__4260 (
            .O(N__22918),
            .I(\POWERLED.dutycycle_RNI9NTJ2Z0Z_2 ));
    CascadeMux I__4259 (
            .O(N__22915),
            .I(\POWERLED.dutycycle_RNI9NTJ2Z0Z_2_cascade_ ));
    InMux I__4258 (
            .O(N__22912),
            .I(N__22906));
    InMux I__4257 (
            .O(N__22911),
            .I(N__22906));
    LocalMux I__4256 (
            .O(N__22906),
            .I(\POWERLED.dutycycleZ1Z_2 ));
    CascadeMux I__4255 (
            .O(N__22903),
            .I(N_2145_i_cascade_));
    CascadeMux I__4254 (
            .O(N__22900),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_6_cascade_ ));
    CascadeMux I__4253 (
            .O(N__22897),
            .I(N__22890));
    CascadeMux I__4252 (
            .O(N__22896),
            .I(N__22886));
    InMux I__4251 (
            .O(N__22895),
            .I(N__22880));
    InMux I__4250 (
            .O(N__22894),
            .I(N__22880));
    InMux I__4249 (
            .O(N__22893),
            .I(N__22875));
    InMux I__4248 (
            .O(N__22890),
            .I(N__22875));
    InMux I__4247 (
            .O(N__22889),
            .I(N__22871));
    InMux I__4246 (
            .O(N__22886),
            .I(N__22866));
    InMux I__4245 (
            .O(N__22885),
            .I(N__22866));
    LocalMux I__4244 (
            .O(N__22880),
            .I(N__22863));
    LocalMux I__4243 (
            .O(N__22875),
            .I(N__22858));
    CascadeMux I__4242 (
            .O(N__22874),
            .I(N__22854));
    LocalMux I__4241 (
            .O(N__22871),
            .I(N__22849));
    LocalMux I__4240 (
            .O(N__22866),
            .I(N__22849));
    Span4Mux_h I__4239 (
            .O(N__22863),
            .I(N__22846));
    InMux I__4238 (
            .O(N__22862),
            .I(N__22841));
    InMux I__4237 (
            .O(N__22861),
            .I(N__22841));
    Span4Mux_h I__4236 (
            .O(N__22858),
            .I(N__22838));
    InMux I__4235 (
            .O(N__22857),
            .I(N__22833));
    InMux I__4234 (
            .O(N__22854),
            .I(N__22833));
    Odrv12 I__4233 (
            .O(N__22849),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv4 I__4232 (
            .O(N__22846),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__4231 (
            .O(N__22841),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv4 I__4230 (
            .O(N__22838),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__4229 (
            .O(N__22833),
            .I(\POWERLED.func_stateZ0Z_0 ));
    InMux I__4228 (
            .O(N__22822),
            .I(N__22819));
    LocalMux I__4227 (
            .O(N__22819),
            .I(\RSMRST_PWRGD.N_13 ));
    InMux I__4226 (
            .O(N__22816),
            .I(N__22813));
    LocalMux I__4225 (
            .O(N__22813),
            .I(POWERLED_dutycycle_eena_14_0));
    InMux I__4224 (
            .O(N__22810),
            .I(N__22806));
    InMux I__4223 (
            .O(N__22809),
            .I(N__22803));
    LocalMux I__4222 (
            .O(N__22806),
            .I(\POWERLED.dutycycle_0_5 ));
    LocalMux I__4221 (
            .O(N__22803),
            .I(\POWERLED.dutycycle_0_5 ));
    CascadeMux I__4220 (
            .O(N__22798),
            .I(POWERLED_dutycycle_eena_14_0_cascade_));
    CascadeMux I__4219 (
            .O(N__22795),
            .I(dutycycle_RNIKBMSJ_0_5_cascade_));
    InMux I__4218 (
            .O(N__22792),
            .I(N__22789));
    LocalMux I__4217 (
            .O(N__22789),
            .I(\POWERLED.dutycycle_eena ));
    CascadeMux I__4216 (
            .O(N__22786),
            .I(\POWERLED.dutycycle_eena_cascade_ ));
    InMux I__4215 (
            .O(N__22783),
            .I(N__22780));
    LocalMux I__4214 (
            .O(N__22780),
            .I(\POWERLED.N_81 ));
    InMux I__4213 (
            .O(N__22777),
            .I(N__22773));
    InMux I__4212 (
            .O(N__22776),
            .I(N__22770));
    LocalMux I__4211 (
            .O(N__22773),
            .I(\POWERLED.dutycycleZ1Z_0 ));
    LocalMux I__4210 (
            .O(N__22770),
            .I(\POWERLED.dutycycleZ1Z_0 ));
    CascadeMux I__4209 (
            .O(N__22765),
            .I(\POWERLED.N_441_cascade_ ));
    InMux I__4208 (
            .O(N__22762),
            .I(N__22759));
    LocalMux I__4207 (
            .O(N__22759),
            .I(N__22756));
    Sp12to4 I__4206 (
            .O(N__22756),
            .I(N__22753));
    Odrv12 I__4205 (
            .O(N__22753),
            .I(\POWERLED.dutycycle_eena_13 ));
    InMux I__4204 (
            .O(N__22750),
            .I(N__22747));
    LocalMux I__4203 (
            .O(N__22747),
            .I(N__22743));
    InMux I__4202 (
            .O(N__22746),
            .I(N__22740));
    Span4Mux_v I__4201 (
            .O(N__22743),
            .I(N__22737));
    LocalMux I__4200 (
            .O(N__22740),
            .I(\POWERLED.dutycycle_0_6 ));
    Odrv4 I__4199 (
            .O(N__22737),
            .I(\POWERLED.dutycycle_0_6 ));
    CascadeMux I__4198 (
            .O(N__22732),
            .I(\POWERLED.dutycycle_eena_13_cascade_ ));
    CascadeMux I__4197 (
            .O(N__22729),
            .I(\POWERLED.dutycycleZ1Z_6_cascade_ ));
    InMux I__4196 (
            .O(N__22726),
            .I(N__22723));
    LocalMux I__4195 (
            .O(N__22723),
            .I(\POWERLED.N_442 ));
    CascadeMux I__4194 (
            .O(N__22720),
            .I(\POWERLED.N_429_cascade_ ));
    InMux I__4193 (
            .O(N__22717),
            .I(N__22714));
    LocalMux I__4192 (
            .O(N__22714),
            .I(\POWERLED.dutycycle_RNI_8Z0Z_10 ));
    InMux I__4191 (
            .O(N__22711),
            .I(N__22705));
    InMux I__4190 (
            .O(N__22710),
            .I(N__22705));
    LocalMux I__4189 (
            .O(N__22705),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    CascadeMux I__4188 (
            .O(N__22702),
            .I(\POWERLED.dutycycleZ0Z_12_cascade_ ));
    InMux I__4187 (
            .O(N__22699),
            .I(N__22696));
    LocalMux I__4186 (
            .O(N__22696),
            .I(\POWERLED.dutycycle_RNIZ0Z_15 ));
    InMux I__4185 (
            .O(N__22693),
            .I(N__22690));
    LocalMux I__4184 (
            .O(N__22690),
            .I(N__22687));
    Odrv4 I__4183 (
            .O(N__22687),
            .I(\POWERLED.m69_0_o2_7 ));
    CascadeMux I__4182 (
            .O(N__22684),
            .I(\POWERLED.N_81_cascade_ ));
    InMux I__4181 (
            .O(N__22681),
            .I(N__22678));
    LocalMux I__4180 (
            .O(N__22678),
            .I(\POWERLED.N_85 ));
    InMux I__4179 (
            .O(N__22675),
            .I(N__22671));
    InMux I__4178 (
            .O(N__22674),
            .I(N__22668));
    LocalMux I__4177 (
            .O(N__22671),
            .I(\POWERLED.dutycycleZ1Z_1 ));
    LocalMux I__4176 (
            .O(N__22668),
            .I(\POWERLED.dutycycleZ1Z_1 ));
    CascadeMux I__4175 (
            .O(N__22663),
            .I(\POWERLED.N_85_cascade_ ));
    CascadeMux I__4174 (
            .O(N__22660),
            .I(\POWERLED.dutycycle_cascade_ ));
    InMux I__4173 (
            .O(N__22657),
            .I(N__22651));
    InMux I__4172 (
            .O(N__22656),
            .I(N__22651));
    LocalMux I__4171 (
            .O(N__22651),
            .I(\POWERLED.dutycycle_eena_0 ));
    CascadeMux I__4170 (
            .O(N__22648),
            .I(\POWERLED.N_9_i_1_cascade_ ));
    InMux I__4169 (
            .O(N__22645),
            .I(N__22642));
    LocalMux I__4168 (
            .O(N__22642),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_7 ));
    CascadeMux I__4167 (
            .O(N__22639),
            .I(N__22636));
    InMux I__4166 (
            .O(N__22636),
            .I(N__22632));
    InMux I__4165 (
            .O(N__22635),
            .I(N__22629));
    LocalMux I__4164 (
            .O(N__22632),
            .I(\POWERLED.dutycycleZ1Z_4 ));
    LocalMux I__4163 (
            .O(N__22629),
            .I(\POWERLED.dutycycleZ1Z_4 ));
    InMux I__4162 (
            .O(N__22624),
            .I(N__22620));
    InMux I__4161 (
            .O(N__22623),
            .I(N__22617));
    LocalMux I__4160 (
            .O(N__22620),
            .I(\POWERLED.dutycycle_en_6 ));
    LocalMux I__4159 (
            .O(N__22617),
            .I(\POWERLED.dutycycle_en_6 ));
    CascadeMux I__4158 (
            .O(N__22612),
            .I(\POWERLED.dutycycleZ0Z_8_cascade_ ));
    CascadeMux I__4157 (
            .O(N__22609),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_4_cascade_ ));
    CascadeMux I__4156 (
            .O(N__22606),
            .I(\POWERLED.un1_dutycycle_53_axb_12_cascade_ ));
    CascadeMux I__4155 (
            .O(N__22603),
            .I(N__22600));
    InMux I__4154 (
            .O(N__22600),
            .I(N__22597));
    LocalMux I__4153 (
            .O(N__22597),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_15 ));
    InMux I__4152 (
            .O(N__22594),
            .I(N__22591));
    LocalMux I__4151 (
            .O(N__22591),
            .I(N__22588));
    Odrv4 I__4150 (
            .O(N__22588),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_1 ));
    CascadeMux I__4149 (
            .O(N__22585),
            .I(\POWERLED.g0_1_1_cascade_ ));
    CascadeMux I__4148 (
            .O(N__22582),
            .I(N__22579));
    InMux I__4147 (
            .O(N__22579),
            .I(N__22576));
    LocalMux I__4146 (
            .O(N__22576),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_3 ));
    CascadeMux I__4145 (
            .O(N__22573),
            .I(N__22570));
    InMux I__4144 (
            .O(N__22570),
            .I(N__22567));
    LocalMux I__4143 (
            .O(N__22567),
            .I(\POWERLED.g0_1_1 ));
    CascadeMux I__4142 (
            .O(N__22564),
            .I(\POWERLED.dutycycle_RNIZ0Z_7_cascade_ ));
    InMux I__4141 (
            .O(N__22561),
            .I(N__22558));
    LocalMux I__4140 (
            .O(N__22558),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_7 ));
    CascadeMux I__4139 (
            .O(N__22555),
            .I(\POWERLED.dutycycle_RNI_9Z0Z_7_cascade_ ));
    CascadeMux I__4138 (
            .O(N__22552),
            .I(N__22549));
    InMux I__4137 (
            .O(N__22549),
            .I(N__22546));
    LocalMux I__4136 (
            .O(N__22546),
            .I(\POWERLED.dutycycle_RNIZ0Z_11 ));
    InMux I__4135 (
            .O(N__22543),
            .I(N__22540));
    LocalMux I__4134 (
            .O(N__22540),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_13 ));
    CascadeMux I__4133 (
            .O(N__22537),
            .I(N__22534));
    InMux I__4132 (
            .O(N__22534),
            .I(N__22531));
    LocalMux I__4131 (
            .O(N__22531),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_12 ));
    InMux I__4130 (
            .O(N__22528),
            .I(N__22525));
    LocalMux I__4129 (
            .O(N__22525),
            .I(\POWERLED.mult1_un96_sum_cry_6_s ));
    CascadeMux I__4128 (
            .O(N__22522),
            .I(N__22519));
    InMux I__4127 (
            .O(N__22519),
            .I(N__22516));
    LocalMux I__4126 (
            .O(N__22516),
            .I(\POWERLED.mult1_un110_sum_axb_8 ));
    InMux I__4125 (
            .O(N__22513),
            .I(\POWERLED.mult1_un103_sum_cry_6 ));
    CascadeMux I__4124 (
            .O(N__22510),
            .I(N__22507));
    InMux I__4123 (
            .O(N__22507),
            .I(N__22504));
    LocalMux I__4122 (
            .O(N__22504),
            .I(\POWERLED.mult1_un103_sum_axb_8 ));
    InMux I__4121 (
            .O(N__22501),
            .I(\POWERLED.mult1_un103_sum_cry_7 ));
    CascadeMux I__4120 (
            .O(N__22498),
            .I(N__22494));
    InMux I__4119 (
            .O(N__22497),
            .I(N__22486));
    InMux I__4118 (
            .O(N__22494),
            .I(N__22486));
    InMux I__4117 (
            .O(N__22493),
            .I(N__22483));
    InMux I__4116 (
            .O(N__22492),
            .I(N__22478));
    InMux I__4115 (
            .O(N__22491),
            .I(N__22478));
    LocalMux I__4114 (
            .O(N__22486),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__4113 (
            .O(N__22483),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__4112 (
            .O(N__22478),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    CascadeMux I__4111 (
            .O(N__22471),
            .I(N__22466));
    InMux I__4110 (
            .O(N__22470),
            .I(N__22461));
    InMux I__4109 (
            .O(N__22469),
            .I(N__22458));
    InMux I__4108 (
            .O(N__22466),
            .I(N__22451));
    InMux I__4107 (
            .O(N__22465),
            .I(N__22451));
    InMux I__4106 (
            .O(N__22464),
            .I(N__22451));
    LocalMux I__4105 (
            .O(N__22461),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__4104 (
            .O(N__22458),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__4103 (
            .O(N__22451),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    CascadeMux I__4102 (
            .O(N__22444),
            .I(N__22440));
    CascadeMux I__4101 (
            .O(N__22443),
            .I(N__22436));
    InMux I__4100 (
            .O(N__22440),
            .I(N__22429));
    InMux I__4099 (
            .O(N__22439),
            .I(N__22429));
    InMux I__4098 (
            .O(N__22436),
            .I(N__22429));
    LocalMux I__4097 (
            .O(N__22429),
            .I(\POWERLED.mult1_un96_sum_i_0_8 ));
    CascadeMux I__4096 (
            .O(N__22426),
            .I(N__22422));
    InMux I__4095 (
            .O(N__22425),
            .I(N__22417));
    InMux I__4094 (
            .O(N__22422),
            .I(N__22410));
    InMux I__4093 (
            .O(N__22421),
            .I(N__22410));
    InMux I__4092 (
            .O(N__22420),
            .I(N__22410));
    LocalMux I__4091 (
            .O(N__22417),
            .I(N__22407));
    LocalMux I__4090 (
            .O(N__22410),
            .I(N__22404));
    Span4Mux_v I__4089 (
            .O(N__22407),
            .I(N__22401));
    Span4Mux_h I__4088 (
            .O(N__22404),
            .I(N__22398));
    Odrv4 I__4087 (
            .O(N__22401),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    Odrv4 I__4086 (
            .O(N__22398),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    CascadeMux I__4085 (
            .O(N__22393),
            .I(N__22390));
    InMux I__4084 (
            .O(N__22390),
            .I(N__22387));
    LocalMux I__4083 (
            .O(N__22387),
            .I(N__22384));
    Span4Mux_v I__4082 (
            .O(N__22384),
            .I(N__22377));
    InMux I__4081 (
            .O(N__22383),
            .I(N__22372));
    InMux I__4080 (
            .O(N__22382),
            .I(N__22372));
    InMux I__4079 (
            .O(N__22381),
            .I(N__22367));
    InMux I__4078 (
            .O(N__22380),
            .I(N__22367));
    Odrv4 I__4077 (
            .O(N__22377),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    LocalMux I__4076 (
            .O(N__22372),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    LocalMux I__4075 (
            .O(N__22367),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    InMux I__4074 (
            .O(N__22360),
            .I(N__22357));
    LocalMux I__4073 (
            .O(N__22357),
            .I(N__22354));
    Span4Mux_h I__4072 (
            .O(N__22354),
            .I(N__22348));
    InMux I__4071 (
            .O(N__22353),
            .I(N__22345));
    InMux I__4070 (
            .O(N__22352),
            .I(N__22340));
    InMux I__4069 (
            .O(N__22351),
            .I(N__22340));
    Odrv4 I__4068 (
            .O(N__22348),
            .I(\POWERLED.count_RNIZ0Z_8 ));
    LocalMux I__4067 (
            .O(N__22345),
            .I(\POWERLED.count_RNIZ0Z_8 ));
    LocalMux I__4066 (
            .O(N__22340),
            .I(\POWERLED.count_RNIZ0Z_8 ));
    InMux I__4065 (
            .O(N__22333),
            .I(N__22330));
    LocalMux I__4064 (
            .O(N__22330),
            .I(N__22327));
    Span4Mux_h I__4063 (
            .O(N__22327),
            .I(N__22324));
    Odrv4 I__4062 (
            .O(N__22324),
            .I(\POWERLED.curr_state_2_0 ));
    CascadeMux I__4061 (
            .O(N__22321),
            .I(N__22317));
    CascadeMux I__4060 (
            .O(N__22320),
            .I(N__22314));
    InMux I__4059 (
            .O(N__22317),
            .I(N__22311));
    InMux I__4058 (
            .O(N__22314),
            .I(N__22308));
    LocalMux I__4057 (
            .O(N__22311),
            .I(N__22305));
    LocalMux I__4056 (
            .O(N__22308),
            .I(\POWERLED.CO2_THRU_CO ));
    Odrv4 I__4055 (
            .O(N__22305),
            .I(\POWERLED.CO2_THRU_CO ));
    InMux I__4054 (
            .O(N__22300),
            .I(N__22293));
    InMux I__4053 (
            .O(N__22299),
            .I(N__22293));
    InMux I__4052 (
            .O(N__22298),
            .I(N__22290));
    LocalMux I__4051 (
            .O(N__22293),
            .I(N__22287));
    LocalMux I__4050 (
            .O(N__22290),
            .I(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ));
    Odrv4 I__4049 (
            .O(N__22287),
            .I(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ));
    CascadeMux I__4048 (
            .O(N__22282),
            .I(N__22278));
    InMux I__4047 (
            .O(N__22281),
            .I(N__22269));
    InMux I__4046 (
            .O(N__22278),
            .I(N__22269));
    InMux I__4045 (
            .O(N__22277),
            .I(N__22269));
    InMux I__4044 (
            .O(N__22276),
            .I(N__22266));
    LocalMux I__4043 (
            .O(N__22269),
            .I(N__22263));
    LocalMux I__4042 (
            .O(N__22266),
            .I(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ));
    Odrv4 I__4041 (
            .O(N__22263),
            .I(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ));
    InMux I__4040 (
            .O(N__22258),
            .I(N__22255));
    LocalMux I__4039 (
            .O(N__22255),
            .I(\POWERLED.mult1_un89_sum_cry_6_s ));
    CascadeMux I__4038 (
            .O(N__22252),
            .I(N__22248));
    CascadeMux I__4037 (
            .O(N__22251),
            .I(N__22244));
    InMux I__4036 (
            .O(N__22248),
            .I(N__22237));
    InMux I__4035 (
            .O(N__22247),
            .I(N__22237));
    InMux I__4034 (
            .O(N__22244),
            .I(N__22237));
    LocalMux I__4033 (
            .O(N__22237),
            .I(\POWERLED.mult1_un89_sum_i_0_8 ));
    InMux I__4032 (
            .O(N__22234),
            .I(\POWERLED.mult1_un96_sum_cry_6 ));
    CascadeMux I__4031 (
            .O(N__22231),
            .I(N__22228));
    InMux I__4030 (
            .O(N__22228),
            .I(N__22225));
    LocalMux I__4029 (
            .O(N__22225),
            .I(\POWERLED.mult1_un96_sum_axb_8 ));
    InMux I__4028 (
            .O(N__22222),
            .I(\POWERLED.mult1_un96_sum_cry_7 ));
    CascadeMux I__4027 (
            .O(N__22219),
            .I(N__22215));
    CascadeMux I__4026 (
            .O(N__22218),
            .I(N__22211));
    InMux I__4025 (
            .O(N__22215),
            .I(N__22204));
    InMux I__4024 (
            .O(N__22214),
            .I(N__22204));
    InMux I__4023 (
            .O(N__22211),
            .I(N__22204));
    LocalMux I__4022 (
            .O(N__22204),
            .I(\POWERLED.mult1_un82_sum_i_0_8 ));
    InMux I__4021 (
            .O(N__22201),
            .I(N__22197));
    InMux I__4020 (
            .O(N__22200),
            .I(N__22194));
    LocalMux I__4019 (
            .O(N__22197),
            .I(N__22189));
    LocalMux I__4018 (
            .O(N__22194),
            .I(N__22189));
    Odrv4 I__4017 (
            .O(N__22189),
            .I(\POWERLED.mult1_un103_sum ));
    InMux I__4016 (
            .O(N__22186),
            .I(N__22183));
    LocalMux I__4015 (
            .O(N__22183),
            .I(N__22180));
    Odrv4 I__4014 (
            .O(N__22180),
            .I(\POWERLED.mult1_un96_sum_i ));
    CascadeMux I__4013 (
            .O(N__22177),
            .I(N__22174));
    InMux I__4012 (
            .O(N__22174),
            .I(N__22171));
    LocalMux I__4011 (
            .O(N__22171),
            .I(\POWERLED.mult1_un103_sum_cry_3_s ));
    InMux I__4010 (
            .O(N__22168),
            .I(\POWERLED.mult1_un103_sum_cry_2 ));
    CascadeMux I__4009 (
            .O(N__22165),
            .I(N__22162));
    InMux I__4008 (
            .O(N__22162),
            .I(N__22159));
    LocalMux I__4007 (
            .O(N__22159),
            .I(\POWERLED.mult1_un96_sum_cry_3_s ));
    InMux I__4006 (
            .O(N__22156),
            .I(N__22153));
    LocalMux I__4005 (
            .O(N__22153),
            .I(\POWERLED.mult1_un103_sum_cry_4_s ));
    InMux I__4004 (
            .O(N__22150),
            .I(\POWERLED.mult1_un103_sum_cry_3 ));
    CascadeMux I__4003 (
            .O(N__22147),
            .I(N__22144));
    InMux I__4002 (
            .O(N__22144),
            .I(N__22141));
    LocalMux I__4001 (
            .O(N__22141),
            .I(\POWERLED.mult1_un96_sum_cry_4_s ));
    CascadeMux I__4000 (
            .O(N__22138),
            .I(N__22135));
    InMux I__3999 (
            .O(N__22135),
            .I(N__22132));
    LocalMux I__3998 (
            .O(N__22132),
            .I(\POWERLED.mult1_un103_sum_cry_5_s ));
    InMux I__3997 (
            .O(N__22129),
            .I(\POWERLED.mult1_un103_sum_cry_4 ));
    InMux I__3996 (
            .O(N__22126),
            .I(N__22123));
    LocalMux I__3995 (
            .O(N__22123),
            .I(\POWERLED.mult1_un96_sum_cry_5_s ));
    InMux I__3994 (
            .O(N__22120),
            .I(N__22117));
    LocalMux I__3993 (
            .O(N__22117),
            .I(\POWERLED.mult1_un103_sum_cry_6_s ));
    InMux I__3992 (
            .O(N__22114),
            .I(\POWERLED.mult1_un103_sum_cry_5 ));
    InMux I__3991 (
            .O(N__22111),
            .I(\POWERLED.mult1_un89_sum_cry_6 ));
    InMux I__3990 (
            .O(N__22108),
            .I(\POWERLED.mult1_un89_sum_cry_7 ));
    CascadeMux I__3989 (
            .O(N__22105),
            .I(\POWERLED.mult1_un89_sum_s_8_cascade_ ));
    InMux I__3988 (
            .O(N__22102),
            .I(N__22098));
    InMux I__3987 (
            .O(N__22101),
            .I(N__22095));
    LocalMux I__3986 (
            .O(N__22098),
            .I(N__22090));
    LocalMux I__3985 (
            .O(N__22095),
            .I(N__22090));
    Span4Mux_s1_v I__3984 (
            .O(N__22090),
            .I(N__22087));
    Odrv4 I__3983 (
            .O(N__22087),
            .I(\POWERLED.mult1_un96_sum ));
    InMux I__3982 (
            .O(N__22084),
            .I(N__22081));
    LocalMux I__3981 (
            .O(N__22081),
            .I(\POWERLED.mult1_un89_sum_i ));
    InMux I__3980 (
            .O(N__22078),
            .I(\POWERLED.mult1_un96_sum_cry_2 ));
    CascadeMux I__3979 (
            .O(N__22075),
            .I(N__22072));
    InMux I__3978 (
            .O(N__22072),
            .I(N__22069));
    LocalMux I__3977 (
            .O(N__22069),
            .I(\POWERLED.mult1_un89_sum_cry_3_s ));
    InMux I__3976 (
            .O(N__22066),
            .I(\POWERLED.mult1_un96_sum_cry_3 ));
    InMux I__3975 (
            .O(N__22063),
            .I(N__22060));
    LocalMux I__3974 (
            .O(N__22060),
            .I(\POWERLED.mult1_un89_sum_cry_4_s ));
    InMux I__3973 (
            .O(N__22057),
            .I(\POWERLED.mult1_un96_sum_cry_4 ));
    CascadeMux I__3972 (
            .O(N__22054),
            .I(N__22049));
    InMux I__3971 (
            .O(N__22053),
            .I(N__22045));
    InMux I__3970 (
            .O(N__22052),
            .I(N__22040));
    InMux I__3969 (
            .O(N__22049),
            .I(N__22040));
    InMux I__3968 (
            .O(N__22048),
            .I(N__22037));
    LocalMux I__3967 (
            .O(N__22045),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__3966 (
            .O(N__22040),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__3965 (
            .O(N__22037),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    CascadeMux I__3964 (
            .O(N__22030),
            .I(N__22027));
    InMux I__3963 (
            .O(N__22027),
            .I(N__22024));
    LocalMux I__3962 (
            .O(N__22024),
            .I(\POWERLED.mult1_un89_sum_cry_5_s ));
    InMux I__3961 (
            .O(N__22021),
            .I(\POWERLED.mult1_un96_sum_cry_5 ));
    InMux I__3960 (
            .O(N__22018),
            .I(\VPP_VDDQ.un1_count_1_cry_12 ));
    InMux I__3959 (
            .O(N__22015),
            .I(\VPP_VDDQ.un1_count_1_cry_13 ));
    InMux I__3958 (
            .O(N__22012),
            .I(bfn_7_16_0_));
    CEMux I__3957 (
            .O(N__22009),
            .I(N__22006));
    LocalMux I__3956 (
            .O(N__22006),
            .I(N__22003));
    Span4Mux_s1_v I__3955 (
            .O(N__22003),
            .I(N__22000));
    Odrv4 I__3954 (
            .O(N__22000),
            .I(\VPP_VDDQ.N_42_0 ));
    SRMux I__3953 (
            .O(N__21997),
            .I(N__21994));
    LocalMux I__3952 (
            .O(N__21994),
            .I(N__21990));
    SRMux I__3951 (
            .O(N__21993),
            .I(N__21987));
    Span4Mux_v I__3950 (
            .O(N__21990),
            .I(N__21983));
    LocalMux I__3949 (
            .O(N__21987),
            .I(N__21980));
    SRMux I__3948 (
            .O(N__21986),
            .I(N__21977));
    Span4Mux_s2_v I__3947 (
            .O(N__21983),
            .I(N__21972));
    Span4Mux_s2_v I__3946 (
            .O(N__21980),
            .I(N__21972));
    LocalMux I__3945 (
            .O(N__21977),
            .I(N__21969));
    Odrv4 I__3944 (
            .O(N__21972),
            .I(G_44));
    Odrv12 I__3943 (
            .O(N__21969),
            .I(G_44));
    InMux I__3942 (
            .O(N__21964),
            .I(N__21960));
    InMux I__3941 (
            .O(N__21963),
            .I(N__21957));
    LocalMux I__3940 (
            .O(N__21960),
            .I(N__21952));
    LocalMux I__3939 (
            .O(N__21957),
            .I(N__21952));
    Span4Mux_s1_v I__3938 (
            .O(N__21952),
            .I(N__21949));
    Odrv4 I__3937 (
            .O(N__21949),
            .I(\POWERLED.mult1_un89_sum ));
    InMux I__3936 (
            .O(N__21946),
            .I(N__21943));
    LocalMux I__3935 (
            .O(N__21943),
            .I(\POWERLED.mult1_un82_sum_i ));
    InMux I__3934 (
            .O(N__21940),
            .I(\POWERLED.mult1_un89_sum_cry_2 ));
    InMux I__3933 (
            .O(N__21937),
            .I(\POWERLED.mult1_un89_sum_cry_3 ));
    InMux I__3932 (
            .O(N__21934),
            .I(\POWERLED.mult1_un89_sum_cry_4 ));
    InMux I__3931 (
            .O(N__21931),
            .I(\POWERLED.mult1_un89_sum_cry_5 ));
    InMux I__3930 (
            .O(N__21928),
            .I(\VPP_VDDQ.un1_count_1_cry_3 ));
    InMux I__3929 (
            .O(N__21925),
            .I(\VPP_VDDQ.un1_count_1_cry_4 ));
    InMux I__3928 (
            .O(N__21922),
            .I(\VPP_VDDQ.un1_count_1_cry_5 ));
    InMux I__3927 (
            .O(N__21919),
            .I(\VPP_VDDQ.un1_count_1_cry_6 ));
    InMux I__3926 (
            .O(N__21916),
            .I(bfn_7_15_0_));
    InMux I__3925 (
            .O(N__21913),
            .I(\VPP_VDDQ.un1_count_1_cry_8 ));
    InMux I__3924 (
            .O(N__21910),
            .I(\VPP_VDDQ.un1_count_1_cry_9 ));
    InMux I__3923 (
            .O(N__21907),
            .I(\VPP_VDDQ.un1_count_1_cry_10 ));
    InMux I__3922 (
            .O(N__21904),
            .I(\VPP_VDDQ.un1_count_1_cry_11 ));
    CascadeMux I__3921 (
            .O(N__21901),
            .I(G_44_cascade_));
    CascadeMux I__3920 (
            .O(N__21898),
            .I(N__21895));
    InMux I__3919 (
            .O(N__21895),
            .I(N__21892));
    LocalMux I__3918 (
            .O(N__21892),
            .I(N_365));
    CascadeMux I__3917 (
            .O(N__21889),
            .I(N__21885));
    InMux I__3916 (
            .O(N__21888),
            .I(N__21882));
    InMux I__3915 (
            .O(N__21885),
            .I(N__21879));
    LocalMux I__3914 (
            .O(N__21882),
            .I(\VPP_VDDQ.N_464_i ));
    LocalMux I__3913 (
            .O(N__21879),
            .I(\VPP_VDDQ.N_464_i ));
    InMux I__3912 (
            .O(N__21874),
            .I(\VPP_VDDQ.un1_count_1_cry_0 ));
    InMux I__3911 (
            .O(N__21871),
            .I(\VPP_VDDQ.un1_count_1_cry_1 ));
    InMux I__3910 (
            .O(N__21868),
            .I(\VPP_VDDQ.un1_count_1_cry_2 ));
    CascadeMux I__3909 (
            .O(N__21865),
            .I(\POWERLED.dutycycle_RNI79E14Z0Z_3_cascade_ ));
    CascadeMux I__3908 (
            .O(N__21862),
            .I(\POWERLED.dutycycleZ0Z_6_cascade_ ));
    InMux I__3907 (
            .O(N__21859),
            .I(N__21856));
    LocalMux I__3906 (
            .O(N__21856),
            .I(\POWERLED.dutycycle_eena_8_c ));
    InMux I__3905 (
            .O(N__21853),
            .I(N__21850));
    LocalMux I__3904 (
            .O(N__21850),
            .I(\POWERLED.dutycycle_RNI79E14Z0Z_3 ));
    CascadeMux I__3903 (
            .O(N__21847),
            .I(N__21844));
    InMux I__3902 (
            .O(N__21844),
            .I(N__21840));
    InMux I__3901 (
            .O(N__21843),
            .I(N__21837));
    LocalMux I__3900 (
            .O(N__21840),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__3899 (
            .O(N__21837),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    InMux I__3898 (
            .O(N__21832),
            .I(N__21829));
    LocalMux I__3897 (
            .O(N__21829),
            .I(N__21825));
    CascadeMux I__3896 (
            .O(N__21828),
            .I(N__21822));
    Span4Mux_v I__3895 (
            .O(N__21825),
            .I(N__21819));
    InMux I__3894 (
            .O(N__21822),
            .I(N__21816));
    Odrv4 I__3893 (
            .O(N__21819),
            .I(\POWERLED.N_2168_i ));
    LocalMux I__3892 (
            .O(N__21816),
            .I(\POWERLED.N_2168_i ));
    CascadeMux I__3891 (
            .O(N__21811),
            .I(\POWERLED.N_231_i_cascade_ ));
    InMux I__3890 (
            .O(N__21808),
            .I(N__21804));
    InMux I__3889 (
            .O(N__21807),
            .I(N__21801));
    LocalMux I__3888 (
            .O(N__21804),
            .I(N__21798));
    LocalMux I__3887 (
            .O(N__21801),
            .I(N__21795));
    Span4Mux_h I__3886 (
            .O(N__21798),
            .I(N__21790));
    Span4Mux_h I__3885 (
            .O(N__21795),
            .I(N__21790));
    Odrv4 I__3884 (
            .O(N__21790),
            .I(\POWERLED.N_321 ));
    InMux I__3883 (
            .O(N__21787),
            .I(N__21784));
    LocalMux I__3882 (
            .O(N__21784),
            .I(\POWERLED.N_52_i_i_0 ));
    CascadeMux I__3881 (
            .O(N__21781),
            .I(\POWERLED.N_410_cascade_ ));
    InMux I__3880 (
            .O(N__21778),
            .I(N__21775));
    LocalMux I__3879 (
            .O(N__21775),
            .I(N__21771));
    InMux I__3878 (
            .O(N__21774),
            .I(N__21768));
    Span4Mux_v I__3877 (
            .O(N__21771),
            .I(N__21765));
    LocalMux I__3876 (
            .O(N__21768),
            .I(N__21762));
    Odrv4 I__3875 (
            .O(N__21765),
            .I(\POWERLED.func_state_RNI1J4E2Z0Z_1 ));
    Odrv4 I__3874 (
            .O(N__21762),
            .I(\POWERLED.func_state_RNI1J4E2Z0Z_1 ));
    InMux I__3873 (
            .O(N__21757),
            .I(N__21754));
    LocalMux I__3872 (
            .O(N__21754),
            .I(N__21744));
    InMux I__3871 (
            .O(N__21753),
            .I(N__21741));
    InMux I__3870 (
            .O(N__21752),
            .I(N__21738));
    InMux I__3869 (
            .O(N__21751),
            .I(N__21735));
    InMux I__3868 (
            .O(N__21750),
            .I(N__21730));
    InMux I__3867 (
            .O(N__21749),
            .I(N__21730));
    InMux I__3866 (
            .O(N__21748),
            .I(N__21727));
    CascadeMux I__3865 (
            .O(N__21747),
            .I(N__21719));
    Span4Mux_v I__3864 (
            .O(N__21744),
            .I(N__21713));
    LocalMux I__3863 (
            .O(N__21741),
            .I(N__21713));
    LocalMux I__3862 (
            .O(N__21738),
            .I(N__21710));
    LocalMux I__3861 (
            .O(N__21735),
            .I(N__21705));
    LocalMux I__3860 (
            .O(N__21730),
            .I(N__21705));
    LocalMux I__3859 (
            .O(N__21727),
            .I(N__21702));
    InMux I__3858 (
            .O(N__21726),
            .I(N__21697));
    InMux I__3857 (
            .O(N__21725),
            .I(N__21697));
    InMux I__3856 (
            .O(N__21724),
            .I(N__21686));
    InMux I__3855 (
            .O(N__21723),
            .I(N__21686));
    InMux I__3854 (
            .O(N__21722),
            .I(N__21686));
    InMux I__3853 (
            .O(N__21719),
            .I(N__21686));
    InMux I__3852 (
            .O(N__21718),
            .I(N__21686));
    Span4Mux_h I__3851 (
            .O(N__21713),
            .I(N__21681));
    Span4Mux_h I__3850 (
            .O(N__21710),
            .I(N__21681));
    Span4Mux_h I__3849 (
            .O(N__21705),
            .I(N__21678));
    Odrv4 I__3848 (
            .O(N__21702),
            .I(COUNTER_un4_counter_7_THRU_CO));
    LocalMux I__3847 (
            .O(N__21697),
            .I(COUNTER_un4_counter_7_THRU_CO));
    LocalMux I__3846 (
            .O(N__21686),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv4 I__3845 (
            .O(N__21681),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv4 I__3844 (
            .O(N__21678),
            .I(COUNTER_un4_counter_7_THRU_CO));
    CascadeMux I__3843 (
            .O(N__21667),
            .I(N__21663));
    InMux I__3842 (
            .O(N__21666),
            .I(N__21660));
    InMux I__3841 (
            .O(N__21663),
            .I(N__21657));
    LocalMux I__3840 (
            .O(N__21660),
            .I(N__21654));
    LocalMux I__3839 (
            .O(N__21657),
            .I(\POWERLED.dutycycleZ1Z_7 ));
    Odrv12 I__3838 (
            .O(N__21654),
            .I(\POWERLED.dutycycleZ1Z_7 ));
    CascadeMux I__3837 (
            .O(N__21649),
            .I(\POWERLED.dutycycle_RNI375F3Z0Z_7_cascade_ ));
    CascadeMux I__3836 (
            .O(N__21646),
            .I(\POWERLED.dutycycleZ0Z_4_cascade_ ));
    InMux I__3835 (
            .O(N__21643),
            .I(N__21640));
    LocalMux I__3834 (
            .O(N__21640),
            .I(\RSMRST_PWRGD.N_8_mux ));
    CascadeMux I__3833 (
            .O(N__21637),
            .I(m57_i_o2_2_cascade_));
    CascadeMux I__3832 (
            .O(N__21634),
            .I(\RSMRST_PWRGD.N_4713_0_0_0_cascade_ ));
    CascadeMux I__3831 (
            .O(N__21631),
            .I(\POWERLED.N_569_N_cascade_ ));
    CascadeMux I__3830 (
            .O(N__21628),
            .I(\POWERLED.N_220_N_cascade_ ));
    CascadeMux I__3829 (
            .O(N__21625),
            .I(\POWERLED.N_282_N_cascade_ ));
    CascadeMux I__3828 (
            .O(N__21622),
            .I(\POWERLED.dutycycle_eena_8_d_cascade_ ));
    CascadeMux I__3827 (
            .O(N__21619),
            .I(func_state_RNITGMHB_0_1_cascade_));
    CascadeMux I__3826 (
            .O(N__21616),
            .I(N__21613));
    InMux I__3825 (
            .O(N__21613),
            .I(N__21610));
    LocalMux I__3824 (
            .O(N__21610),
            .I(N__21607));
    Odrv12 I__3823 (
            .O(N__21607),
            .I(\POWERLED.dutycycle_RNIZ0Z_3 ));
    InMux I__3822 (
            .O(N__21604),
            .I(N__21598));
    InMux I__3821 (
            .O(N__21603),
            .I(N__21598));
    LocalMux I__3820 (
            .O(N__21598),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_1 ));
    CascadeMux I__3819 (
            .O(N__21595),
            .I(N__21592));
    InMux I__3818 (
            .O(N__21592),
            .I(N__21589));
    LocalMux I__3817 (
            .O(N__21589),
            .I(N__21586));
    Odrv12 I__3816 (
            .O(N__21586),
            .I(\POWERLED.dutycycle_RNIZ0Z_2 ));
    InMux I__3815 (
            .O(N__21583),
            .I(N__21577));
    InMux I__3814 (
            .O(N__21582),
            .I(N__21577));
    LocalMux I__3813 (
            .O(N__21577),
            .I(\POWERLED.func_state_RNICK8N9Z0Z_1 ));
    CascadeMux I__3812 (
            .O(N__21574),
            .I(N__21570));
    InMux I__3811 (
            .O(N__21573),
            .I(N__21565));
    InMux I__3810 (
            .O(N__21570),
            .I(N__21565));
    LocalMux I__3809 (
            .O(N__21565),
            .I(\POWERLED.func_stateZ0Z_1 ));
    InMux I__3808 (
            .O(N__21562),
            .I(N__21558));
    InMux I__3807 (
            .O(N__21561),
            .I(N__21555));
    LocalMux I__3806 (
            .O(N__21558),
            .I(N__21552));
    LocalMux I__3805 (
            .O(N__21555),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_3 ));
    Odrv12 I__3804 (
            .O(N__21552),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_3 ));
    CascadeMux I__3803 (
            .O(N__21547),
            .I(\POWERLED.N_80_f0_cascade_ ));
    InMux I__3802 (
            .O(N__21544),
            .I(N__21541));
    LocalMux I__3801 (
            .O(N__21541),
            .I(N__21538));
    Odrv12 I__3800 (
            .O(N__21538),
            .I(\POWERLED.dutycycle_RNI375F3Z0Z_7 ));
    CascadeMux I__3799 (
            .O(N__21535),
            .I(N__21532));
    InMux I__3798 (
            .O(N__21532),
            .I(N__21529));
    LocalMux I__3797 (
            .O(N__21529),
            .I(N__21526));
    Odrv4 I__3796 (
            .O(N__21526),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_1 ));
    InMux I__3795 (
            .O(N__21523),
            .I(N__21520));
    LocalMux I__3794 (
            .O(N__21520),
            .I(\POWERLED.mult1_un159_sum_i ));
    InMux I__3793 (
            .O(N__21517),
            .I(N__21514));
    LocalMux I__3792 (
            .O(N__21514),
            .I(N__21511));
    Odrv12 I__3791 (
            .O(N__21511),
            .I(\POWERLED.mult1_un152_sum_i ));
    InMux I__3790 (
            .O(N__21508),
            .I(N__21505));
    LocalMux I__3789 (
            .O(N__21505),
            .I(\POWERLED.func_state_1_m0_i_o2_0_1 ));
    InMux I__3788 (
            .O(N__21502),
            .I(N__21499));
    LocalMux I__3787 (
            .O(N__21499),
            .I(N_21));
    InMux I__3786 (
            .O(N__21496),
            .I(\POWERLED.un1_dutycycle_53_cry_10 ));
    InMux I__3785 (
            .O(N__21493),
            .I(\POWERLED.un1_dutycycle_53_cry_11 ));
    InMux I__3784 (
            .O(N__21490),
            .I(\POWERLED.un1_dutycycle_53_cry_12 ));
    InMux I__3783 (
            .O(N__21487),
            .I(\POWERLED.un1_dutycycle_53_cry_13 ));
    InMux I__3782 (
            .O(N__21484),
            .I(\POWERLED.un1_dutycycle_53_cry_14 ));
    InMux I__3781 (
            .O(N__21481),
            .I(bfn_7_7_0_));
    InMux I__3780 (
            .O(N__21478),
            .I(\POWERLED.CO2 ));
    InMux I__3779 (
            .O(N__21475),
            .I(N__21472));
    LocalMux I__3778 (
            .O(N__21472),
            .I(\POWERLED.N_76_f0 ));
    InMux I__3777 (
            .O(N__21469),
            .I(N__21465));
    InMux I__3776 (
            .O(N__21468),
            .I(N__21462));
    LocalMux I__3775 (
            .O(N__21465),
            .I(N__21459));
    LocalMux I__3774 (
            .O(N__21462),
            .I(N__21454));
    Span4Mux_v I__3773 (
            .O(N__21459),
            .I(N__21454));
    Odrv4 I__3772 (
            .O(N__21454),
            .I(\POWERLED.mult1_un124_sum ));
    InMux I__3771 (
            .O(N__21451),
            .I(\POWERLED.un1_dutycycle_53_cry_2_cZ0 ));
    InMux I__3770 (
            .O(N__21448),
            .I(N__21444));
    InMux I__3769 (
            .O(N__21447),
            .I(N__21441));
    LocalMux I__3768 (
            .O(N__21444),
            .I(\POWERLED.mult1_un117_sum ));
    LocalMux I__3767 (
            .O(N__21441),
            .I(\POWERLED.mult1_un117_sum ));
    InMux I__3766 (
            .O(N__21436),
            .I(\POWERLED.un1_dutycycle_53_cry_3_cZ0 ));
    InMux I__3765 (
            .O(N__21433),
            .I(N__21429));
    InMux I__3764 (
            .O(N__21432),
            .I(N__21426));
    LocalMux I__3763 (
            .O(N__21429),
            .I(N__21423));
    LocalMux I__3762 (
            .O(N__21426),
            .I(\POWERLED.mult1_un110_sum ));
    Odrv4 I__3761 (
            .O(N__21423),
            .I(\POWERLED.mult1_un110_sum ));
    InMux I__3760 (
            .O(N__21418),
            .I(\POWERLED.un1_dutycycle_53_cry_4_cZ0 ));
    InMux I__3759 (
            .O(N__21415),
            .I(\POWERLED.un1_dutycycle_53_cry_5_cZ0 ));
    InMux I__3758 (
            .O(N__21412),
            .I(\POWERLED.un1_dutycycle_53_cry_6_cZ0 ));
    InMux I__3757 (
            .O(N__21409),
            .I(bfn_7_6_0_));
    InMux I__3756 (
            .O(N__21406),
            .I(\POWERLED.un1_dutycycle_53_cry_8 ));
    InMux I__3755 (
            .O(N__21403),
            .I(\POWERLED.un1_dutycycle_53_cry_9 ));
    InMux I__3754 (
            .O(N__21400),
            .I(N__21397));
    LocalMux I__3753 (
            .O(N__21397),
            .I(N__21394));
    Odrv4 I__3752 (
            .O(N__21394),
            .I(\POWERLED.mult1_un110_sum_cry_4_s ));
    InMux I__3751 (
            .O(N__21391),
            .I(\POWERLED.mult1_un110_sum_cry_3 ));
    CascadeMux I__3750 (
            .O(N__21388),
            .I(N__21385));
    InMux I__3749 (
            .O(N__21385),
            .I(N__21382));
    LocalMux I__3748 (
            .O(N__21382),
            .I(N__21379));
    Odrv4 I__3747 (
            .O(N__21379),
            .I(\POWERLED.mult1_un110_sum_cry_5_s ));
    InMux I__3746 (
            .O(N__21376),
            .I(\POWERLED.mult1_un110_sum_cry_4 ));
    InMux I__3745 (
            .O(N__21373),
            .I(N__21370));
    LocalMux I__3744 (
            .O(N__21370),
            .I(N__21367));
    Span4Mux_h I__3743 (
            .O(N__21367),
            .I(N__21364));
    Odrv4 I__3742 (
            .O(N__21364),
            .I(\POWERLED.mult1_un110_sum_cry_6_s ));
    InMux I__3741 (
            .O(N__21361),
            .I(\POWERLED.mult1_un110_sum_cry_5 ));
    CascadeMux I__3740 (
            .O(N__21358),
            .I(N__21354));
    CascadeMux I__3739 (
            .O(N__21357),
            .I(N__21350));
    InMux I__3738 (
            .O(N__21354),
            .I(N__21343));
    InMux I__3737 (
            .O(N__21353),
            .I(N__21343));
    InMux I__3736 (
            .O(N__21350),
            .I(N__21343));
    LocalMux I__3735 (
            .O(N__21343),
            .I(\POWERLED.mult1_un103_sum_i_0_8 ));
    InMux I__3734 (
            .O(N__21340),
            .I(N__21337));
    LocalMux I__3733 (
            .O(N__21337),
            .I(N__21334));
    Odrv4 I__3732 (
            .O(N__21334),
            .I(\POWERLED.mult1_un117_sum_axb_8 ));
    InMux I__3731 (
            .O(N__21331),
            .I(\POWERLED.mult1_un110_sum_cry_6 ));
    InMux I__3730 (
            .O(N__21328),
            .I(\POWERLED.mult1_un110_sum_cry_7 ));
    CascadeMux I__3729 (
            .O(N__21325),
            .I(N__21321));
    InMux I__3728 (
            .O(N__21324),
            .I(N__21315));
    InMux I__3727 (
            .O(N__21321),
            .I(N__21315));
    InMux I__3726 (
            .O(N__21320),
            .I(N__21310));
    LocalMux I__3725 (
            .O(N__21315),
            .I(N__21307));
    InMux I__3724 (
            .O(N__21314),
            .I(N__21304));
    InMux I__3723 (
            .O(N__21313),
            .I(N__21301));
    LocalMux I__3722 (
            .O(N__21310),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    Odrv4 I__3721 (
            .O(N__21307),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__3720 (
            .O(N__21304),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__3719 (
            .O(N__21301),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    InMux I__3718 (
            .O(N__21292),
            .I(N__21289));
    LocalMux I__3717 (
            .O(N__21289),
            .I(\POWERLED.un85_clk_100khz_12 ));
    InMux I__3716 (
            .O(N__21286),
            .I(N__21283));
    LocalMux I__3715 (
            .O(N__21283),
            .I(N__21279));
    InMux I__3714 (
            .O(N__21282),
            .I(N__21276));
    Span4Mux_v I__3713 (
            .O(N__21279),
            .I(N__21271));
    LocalMux I__3712 (
            .O(N__21276),
            .I(N__21271));
    Odrv4 I__3711 (
            .O(N__21271),
            .I(\POWERLED.mult1_un145_sum ));
    InMux I__3710 (
            .O(N__21268),
            .I(N__21264));
    InMux I__3709 (
            .O(N__21267),
            .I(N__21261));
    LocalMux I__3708 (
            .O(N__21264),
            .I(N__21258));
    LocalMux I__3707 (
            .O(N__21261),
            .I(\POWERLED.mult1_un138_sum ));
    Odrv12 I__3706 (
            .O(N__21258),
            .I(\POWERLED.mult1_un138_sum ));
    InMux I__3705 (
            .O(N__21253),
            .I(\POWERLED.un1_dutycycle_53_cry_0_cZ0 ));
    InMux I__3704 (
            .O(N__21250),
            .I(N__21247));
    LocalMux I__3703 (
            .O(N__21247),
            .I(N__21243));
    InMux I__3702 (
            .O(N__21246),
            .I(N__21240));
    Span4Mux_h I__3701 (
            .O(N__21243),
            .I(N__21237));
    LocalMux I__3700 (
            .O(N__21240),
            .I(\POWERLED.mult1_un131_sum ));
    Odrv4 I__3699 (
            .O(N__21237),
            .I(\POWERLED.mult1_un131_sum ));
    InMux I__3698 (
            .O(N__21232),
            .I(\POWERLED.un1_dutycycle_53_cry_1_cZ0 ));
    InMux I__3697 (
            .O(N__21229),
            .I(N__21226));
    LocalMux I__3696 (
            .O(N__21226),
            .I(\POWERLED.un85_clk_100khz_9 ));
    InMux I__3695 (
            .O(N__21223),
            .I(N__21220));
    LocalMux I__3694 (
            .O(N__21220),
            .I(\POWERLED.un85_clk_100khz_8 ));
    InMux I__3693 (
            .O(N__21217),
            .I(N__21214));
    LocalMux I__3692 (
            .O(N__21214),
            .I(N__21211));
    Odrv4 I__3691 (
            .O(N__21211),
            .I(\POWERLED.mult1_un103_sum_i ));
    CascadeMux I__3690 (
            .O(N__21208),
            .I(N__21205));
    InMux I__3689 (
            .O(N__21205),
            .I(N__21202));
    LocalMux I__3688 (
            .O(N__21202),
            .I(N__21199));
    Odrv4 I__3687 (
            .O(N__21199),
            .I(\POWERLED.mult1_un110_sum_cry_3_s ));
    InMux I__3686 (
            .O(N__21196),
            .I(\POWERLED.mult1_un110_sum_cry_2 ));
    InMux I__3685 (
            .O(N__21193),
            .I(N__21190));
    LocalMux I__3684 (
            .O(N__21190),
            .I(N__21187));
    Span4Mux_s1_v I__3683 (
            .O(N__21187),
            .I(N__21184));
    Span4Mux_h I__3682 (
            .O(N__21184),
            .I(N__21180));
    InMux I__3681 (
            .O(N__21183),
            .I(N__21177));
    Odrv4 I__3680 (
            .O(N__21180),
            .I(\PCH_PWRGD.count_rst_8 ));
    LocalMux I__3679 (
            .O(N__21177),
            .I(\PCH_PWRGD.count_rst_8 ));
    InMux I__3678 (
            .O(N__21172),
            .I(N__21169));
    LocalMux I__3677 (
            .O(N__21169),
            .I(N__21166));
    Span4Mux_s2_h I__3676 (
            .O(N__21166),
            .I(N__21163));
    Span4Mux_h I__3675 (
            .O(N__21163),
            .I(N__21160));
    Odrv4 I__3674 (
            .O(N__21160),
            .I(\PCH_PWRGD.count_0_6 ));
    CEMux I__3673 (
            .O(N__21157),
            .I(N__21147));
    InMux I__3672 (
            .O(N__21156),
            .I(N__21139));
    CEMux I__3671 (
            .O(N__21155),
            .I(N__21139));
    InMux I__3670 (
            .O(N__21154),
            .I(N__21134));
    CEMux I__3669 (
            .O(N__21153),
            .I(N__21134));
    InMux I__3668 (
            .O(N__21152),
            .I(N__21127));
    InMux I__3667 (
            .O(N__21151),
            .I(N__21127));
    CEMux I__3666 (
            .O(N__21150),
            .I(N__21127));
    LocalMux I__3665 (
            .O(N__21147),
            .I(N__21122));
    CEMux I__3664 (
            .O(N__21146),
            .I(N__21119));
    InMux I__3663 (
            .O(N__21145),
            .I(N__21114));
    InMux I__3662 (
            .O(N__21144),
            .I(N__21114));
    LocalMux I__3661 (
            .O(N__21139),
            .I(N__21109));
    LocalMux I__3660 (
            .O(N__21134),
            .I(N__21106));
    LocalMux I__3659 (
            .O(N__21127),
            .I(N__21103));
    InMux I__3658 (
            .O(N__21126),
            .I(N__21091));
    InMux I__3657 (
            .O(N__21125),
            .I(N__21091));
    Span4Mux_h I__3656 (
            .O(N__21122),
            .I(N__21088));
    LocalMux I__3655 (
            .O(N__21119),
            .I(N__21085));
    LocalMux I__3654 (
            .O(N__21114),
            .I(N__21082));
    InMux I__3653 (
            .O(N__21113),
            .I(N__21077));
    InMux I__3652 (
            .O(N__21112),
            .I(N__21077));
    Span4Mux_s2_v I__3651 (
            .O(N__21109),
            .I(N__21065));
    Span4Mux_h I__3650 (
            .O(N__21106),
            .I(N__21065));
    Span4Mux_s2_v I__3649 (
            .O(N__21103),
            .I(N__21065));
    InMux I__3648 (
            .O(N__21102),
            .I(N__21062));
    CEMux I__3647 (
            .O(N__21101),
            .I(N__21053));
    InMux I__3646 (
            .O(N__21100),
            .I(N__21053));
    InMux I__3645 (
            .O(N__21099),
            .I(N__21053));
    InMux I__3644 (
            .O(N__21098),
            .I(N__21053));
    CEMux I__3643 (
            .O(N__21097),
            .I(N__21048));
    InMux I__3642 (
            .O(N__21096),
            .I(N__21048));
    LocalMux I__3641 (
            .O(N__21091),
            .I(N__21045));
    Span4Mux_h I__3640 (
            .O(N__21088),
            .I(N__21036));
    Span4Mux_s0_v I__3639 (
            .O(N__21085),
            .I(N__21036));
    Span4Mux_s1_h I__3638 (
            .O(N__21082),
            .I(N__21036));
    LocalMux I__3637 (
            .O(N__21077),
            .I(N__21036));
    CEMux I__3636 (
            .O(N__21076),
            .I(N__21025));
    InMux I__3635 (
            .O(N__21075),
            .I(N__21025));
    InMux I__3634 (
            .O(N__21074),
            .I(N__21025));
    InMux I__3633 (
            .O(N__21073),
            .I(N__21025));
    InMux I__3632 (
            .O(N__21072),
            .I(N__21025));
    Odrv4 I__3631 (
            .O(N__21065),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    LocalMux I__3630 (
            .O(N__21062),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    LocalMux I__3629 (
            .O(N__21053),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    LocalMux I__3628 (
            .O(N__21048),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    Odrv4 I__3627 (
            .O(N__21045),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    Odrv4 I__3626 (
            .O(N__21036),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    LocalMux I__3625 (
            .O(N__21025),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    SRMux I__3624 (
            .O(N__21010),
            .I(N__21007));
    LocalMux I__3623 (
            .O(N__21007),
            .I(N__21002));
    SRMux I__3622 (
            .O(N__21006),
            .I(N__20999));
    SRMux I__3621 (
            .O(N__21005),
            .I(N__20993));
    Span4Mux_v I__3620 (
            .O(N__21002),
            .I(N__20988));
    LocalMux I__3619 (
            .O(N__20999),
            .I(N__20988));
    InMux I__3618 (
            .O(N__20998),
            .I(N__20979));
    SRMux I__3617 (
            .O(N__20997),
            .I(N__20979));
    SRMux I__3616 (
            .O(N__20996),
            .I(N__20973));
    LocalMux I__3615 (
            .O(N__20993),
            .I(N__20962));
    Span4Mux_s1_v I__3614 (
            .O(N__20988),
            .I(N__20959));
    InMux I__3613 (
            .O(N__20987),
            .I(N__20950));
    InMux I__3612 (
            .O(N__20986),
            .I(N__20950));
    InMux I__3611 (
            .O(N__20985),
            .I(N__20950));
    InMux I__3610 (
            .O(N__20984),
            .I(N__20950));
    LocalMux I__3609 (
            .O(N__20979),
            .I(N__20944));
    SRMux I__3608 (
            .O(N__20978),
            .I(N__20941));
    SRMux I__3607 (
            .O(N__20977),
            .I(N__20938));
    SRMux I__3606 (
            .O(N__20976),
            .I(N__20935));
    LocalMux I__3605 (
            .O(N__20973),
            .I(N__20932));
    CascadeMux I__3604 (
            .O(N__20972),
            .I(N__20926));
    InMux I__3603 (
            .O(N__20971),
            .I(N__20922));
    InMux I__3602 (
            .O(N__20970),
            .I(N__20911));
    InMux I__3601 (
            .O(N__20969),
            .I(N__20911));
    InMux I__3600 (
            .O(N__20968),
            .I(N__20911));
    InMux I__3599 (
            .O(N__20967),
            .I(N__20911));
    InMux I__3598 (
            .O(N__20966),
            .I(N__20911));
    CascadeMux I__3597 (
            .O(N__20965),
            .I(N__20908));
    Span4Mux_s1_v I__3596 (
            .O(N__20962),
            .I(N__20901));
    Span4Mux_s1_h I__3595 (
            .O(N__20959),
            .I(N__20901));
    LocalMux I__3594 (
            .O(N__20950),
            .I(N__20901));
    InMux I__3593 (
            .O(N__20949),
            .I(N__20896));
    InMux I__3592 (
            .O(N__20948),
            .I(N__20896));
    CascadeMux I__3591 (
            .O(N__20947),
            .I(N__20893));
    Span4Mux_s2_v I__3590 (
            .O(N__20944),
            .I(N__20886));
    LocalMux I__3589 (
            .O(N__20941),
            .I(N__20886));
    LocalMux I__3588 (
            .O(N__20938),
            .I(N__20883));
    LocalMux I__3587 (
            .O(N__20935),
            .I(N__20880));
    Span4Mux_s3_v I__3586 (
            .O(N__20932),
            .I(N__20877));
    CascadeMux I__3585 (
            .O(N__20931),
            .I(N__20869));
    InMux I__3584 (
            .O(N__20930),
            .I(N__20860));
    InMux I__3583 (
            .O(N__20929),
            .I(N__20860));
    InMux I__3582 (
            .O(N__20926),
            .I(N__20860));
    InMux I__3581 (
            .O(N__20925),
            .I(N__20860));
    LocalMux I__3580 (
            .O(N__20922),
            .I(N__20855));
    LocalMux I__3579 (
            .O(N__20911),
            .I(N__20855));
    InMux I__3578 (
            .O(N__20908),
            .I(N__20852));
    Span4Mux_v I__3577 (
            .O(N__20901),
            .I(N__20847));
    LocalMux I__3576 (
            .O(N__20896),
            .I(N__20847));
    InMux I__3575 (
            .O(N__20893),
            .I(N__20842));
    InMux I__3574 (
            .O(N__20892),
            .I(N__20842));
    InMux I__3573 (
            .O(N__20891),
            .I(N__20839));
    Span4Mux_h I__3572 (
            .O(N__20886),
            .I(N__20836));
    Span4Mux_s2_h I__3571 (
            .O(N__20883),
            .I(N__20829));
    Span4Mux_s3_v I__3570 (
            .O(N__20880),
            .I(N__20829));
    Span4Mux_h I__3569 (
            .O(N__20877),
            .I(N__20829));
    InMux I__3568 (
            .O(N__20876),
            .I(N__20824));
    InMux I__3567 (
            .O(N__20875),
            .I(N__20824));
    InMux I__3566 (
            .O(N__20874),
            .I(N__20815));
    InMux I__3565 (
            .O(N__20873),
            .I(N__20815));
    InMux I__3564 (
            .O(N__20872),
            .I(N__20815));
    InMux I__3563 (
            .O(N__20869),
            .I(N__20815));
    LocalMux I__3562 (
            .O(N__20860),
            .I(N__20812));
    Span4Mux_s1_v I__3561 (
            .O(N__20855),
            .I(N__20801));
    LocalMux I__3560 (
            .O(N__20852),
            .I(N__20801));
    Span4Mux_s1_h I__3559 (
            .O(N__20847),
            .I(N__20801));
    LocalMux I__3558 (
            .O(N__20842),
            .I(N__20801));
    LocalMux I__3557 (
            .O(N__20839),
            .I(N__20801));
    Odrv4 I__3556 (
            .O(N__20836),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__3555 (
            .O(N__20829),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    LocalMux I__3554 (
            .O(N__20824),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    LocalMux I__3553 (
            .O(N__20815),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv12 I__3552 (
            .O(N__20812),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__3551 (
            .O(N__20801),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    InMux I__3550 (
            .O(N__20788),
            .I(N__20785));
    LocalMux I__3549 (
            .O(N__20785),
            .I(N__20781));
    InMux I__3548 (
            .O(N__20784),
            .I(N__20778));
    Span4Mux_h I__3547 (
            .O(N__20781),
            .I(N__20773));
    LocalMux I__3546 (
            .O(N__20778),
            .I(N__20773));
    Span4Mux_v I__3545 (
            .O(N__20773),
            .I(N__20767));
    InMux I__3544 (
            .O(N__20772),
            .I(N__20762));
    InMux I__3543 (
            .O(N__20771),
            .I(N__20762));
    InMux I__3542 (
            .O(N__20770),
            .I(N__20759));
    Odrv4 I__3541 (
            .O(N__20767),
            .I(N_355));
    LocalMux I__3540 (
            .O(N__20762),
            .I(N_355));
    LocalMux I__3539 (
            .O(N__20759),
            .I(N_355));
    IoInMux I__3538 (
            .O(N__20752),
            .I(N__20749));
    LocalMux I__3537 (
            .O(N__20749),
            .I(N__20746));
    IoSpan4Mux I__3536 (
            .O(N__20746),
            .I(N__20743));
    Span4Mux_s2_h I__3535 (
            .O(N__20743),
            .I(N__20740));
    Span4Mux_v I__3534 (
            .O(N__20740),
            .I(N__20736));
    IoInMux I__3533 (
            .O(N__20739),
            .I(N__20733));
    Span4Mux_v I__3532 (
            .O(N__20736),
            .I(N__20730));
    LocalMux I__3531 (
            .O(N__20733),
            .I(N__20727));
    Span4Mux_v I__3530 (
            .O(N__20730),
            .I(N__20724));
    Span12Mux_s6_h I__3529 (
            .O(N__20727),
            .I(N__20721));
    Odrv4 I__3528 (
            .O(N__20724),
            .I(pch_pwrok));
    Odrv12 I__3527 (
            .O(N__20721),
            .I(pch_pwrok));
    InMux I__3526 (
            .O(N__20716),
            .I(N__20713));
    LocalMux I__3525 (
            .O(N__20713),
            .I(N__20710));
    Odrv4 I__3524 (
            .O(N__20710),
            .I(\POWERLED.mult1_un68_sum_i_8 ));
    CascadeMux I__3523 (
            .O(N__20707),
            .I(N__20704));
    InMux I__3522 (
            .O(N__20704),
            .I(N__20701));
    LocalMux I__3521 (
            .O(N__20701),
            .I(N__20698));
    Odrv4 I__3520 (
            .O(N__20698),
            .I(\POWERLED.mult1_un75_sum_i_8 ));
    InMux I__3519 (
            .O(N__20695),
            .I(N__20689));
    InMux I__3518 (
            .O(N__20694),
            .I(N__20689));
    LocalMux I__3517 (
            .O(N__20689),
            .I(N__20686));
    Odrv4 I__3516 (
            .O(N__20686),
            .I(\POWERLED.count_off_1_7 ));
    InMux I__3515 (
            .O(N__20683),
            .I(N__20680));
    LocalMux I__3514 (
            .O(N__20680),
            .I(\POWERLED.count_off_0_7 ));
    InMux I__3513 (
            .O(N__20677),
            .I(N__20673));
    InMux I__3512 (
            .O(N__20676),
            .I(N__20670));
    LocalMux I__3511 (
            .O(N__20673),
            .I(N__20665));
    LocalMux I__3510 (
            .O(N__20670),
            .I(N__20665));
    Odrv4 I__3509 (
            .O(N__20665),
            .I(\POWERLED.count_offZ0Z_8 ));
    InMux I__3508 (
            .O(N__20662),
            .I(N__20656));
    InMux I__3507 (
            .O(N__20661),
            .I(N__20656));
    LocalMux I__3506 (
            .O(N__20656),
            .I(N__20653));
    Odrv4 I__3505 (
            .O(N__20653),
            .I(\POWERLED.count_off_1_8 ));
    InMux I__3504 (
            .O(N__20650),
            .I(N__20647));
    LocalMux I__3503 (
            .O(N__20647),
            .I(\POWERLED.count_off_0_8 ));
    InMux I__3502 (
            .O(N__20644),
            .I(N__20640));
    InMux I__3501 (
            .O(N__20643),
            .I(N__20637));
    LocalMux I__3500 (
            .O(N__20640),
            .I(\POWERLED.count_off_1_9 ));
    LocalMux I__3499 (
            .O(N__20637),
            .I(\POWERLED.count_off_1_9 ));
    InMux I__3498 (
            .O(N__20632),
            .I(N__20629));
    LocalMux I__3497 (
            .O(N__20629),
            .I(\POWERLED.count_off_0_9 ));
    CEMux I__3496 (
            .O(N__20626),
            .I(N__20622));
    CEMux I__3495 (
            .O(N__20625),
            .I(N__20618));
    LocalMux I__3494 (
            .O(N__20622),
            .I(N__20614));
    CEMux I__3493 (
            .O(N__20621),
            .I(N__20611));
    LocalMux I__3492 (
            .O(N__20618),
            .I(N__20607));
    CEMux I__3491 (
            .O(N__20617),
            .I(N__20602));
    Span4Mux_h I__3490 (
            .O(N__20614),
            .I(N__20597));
    LocalMux I__3489 (
            .O(N__20611),
            .I(N__20597));
    CEMux I__3488 (
            .O(N__20610),
            .I(N__20583));
    Span4Mux_v I__3487 (
            .O(N__20607),
            .I(N__20580));
    InMux I__3486 (
            .O(N__20606),
            .I(N__20577));
    InMux I__3485 (
            .O(N__20605),
            .I(N__20574));
    LocalMux I__3484 (
            .O(N__20602),
            .I(N__20571));
    Span4Mux_v I__3483 (
            .O(N__20597),
            .I(N__20568));
    InMux I__3482 (
            .O(N__20596),
            .I(N__20559));
    InMux I__3481 (
            .O(N__20595),
            .I(N__20559));
    InMux I__3480 (
            .O(N__20594),
            .I(N__20559));
    InMux I__3479 (
            .O(N__20593),
            .I(N__20559));
    InMux I__3478 (
            .O(N__20592),
            .I(N__20550));
    InMux I__3477 (
            .O(N__20591),
            .I(N__20550));
    InMux I__3476 (
            .O(N__20590),
            .I(N__20550));
    InMux I__3475 (
            .O(N__20589),
            .I(N__20550));
    InMux I__3474 (
            .O(N__20588),
            .I(N__20547));
    InMux I__3473 (
            .O(N__20587),
            .I(N__20542));
    InMux I__3472 (
            .O(N__20586),
            .I(N__20542));
    LocalMux I__3471 (
            .O(N__20583),
            .I(N__20536));
    Span4Mux_v I__3470 (
            .O(N__20580),
            .I(N__20533));
    LocalMux I__3469 (
            .O(N__20577),
            .I(N__20530));
    LocalMux I__3468 (
            .O(N__20574),
            .I(N__20515));
    Span4Mux_h I__3467 (
            .O(N__20571),
            .I(N__20515));
    Span4Mux_s2_v I__3466 (
            .O(N__20568),
            .I(N__20515));
    LocalMux I__3465 (
            .O(N__20559),
            .I(N__20515));
    LocalMux I__3464 (
            .O(N__20550),
            .I(N__20515));
    LocalMux I__3463 (
            .O(N__20547),
            .I(N__20515));
    LocalMux I__3462 (
            .O(N__20542),
            .I(N__20515));
    InMux I__3461 (
            .O(N__20541),
            .I(N__20508));
    InMux I__3460 (
            .O(N__20540),
            .I(N__20508));
    InMux I__3459 (
            .O(N__20539),
            .I(N__20508));
    Span4Mux_v I__3458 (
            .O(N__20536),
            .I(N__20501));
    Span4Mux_h I__3457 (
            .O(N__20533),
            .I(N__20501));
    Span4Mux_v I__3456 (
            .O(N__20530),
            .I(N__20501));
    Sp12to4 I__3455 (
            .O(N__20515),
            .I(N__20496));
    LocalMux I__3454 (
            .O(N__20508),
            .I(N__20496));
    Odrv4 I__3453 (
            .O(N__20501),
            .I(\POWERLED.count_off_enZ0 ));
    Odrv12 I__3452 (
            .O(N__20496),
            .I(\POWERLED.count_off_enZ0 ));
    IoInMux I__3451 (
            .O(N__20491),
            .I(N__20488));
    LocalMux I__3450 (
            .O(N__20488),
            .I(N__20485));
    Odrv4 I__3449 (
            .O(N__20485),
            .I(G_10));
    InMux I__3448 (
            .O(N__20482),
            .I(N__20479));
    LocalMux I__3447 (
            .O(N__20479),
            .I(N__20476));
    Odrv4 I__3446 (
            .O(N__20476),
            .I(\POWERLED.un85_clk_100khz_11 ));
    CascadeMux I__3445 (
            .O(N__20473),
            .I(N__20470));
    InMux I__3444 (
            .O(N__20470),
            .I(N__20467));
    LocalMux I__3443 (
            .O(N__20467),
            .I(N__20464));
    Odrv4 I__3442 (
            .O(N__20464),
            .I(\POWERLED.un85_clk_100khz_10 ));
    InMux I__3441 (
            .O(N__20461),
            .I(N__20458));
    LocalMux I__3440 (
            .O(N__20458),
            .I(N__20454));
    InMux I__3439 (
            .O(N__20457),
            .I(N__20451));
    Odrv4 I__3438 (
            .O(N__20454),
            .I(\POWERLED.count_offZ0Z_12 ));
    LocalMux I__3437 (
            .O(N__20451),
            .I(\POWERLED.count_offZ0Z_12 ));
    InMux I__3436 (
            .O(N__20446),
            .I(N__20440));
    InMux I__3435 (
            .O(N__20445),
            .I(N__20440));
    LocalMux I__3434 (
            .O(N__20440),
            .I(N__20437));
    Odrv4 I__3433 (
            .O(N__20437),
            .I(\POWERLED.count_off_1_12 ));
    InMux I__3432 (
            .O(N__20434),
            .I(\POWERLED.un3_count_off_1_cry_11 ));
    InMux I__3431 (
            .O(N__20431),
            .I(N__20427));
    InMux I__3430 (
            .O(N__20430),
            .I(N__20424));
    LocalMux I__3429 (
            .O(N__20427),
            .I(\POWERLED.count_offZ0Z_13 ));
    LocalMux I__3428 (
            .O(N__20424),
            .I(\POWERLED.count_offZ0Z_13 ));
    InMux I__3427 (
            .O(N__20419),
            .I(N__20413));
    InMux I__3426 (
            .O(N__20418),
            .I(N__20413));
    LocalMux I__3425 (
            .O(N__20413),
            .I(\POWERLED.count_off_1_13 ));
    InMux I__3424 (
            .O(N__20410),
            .I(\POWERLED.un3_count_off_1_cry_12 ));
    InMux I__3423 (
            .O(N__20407),
            .I(N__20403));
    InMux I__3422 (
            .O(N__20406),
            .I(N__20400));
    LocalMux I__3421 (
            .O(N__20403),
            .I(\POWERLED.count_offZ0Z_14 ));
    LocalMux I__3420 (
            .O(N__20400),
            .I(\POWERLED.count_offZ0Z_14 ));
    InMux I__3419 (
            .O(N__20395),
            .I(N__20389));
    InMux I__3418 (
            .O(N__20394),
            .I(N__20389));
    LocalMux I__3417 (
            .O(N__20389),
            .I(\POWERLED.count_off_1_14 ));
    InMux I__3416 (
            .O(N__20386),
            .I(\POWERLED.un3_count_off_1_cry_13 ));
    InMux I__3415 (
            .O(N__20383),
            .I(N__20374));
    InMux I__3414 (
            .O(N__20382),
            .I(N__20374));
    InMux I__3413 (
            .O(N__20381),
            .I(N__20374));
    LocalMux I__3412 (
            .O(N__20374),
            .I(N__20361));
    InMux I__3411 (
            .O(N__20373),
            .I(N__20352));
    InMux I__3410 (
            .O(N__20372),
            .I(N__20352));
    InMux I__3409 (
            .O(N__20371),
            .I(N__20352));
    InMux I__3408 (
            .O(N__20370),
            .I(N__20352));
    InMux I__3407 (
            .O(N__20369),
            .I(N__20343));
    InMux I__3406 (
            .O(N__20368),
            .I(N__20343));
    InMux I__3405 (
            .O(N__20367),
            .I(N__20336));
    InMux I__3404 (
            .O(N__20366),
            .I(N__20336));
    InMux I__3403 (
            .O(N__20365),
            .I(N__20336));
    InMux I__3402 (
            .O(N__20364),
            .I(N__20333));
    Span4Mux_h I__3401 (
            .O(N__20361),
            .I(N__20327));
    LocalMux I__3400 (
            .O(N__20352),
            .I(N__20327));
    InMux I__3399 (
            .O(N__20351),
            .I(N__20317));
    InMux I__3398 (
            .O(N__20350),
            .I(N__20317));
    InMux I__3397 (
            .O(N__20349),
            .I(N__20317));
    InMux I__3396 (
            .O(N__20348),
            .I(N__20317));
    LocalMux I__3395 (
            .O(N__20343),
            .I(N__20312));
    LocalMux I__3394 (
            .O(N__20336),
            .I(N__20312));
    LocalMux I__3393 (
            .O(N__20333),
            .I(N__20309));
    InMux I__3392 (
            .O(N__20332),
            .I(N__20306));
    Span4Mux_v I__3391 (
            .O(N__20327),
            .I(N__20303));
    InMux I__3390 (
            .O(N__20326),
            .I(N__20300));
    LocalMux I__3389 (
            .O(N__20317),
            .I(N__20291));
    Span4Mux_h I__3388 (
            .O(N__20312),
            .I(N__20291));
    Span4Mux_v I__3387 (
            .O(N__20309),
            .I(N__20291));
    LocalMux I__3386 (
            .O(N__20306),
            .I(N__20291));
    Odrv4 I__3385 (
            .O(N__20303),
            .I(\POWERLED.N_96 ));
    LocalMux I__3384 (
            .O(N__20300),
            .I(\POWERLED.N_96 ));
    Odrv4 I__3383 (
            .O(N__20291),
            .I(\POWERLED.N_96 ));
    InMux I__3382 (
            .O(N__20284),
            .I(\POWERLED.un3_count_off_1_cry_14 ));
    InMux I__3381 (
            .O(N__20281),
            .I(N__20278));
    LocalMux I__3380 (
            .O(N__20278),
            .I(N__20274));
    InMux I__3379 (
            .O(N__20277),
            .I(N__20271));
    Odrv4 I__3378 (
            .O(N__20274),
            .I(\POWERLED.count_offZ0Z_9 ));
    LocalMux I__3377 (
            .O(N__20271),
            .I(\POWERLED.count_offZ0Z_9 ));
    InMux I__3376 (
            .O(N__20266),
            .I(N__20263));
    LocalMux I__3375 (
            .O(N__20263),
            .I(N__20259));
    InMux I__3374 (
            .O(N__20262),
            .I(N__20256));
    Odrv4 I__3373 (
            .O(N__20259),
            .I(\POWERLED.count_offZ0Z_15 ));
    LocalMux I__3372 (
            .O(N__20256),
            .I(\POWERLED.count_offZ0Z_15 ));
    InMux I__3371 (
            .O(N__20251),
            .I(N__20245));
    InMux I__3370 (
            .O(N__20250),
            .I(N__20245));
    LocalMux I__3369 (
            .O(N__20245),
            .I(\POWERLED.un3_count_off_1_cry_14_c_RNIMONZ0Z33 ));
    InMux I__3368 (
            .O(N__20242),
            .I(N__20239));
    LocalMux I__3367 (
            .O(N__20239),
            .I(\POWERLED.count_off_0_15 ));
    InMux I__3366 (
            .O(N__20236),
            .I(N__20233));
    LocalMux I__3365 (
            .O(N__20233),
            .I(N__20229));
    InMux I__3364 (
            .O(N__20232),
            .I(N__20226));
    Span4Mux_v I__3363 (
            .O(N__20229),
            .I(N__20221));
    LocalMux I__3362 (
            .O(N__20226),
            .I(N__20221));
    Odrv4 I__3361 (
            .O(N__20221),
            .I(\POWERLED.count_offZ0Z_7 ));
    InMux I__3360 (
            .O(N__20218),
            .I(N__20214));
    InMux I__3359 (
            .O(N__20217),
            .I(N__20211));
    LocalMux I__3358 (
            .O(N__20214),
            .I(N__20208));
    LocalMux I__3357 (
            .O(N__20211),
            .I(N__20205));
    Span4Mux_v I__3356 (
            .O(N__20208),
            .I(N__20202));
    Odrv4 I__3355 (
            .O(N__20205),
            .I(\POWERLED.count_offZ0Z_4 ));
    Odrv4 I__3354 (
            .O(N__20202),
            .I(\POWERLED.count_offZ0Z_4 ));
    InMux I__3353 (
            .O(N__20197),
            .I(N__20191));
    InMux I__3352 (
            .O(N__20196),
            .I(N__20191));
    LocalMux I__3351 (
            .O(N__20191),
            .I(N__20188));
    Span4Mux_h I__3350 (
            .O(N__20188),
            .I(N__20185));
    Odrv4 I__3349 (
            .O(N__20185),
            .I(\POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ));
    InMux I__3348 (
            .O(N__20182),
            .I(\POWERLED.un3_count_off_1_cry_3 ));
    InMux I__3347 (
            .O(N__20179),
            .I(N__20175));
    InMux I__3346 (
            .O(N__20178),
            .I(N__20172));
    LocalMux I__3345 (
            .O(N__20175),
            .I(N__20169));
    LocalMux I__3344 (
            .O(N__20172),
            .I(N__20166));
    Odrv4 I__3343 (
            .O(N__20169),
            .I(\POWERLED.count_offZ0Z_5 ));
    Odrv4 I__3342 (
            .O(N__20166),
            .I(\POWERLED.count_offZ0Z_5 ));
    InMux I__3341 (
            .O(N__20161),
            .I(N__20155));
    InMux I__3340 (
            .O(N__20160),
            .I(N__20155));
    LocalMux I__3339 (
            .O(N__20155),
            .I(N__20152));
    Odrv4 I__3338 (
            .O(N__20152),
            .I(\POWERLED.count_off_1_5 ));
    InMux I__3337 (
            .O(N__20149),
            .I(\POWERLED.un3_count_off_1_cry_4 ));
    CascadeMux I__3336 (
            .O(N__20146),
            .I(N__20143));
    InMux I__3335 (
            .O(N__20143),
            .I(N__20139));
    InMux I__3334 (
            .O(N__20142),
            .I(N__20136));
    LocalMux I__3333 (
            .O(N__20139),
            .I(N__20133));
    LocalMux I__3332 (
            .O(N__20136),
            .I(N__20130));
    Odrv12 I__3331 (
            .O(N__20133),
            .I(\POWERLED.count_offZ0Z_6 ));
    Odrv4 I__3330 (
            .O(N__20130),
            .I(\POWERLED.count_offZ0Z_6 ));
    InMux I__3329 (
            .O(N__20125),
            .I(N__20119));
    InMux I__3328 (
            .O(N__20124),
            .I(N__20119));
    LocalMux I__3327 (
            .O(N__20119),
            .I(N__20116));
    Odrv4 I__3326 (
            .O(N__20116),
            .I(\POWERLED.count_off_1_6 ));
    InMux I__3325 (
            .O(N__20113),
            .I(\POWERLED.un3_count_off_1_cry_5 ));
    InMux I__3324 (
            .O(N__20110),
            .I(\POWERLED.un3_count_off_1_cry_6 ));
    InMux I__3323 (
            .O(N__20107),
            .I(\POWERLED.un3_count_off_1_cry_7 ));
    InMux I__3322 (
            .O(N__20104),
            .I(bfn_6_13_0_));
    InMux I__3321 (
            .O(N__20101),
            .I(N__20098));
    LocalMux I__3320 (
            .O(N__20098),
            .I(N__20094));
    InMux I__3319 (
            .O(N__20097),
            .I(N__20091));
    Odrv4 I__3318 (
            .O(N__20094),
            .I(\POWERLED.count_offZ0Z_10 ));
    LocalMux I__3317 (
            .O(N__20091),
            .I(\POWERLED.count_offZ0Z_10 ));
    CascadeMux I__3316 (
            .O(N__20086),
            .I(N__20083));
    InMux I__3315 (
            .O(N__20083),
            .I(N__20077));
    InMux I__3314 (
            .O(N__20082),
            .I(N__20077));
    LocalMux I__3313 (
            .O(N__20077),
            .I(N__20074));
    Odrv4 I__3312 (
            .O(N__20074),
            .I(\POWERLED.count_off_1_10 ));
    InMux I__3311 (
            .O(N__20071),
            .I(\POWERLED.un3_count_off_1_cry_9 ));
    InMux I__3310 (
            .O(N__20068),
            .I(N__20064));
    CascadeMux I__3309 (
            .O(N__20067),
            .I(N__20061));
    LocalMux I__3308 (
            .O(N__20064),
            .I(N__20058));
    InMux I__3307 (
            .O(N__20061),
            .I(N__20055));
    Odrv4 I__3306 (
            .O(N__20058),
            .I(\POWERLED.count_offZ0Z_11 ));
    LocalMux I__3305 (
            .O(N__20055),
            .I(\POWERLED.count_offZ0Z_11 ));
    InMux I__3304 (
            .O(N__20050),
            .I(N__20044));
    InMux I__3303 (
            .O(N__20049),
            .I(N__20044));
    LocalMux I__3302 (
            .O(N__20044),
            .I(N__20041));
    Odrv4 I__3301 (
            .O(N__20041),
            .I(\POWERLED.count_off_1_11 ));
    InMux I__3300 (
            .O(N__20038),
            .I(\POWERLED.un3_count_off_1_cry_10 ));
    InMux I__3299 (
            .O(N__20035),
            .I(N__20032));
    LocalMux I__3298 (
            .O(N__20032),
            .I(\POWERLED.count_off_0_11 ));
    InMux I__3297 (
            .O(N__20029),
            .I(N__20026));
    LocalMux I__3296 (
            .O(N__20026),
            .I(\POWERLED.count_off_0_2 ));
    InMux I__3295 (
            .O(N__20023),
            .I(N__20020));
    LocalMux I__3294 (
            .O(N__20020),
            .I(\POWERLED.count_off_0_12 ));
    CascadeMux I__3293 (
            .O(N__20017),
            .I(N__20014));
    InMux I__3292 (
            .O(N__20014),
            .I(N__20008));
    InMux I__3291 (
            .O(N__20013),
            .I(N__20005));
    InMux I__3290 (
            .O(N__20012),
            .I(N__20002));
    InMux I__3289 (
            .O(N__20011),
            .I(N__19999));
    LocalMux I__3288 (
            .O(N__20008),
            .I(\POWERLED.count_offZ0Z_0 ));
    LocalMux I__3287 (
            .O(N__20005),
            .I(\POWERLED.count_offZ0Z_0 ));
    LocalMux I__3286 (
            .O(N__20002),
            .I(\POWERLED.count_offZ0Z_0 ));
    LocalMux I__3285 (
            .O(N__19999),
            .I(\POWERLED.count_offZ0Z_0 ));
    InMux I__3284 (
            .O(N__19990),
            .I(N__19986));
    CascadeMux I__3283 (
            .O(N__19989),
            .I(N__19982));
    LocalMux I__3282 (
            .O(N__19986),
            .I(N__19979));
    InMux I__3281 (
            .O(N__19985),
            .I(N__19976));
    InMux I__3280 (
            .O(N__19982),
            .I(N__19973));
    Odrv4 I__3279 (
            .O(N__19979),
            .I(\POWERLED.count_offZ0Z_1 ));
    LocalMux I__3278 (
            .O(N__19976),
            .I(\POWERLED.count_offZ0Z_1 ));
    LocalMux I__3277 (
            .O(N__19973),
            .I(\POWERLED.count_offZ0Z_1 ));
    InMux I__3276 (
            .O(N__19966),
            .I(N__19962));
    InMux I__3275 (
            .O(N__19965),
            .I(N__19959));
    LocalMux I__3274 (
            .O(N__19962),
            .I(\POWERLED.count_offZ0Z_2 ));
    LocalMux I__3273 (
            .O(N__19959),
            .I(\POWERLED.count_offZ0Z_2 ));
    InMux I__3272 (
            .O(N__19954),
            .I(N__19948));
    InMux I__3271 (
            .O(N__19953),
            .I(N__19948));
    LocalMux I__3270 (
            .O(N__19948),
            .I(\POWERLED.count_off_1_2 ));
    InMux I__3269 (
            .O(N__19945),
            .I(\POWERLED.un3_count_off_1_cry_1 ));
    CascadeMux I__3268 (
            .O(N__19942),
            .I(N__19939));
    InMux I__3267 (
            .O(N__19939),
            .I(N__19935));
    InMux I__3266 (
            .O(N__19938),
            .I(N__19932));
    LocalMux I__3265 (
            .O(N__19935),
            .I(\POWERLED.count_offZ0Z_3 ));
    LocalMux I__3264 (
            .O(N__19932),
            .I(\POWERLED.count_offZ0Z_3 ));
    InMux I__3263 (
            .O(N__19927),
            .I(N__19921));
    InMux I__3262 (
            .O(N__19926),
            .I(N__19921));
    LocalMux I__3261 (
            .O(N__19921),
            .I(\POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ));
    InMux I__3260 (
            .O(N__19918),
            .I(\POWERLED.un3_count_off_1_cry_2 ));
    CascadeMux I__3259 (
            .O(N__19915),
            .I(N__19912));
    InMux I__3258 (
            .O(N__19912),
            .I(N__19909));
    LocalMux I__3257 (
            .O(N__19909),
            .I(m3_1));
    InMux I__3256 (
            .O(N__19906),
            .I(N__19901));
    CascadeMux I__3255 (
            .O(N__19905),
            .I(N__19898));
    CascadeMux I__3254 (
            .O(N__19904),
            .I(N__19892));
    LocalMux I__3253 (
            .O(N__19901),
            .I(N__19883));
    InMux I__3252 (
            .O(N__19898),
            .I(N__19878));
    InMux I__3251 (
            .O(N__19897),
            .I(N__19878));
    InMux I__3250 (
            .O(N__19896),
            .I(N__19875));
    InMux I__3249 (
            .O(N__19895),
            .I(N__19872));
    InMux I__3248 (
            .O(N__19892),
            .I(N__19867));
    InMux I__3247 (
            .O(N__19891),
            .I(N__19867));
    InMux I__3246 (
            .O(N__19890),
            .I(N__19862));
    InMux I__3245 (
            .O(N__19889),
            .I(N__19862));
    InMux I__3244 (
            .O(N__19888),
            .I(N__19859));
    InMux I__3243 (
            .O(N__19887),
            .I(N__19854));
    InMux I__3242 (
            .O(N__19886),
            .I(N__19854));
    Span4Mux_v I__3241 (
            .O(N__19883),
            .I(N__19851));
    LocalMux I__3240 (
            .O(N__19878),
            .I(N__19848));
    LocalMux I__3239 (
            .O(N__19875),
            .I(N__19841));
    LocalMux I__3238 (
            .O(N__19872),
            .I(N__19841));
    LocalMux I__3237 (
            .O(N__19867),
            .I(N__19841));
    LocalMux I__3236 (
            .O(N__19862),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    LocalMux I__3235 (
            .O(N__19859),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    LocalMux I__3234 (
            .O(N__19854),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv4 I__3233 (
            .O(N__19851),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv4 I__3232 (
            .O(N__19848),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv4 I__3231 (
            .O(N__19841),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    InMux I__3230 (
            .O(N__19828),
            .I(N__19824));
    InMux I__3229 (
            .O(N__19827),
            .I(N__19821));
    LocalMux I__3228 (
            .O(N__19824),
            .I(\POWERLED.func_state_RNI5DLR_0Z0Z_0 ));
    LocalMux I__3227 (
            .O(N__19821),
            .I(\POWERLED.func_state_RNI5DLR_0Z0Z_0 ));
    InMux I__3226 (
            .O(N__19816),
            .I(N__19813));
    LocalMux I__3225 (
            .O(N__19813),
            .I(\POWERLED.func_state_1_m0_i_o2_2_1 ));
    InMux I__3224 (
            .O(N__19810),
            .I(N__19807));
    LocalMux I__3223 (
            .O(N__19807),
            .I(N__19803));
    InMux I__3222 (
            .O(N__19806),
            .I(N__19800));
    Span4Mux_v I__3221 (
            .O(N__19803),
            .I(N__19795));
    LocalMux I__3220 (
            .O(N__19800),
            .I(N__19795));
    Odrv4 I__3219 (
            .O(N__19795),
            .I(\POWERLED.func_state_RNILFRF4Z0Z_0 ));
    CascadeMux I__3218 (
            .O(N__19792),
            .I(\POWERLED.N_143_cascade_ ));
    InMux I__3217 (
            .O(N__19789),
            .I(N__19783));
    InMux I__3216 (
            .O(N__19788),
            .I(N__19783));
    LocalMux I__3215 (
            .O(N__19783),
            .I(\POWERLED.func_stateZ1Z_0 ));
    InMux I__3214 (
            .O(N__19780),
            .I(N__19774));
    InMux I__3213 (
            .O(N__19779),
            .I(N__19774));
    LocalMux I__3212 (
            .O(N__19774),
            .I(\POWERLED.func_state_RNIU8CJBZ0Z_0 ));
    CascadeMux I__3211 (
            .O(N__19771),
            .I(\POWERLED.func_stateZ0Z_0_cascade_ ));
    InMux I__3210 (
            .O(N__19768),
            .I(N__19765));
    LocalMux I__3209 (
            .O(N__19765),
            .I(\POWERLED.count_off_0_10 ));
    CascadeMux I__3208 (
            .O(N__19762),
            .I(\POWERLED.N_394_cascade_ ));
    InMux I__3207 (
            .O(N__19759),
            .I(N__19756));
    LocalMux I__3206 (
            .O(N__19756),
            .I(N__19753));
    Odrv4 I__3205 (
            .O(N__19753),
            .I(\POWERLED.N_453 ));
    InMux I__3204 (
            .O(N__19750),
            .I(N__19744));
    InMux I__3203 (
            .O(N__19749),
            .I(N__19744));
    LocalMux I__3202 (
            .O(N__19744),
            .I(N__19741));
    Span4Mux_v I__3201 (
            .O(N__19741),
            .I(N__19737));
    InMux I__3200 (
            .O(N__19740),
            .I(N__19734));
    Odrv4 I__3199 (
            .O(N__19737),
            .I(\POWERLED.func_state_RNI5DLR_1Z0Z_1 ));
    LocalMux I__3198 (
            .O(N__19734),
            .I(\POWERLED.func_state_RNI5DLR_1Z0Z_1 ));
    CascadeMux I__3197 (
            .O(N__19729),
            .I(\POWERLED.un1_func_state25_6_0_0_a3_0_cascade_ ));
    InMux I__3196 (
            .O(N__19726),
            .I(N__19723));
    LocalMux I__3195 (
            .O(N__19723),
            .I(\POWERLED.un1_func_state25_6_0_o_N_422_N ));
    InMux I__3194 (
            .O(N__19720),
            .I(N__19716));
    InMux I__3193 (
            .O(N__19719),
            .I(N__19713));
    LocalMux I__3192 (
            .O(N__19716),
            .I(\POWERLED.un1_func_state25_6_0_o_N_516_N ));
    LocalMux I__3191 (
            .O(N__19713),
            .I(\POWERLED.un1_func_state25_6_0_o_N_516_N ));
    InMux I__3190 (
            .O(N__19708),
            .I(N__19705));
    LocalMux I__3189 (
            .O(N__19705),
            .I(\POWERLED.un1_func_state25_6_0_o_N_425_N ));
    InMux I__3188 (
            .O(N__19702),
            .I(N__19699));
    LocalMux I__3187 (
            .O(N__19699),
            .I(\POWERLED.un1_func_state25_6_0_0_2 ));
    CascadeMux I__3186 (
            .O(N__19696),
            .I(N__19693));
    InMux I__3185 (
            .O(N__19693),
            .I(N__19690));
    LocalMux I__3184 (
            .O(N__19690),
            .I(\POWERLED.un1_func_state25_6_0_0_0 ));
    CascadeMux I__3183 (
            .O(N__19687),
            .I(\POWERLED.N_341_cascade_ ));
    CascadeMux I__3182 (
            .O(N__19684),
            .I(N__19681));
    InMux I__3181 (
            .O(N__19681),
            .I(N__19678));
    LocalMux I__3180 (
            .O(N__19678),
            .I(\POWERLED.mult1_un159_sum_cry_2_s ));
    InMux I__3179 (
            .O(N__19675),
            .I(N__19672));
    LocalMux I__3178 (
            .O(N__19672),
            .I(\POWERLED.mult1_un159_sum_cry_3_s ));
    InMux I__3177 (
            .O(N__19669),
            .I(N__19666));
    LocalMux I__3176 (
            .O(N__19666),
            .I(\POWERLED.mult1_un159_sum_cry_4_s ));
    InMux I__3175 (
            .O(N__19663),
            .I(N__19660));
    LocalMux I__3174 (
            .O(N__19660),
            .I(\POWERLED.mult1_un159_sum_cry_5_s ));
    CascadeMux I__3173 (
            .O(N__19657),
            .I(N__19653));
    CascadeMux I__3172 (
            .O(N__19656),
            .I(N__19649));
    InMux I__3171 (
            .O(N__19653),
            .I(N__19642));
    InMux I__3170 (
            .O(N__19652),
            .I(N__19642));
    InMux I__3169 (
            .O(N__19649),
            .I(N__19642));
    LocalMux I__3168 (
            .O(N__19642),
            .I(N__19639));
    Odrv4 I__3167 (
            .O(N__19639),
            .I(G_2129));
    InMux I__3166 (
            .O(N__19636),
            .I(N__19633));
    LocalMux I__3165 (
            .O(N__19633),
            .I(\POWERLED.mult1_un166_sum_axb_6 ));
    InMux I__3164 (
            .O(N__19630),
            .I(\POWERLED.mult1_un166_sum_cry_5 ));
    CascadeMux I__3163 (
            .O(N__19627),
            .I(N__19624));
    InMux I__3162 (
            .O(N__19624),
            .I(N__19621));
    LocalMux I__3161 (
            .O(N__19621),
            .I(N__19618));
    Odrv12 I__3160 (
            .O(N__19618),
            .I(\POWERLED.un85_clk_100khz_0 ));
    CascadeMux I__3159 (
            .O(N__19615),
            .I(N__19611));
    CascadeMux I__3158 (
            .O(N__19614),
            .I(N__19607));
    InMux I__3157 (
            .O(N__19611),
            .I(N__19602));
    InMux I__3156 (
            .O(N__19610),
            .I(N__19599));
    InMux I__3155 (
            .O(N__19607),
            .I(N__19592));
    InMux I__3154 (
            .O(N__19606),
            .I(N__19592));
    InMux I__3153 (
            .O(N__19605),
            .I(N__19592));
    LocalMux I__3152 (
            .O(N__19602),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__3151 (
            .O(N__19599),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__3150 (
            .O(N__19592),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    CascadeMux I__3149 (
            .O(N__19585),
            .I(N__19582));
    InMux I__3148 (
            .O(N__19582),
            .I(N__19579));
    LocalMux I__3147 (
            .O(N__19579),
            .I(N__19576));
    Span12Mux_s2_v I__3146 (
            .O(N__19576),
            .I(N__19573));
    Odrv12 I__3145 (
            .O(N__19573),
            .I(\POWERLED.un85_clk_100khz_1 ));
    InMux I__3144 (
            .O(N__19570),
            .I(N__19567));
    LocalMux I__3143 (
            .O(N__19567),
            .I(\POWERLED.mult1_un117_sum_cry_5_s ));
    InMux I__3142 (
            .O(N__19564),
            .I(\POWERLED.mult1_un117_sum_cry_4 ));
    InMux I__3141 (
            .O(N__19561),
            .I(N__19555));
    InMux I__3140 (
            .O(N__19560),
            .I(N__19555));
    LocalMux I__3139 (
            .O(N__19555),
            .I(\POWERLED.mult1_un117_sum_cry_6_s ));
    InMux I__3138 (
            .O(N__19552),
            .I(\POWERLED.mult1_un117_sum_cry_5 ));
    CascadeMux I__3137 (
            .O(N__19549),
            .I(N__19545));
    CascadeMux I__3136 (
            .O(N__19548),
            .I(N__19541));
    InMux I__3135 (
            .O(N__19545),
            .I(N__19534));
    InMux I__3134 (
            .O(N__19544),
            .I(N__19534));
    InMux I__3133 (
            .O(N__19541),
            .I(N__19534));
    LocalMux I__3132 (
            .O(N__19534),
            .I(\POWERLED.mult1_un110_sum_i_0_8 ));
    CascadeMux I__3131 (
            .O(N__19531),
            .I(N__19528));
    InMux I__3130 (
            .O(N__19528),
            .I(N__19525));
    LocalMux I__3129 (
            .O(N__19525),
            .I(\POWERLED.mult1_un124_sum_axb_8 ));
    InMux I__3128 (
            .O(N__19522),
            .I(\POWERLED.mult1_un117_sum_cry_6 ));
    InMux I__3127 (
            .O(N__19519),
            .I(\POWERLED.mult1_un117_sum_cry_7 ));
    InMux I__3126 (
            .O(N__19516),
            .I(N__19512));
    InMux I__3125 (
            .O(N__19515),
            .I(N__19509));
    LocalMux I__3124 (
            .O(N__19512),
            .I(\POWERLED.mult1_un117_sum_cry_3_s ));
    LocalMux I__3123 (
            .O(N__19509),
            .I(\POWERLED.mult1_un117_sum_cry_3_s ));
    CascadeMux I__3122 (
            .O(N__19504),
            .I(\POWERLED.mult1_un117_sum_s_8_cascade_ ));
    CascadeMux I__3121 (
            .O(N__19501),
            .I(N__19498));
    InMux I__3120 (
            .O(N__19498),
            .I(N__19495));
    LocalMux I__3119 (
            .O(N__19495),
            .I(\POWERLED.mult1_un124_sum_axb_4_l_fx ));
    InMux I__3118 (
            .O(N__19492),
            .I(N__19489));
    LocalMux I__3117 (
            .O(N__19489),
            .I(N__19486));
    Span4Mux_h I__3116 (
            .O(N__19486),
            .I(N__19483));
    Odrv4 I__3115 (
            .O(N__19483),
            .I(\PCH_PWRGD.N_38_f0 ));
    InMux I__3114 (
            .O(N__19480),
            .I(N__19474));
    InMux I__3113 (
            .O(N__19479),
            .I(N__19471));
    InMux I__3112 (
            .O(N__19478),
            .I(N__19466));
    InMux I__3111 (
            .O(N__19477),
            .I(N__19466));
    LocalMux I__3110 (
            .O(N__19474),
            .I(N__19463));
    LocalMux I__3109 (
            .O(N__19471),
            .I(N__19460));
    LocalMux I__3108 (
            .O(N__19466),
            .I(N__19457));
    Span4Mux_v I__3107 (
            .O(N__19463),
            .I(N__19454));
    Span4Mux_s3_h I__3106 (
            .O(N__19460),
            .I(N__19451));
    Span12Mux_s3_h I__3105 (
            .O(N__19457),
            .I(N__19448));
    Odrv4 I__3104 (
            .O(N__19454),
            .I(\PCH_PWRGD.curr_state_0_sqmuxa ));
    Odrv4 I__3103 (
            .O(N__19451),
            .I(\PCH_PWRGD.curr_state_0_sqmuxa ));
    Odrv12 I__3102 (
            .O(N__19448),
            .I(\PCH_PWRGD.curr_state_0_sqmuxa ));
    InMux I__3101 (
            .O(N__19441),
            .I(N__19438));
    LocalMux I__3100 (
            .O(N__19438),
            .I(N__19434));
    InMux I__3099 (
            .O(N__19437),
            .I(N__19431));
    Span12Mux_s6_v I__3098 (
            .O(N__19434),
            .I(N__19428));
    LocalMux I__3097 (
            .O(N__19431),
            .I(\PCH_PWRGD.delayed_vccin_ok_0 ));
    Odrv12 I__3096 (
            .O(N__19428),
            .I(\PCH_PWRGD.delayed_vccin_ok_0 ));
    CascadeMux I__3095 (
            .O(N__19423),
            .I(N__19418));
    InMux I__3094 (
            .O(N__19422),
            .I(N__19412));
    InMux I__3093 (
            .O(N__19421),
            .I(N__19409));
    InMux I__3092 (
            .O(N__19418),
            .I(N__19402));
    InMux I__3091 (
            .O(N__19417),
            .I(N__19402));
    InMux I__3090 (
            .O(N__19416),
            .I(N__19402));
    InMux I__3089 (
            .O(N__19415),
            .I(N__19399));
    LocalMux I__3088 (
            .O(N__19412),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__3087 (
            .O(N__19409),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__3086 (
            .O(N__19402),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__3085 (
            .O(N__19399),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    CascadeMux I__3084 (
            .O(N__19390),
            .I(N__19387));
    InMux I__3083 (
            .O(N__19387),
            .I(N__19384));
    LocalMux I__3082 (
            .O(N__19384),
            .I(\POWERLED.mult1_un117_sum_i_0_8 ));
    InMux I__3081 (
            .O(N__19381),
            .I(N__19378));
    LocalMux I__3080 (
            .O(N__19378),
            .I(N__19375));
    Odrv4 I__3079 (
            .O(N__19375),
            .I(\POWERLED.un85_clk_100khz_7 ));
    InMux I__3078 (
            .O(N__19372),
            .I(N__19369));
    LocalMux I__3077 (
            .O(N__19369),
            .I(N__19366));
    Odrv12 I__3076 (
            .O(N__19366),
            .I(\POWERLED.mult1_un131_sum_i ));
    InMux I__3075 (
            .O(N__19363),
            .I(N__19360));
    LocalMux I__3074 (
            .O(N__19360),
            .I(\POWERLED.mult1_un138_sum_i ));
    InMux I__3073 (
            .O(N__19357),
            .I(N__19354));
    LocalMux I__3072 (
            .O(N__19354),
            .I(\POWERLED.mult1_un117_sum_i ));
    InMux I__3071 (
            .O(N__19351),
            .I(N__19348));
    LocalMux I__3070 (
            .O(N__19348),
            .I(N__19345));
    Span12Mux_s11_v I__3069 (
            .O(N__19345),
            .I(N__19342));
    Odrv12 I__3068 (
            .O(N__19342),
            .I(\POWERLED.mult1_un124_sum_i ));
    InMux I__3067 (
            .O(N__19339),
            .I(N__19336));
    LocalMux I__3066 (
            .O(N__19336),
            .I(\POWERLED.mult1_un110_sum_i ));
    InMux I__3065 (
            .O(N__19333),
            .I(\POWERLED.mult1_un117_sum_cry_2 ));
    CascadeMux I__3064 (
            .O(N__19330),
            .I(N__19327));
    InMux I__3063 (
            .O(N__19327),
            .I(N__19324));
    LocalMux I__3062 (
            .O(N__19324),
            .I(\POWERLED.mult1_un117_sum_cry_4_s ));
    InMux I__3061 (
            .O(N__19321),
            .I(\POWERLED.mult1_un117_sum_cry_3 ));
    InMux I__3060 (
            .O(N__19318),
            .I(N__19314));
    InMux I__3059 (
            .O(N__19317),
            .I(N__19310));
    LocalMux I__3058 (
            .O(N__19314),
            .I(N__19307));
    InMux I__3057 (
            .O(N__19313),
            .I(N__19304));
    LocalMux I__3056 (
            .O(N__19310),
            .I(\POWERLED.countZ0Z_9 ));
    Odrv4 I__3055 (
            .O(N__19307),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__3054 (
            .O(N__19304),
            .I(\POWERLED.countZ0Z_9 ));
    CascadeMux I__3053 (
            .O(N__19297),
            .I(N__19294));
    InMux I__3052 (
            .O(N__19294),
            .I(N__19291));
    LocalMux I__3051 (
            .O(N__19291),
            .I(\POWERLED.N_4706_i ));
    InMux I__3050 (
            .O(N__19288),
            .I(N__19283));
    InMux I__3049 (
            .O(N__19287),
            .I(N__19280));
    InMux I__3048 (
            .O(N__19286),
            .I(N__19277));
    LocalMux I__3047 (
            .O(N__19283),
            .I(N__19274));
    LocalMux I__3046 (
            .O(N__19280),
            .I(\POWERLED.countZ0Z_10 ));
    LocalMux I__3045 (
            .O(N__19277),
            .I(\POWERLED.countZ0Z_10 ));
    Odrv12 I__3044 (
            .O(N__19274),
            .I(\POWERLED.countZ0Z_10 ));
    InMux I__3043 (
            .O(N__19267),
            .I(N__19264));
    LocalMux I__3042 (
            .O(N__19264),
            .I(\POWERLED.N_4707_i ));
    InMux I__3041 (
            .O(N__19261),
            .I(N__19256));
    InMux I__3040 (
            .O(N__19260),
            .I(N__19253));
    InMux I__3039 (
            .O(N__19259),
            .I(N__19250));
    LocalMux I__3038 (
            .O(N__19256),
            .I(N__19247));
    LocalMux I__3037 (
            .O(N__19253),
            .I(N__19244));
    LocalMux I__3036 (
            .O(N__19250),
            .I(\POWERLED.countZ0Z_11 ));
    Odrv4 I__3035 (
            .O(N__19247),
            .I(\POWERLED.countZ0Z_11 ));
    Odrv4 I__3034 (
            .O(N__19244),
            .I(\POWERLED.countZ0Z_11 ));
    CascadeMux I__3033 (
            .O(N__19237),
            .I(N__19234));
    InMux I__3032 (
            .O(N__19234),
            .I(N__19231));
    LocalMux I__3031 (
            .O(N__19231),
            .I(\POWERLED.N_4708_i ));
    InMux I__3030 (
            .O(N__19228),
            .I(N__19225));
    LocalMux I__3029 (
            .O(N__19225),
            .I(N__19221));
    CascadeMux I__3028 (
            .O(N__19224),
            .I(N__19217));
    Span4Mux_v I__3027 (
            .O(N__19221),
            .I(N__19214));
    InMux I__3026 (
            .O(N__19220),
            .I(N__19211));
    InMux I__3025 (
            .O(N__19217),
            .I(N__19208));
    Odrv4 I__3024 (
            .O(N__19214),
            .I(\POWERLED.countZ0Z_12 ));
    LocalMux I__3023 (
            .O(N__19211),
            .I(\POWERLED.countZ0Z_12 ));
    LocalMux I__3022 (
            .O(N__19208),
            .I(\POWERLED.countZ0Z_12 ));
    CascadeMux I__3021 (
            .O(N__19201),
            .I(N__19198));
    InMux I__3020 (
            .O(N__19198),
            .I(N__19195));
    LocalMux I__3019 (
            .O(N__19195),
            .I(\POWERLED.N_4709_i ));
    InMux I__3018 (
            .O(N__19192),
            .I(N__19189));
    LocalMux I__3017 (
            .O(N__19189),
            .I(N__19185));
    InMux I__3016 (
            .O(N__19188),
            .I(N__19182));
    Span4Mux_v I__3015 (
            .O(N__19185),
            .I(N__19178));
    LocalMux I__3014 (
            .O(N__19182),
            .I(N__19175));
    InMux I__3013 (
            .O(N__19181),
            .I(N__19172));
    Odrv4 I__3012 (
            .O(N__19178),
            .I(\POWERLED.countZ0Z_13 ));
    Odrv4 I__3011 (
            .O(N__19175),
            .I(\POWERLED.countZ0Z_13 ));
    LocalMux I__3010 (
            .O(N__19172),
            .I(\POWERLED.countZ0Z_13 ));
    InMux I__3009 (
            .O(N__19165),
            .I(N__19162));
    LocalMux I__3008 (
            .O(N__19162),
            .I(\POWERLED.N_4710_i ));
    InMux I__3007 (
            .O(N__19159),
            .I(N__19156));
    LocalMux I__3006 (
            .O(N__19156),
            .I(N__19152));
    InMux I__3005 (
            .O(N__19155),
            .I(N__19149));
    Span4Mux_h I__3004 (
            .O(N__19152),
            .I(N__19143));
    LocalMux I__3003 (
            .O(N__19149),
            .I(N__19143));
    InMux I__3002 (
            .O(N__19148),
            .I(N__19140));
    Odrv4 I__3001 (
            .O(N__19143),
            .I(\POWERLED.countZ0Z_14 ));
    LocalMux I__3000 (
            .O(N__19140),
            .I(\POWERLED.countZ0Z_14 ));
    CascadeMux I__2999 (
            .O(N__19135),
            .I(N__19132));
    InMux I__2998 (
            .O(N__19132),
            .I(N__19129));
    LocalMux I__2997 (
            .O(N__19129),
            .I(\POWERLED.N_4711_i ));
    InMux I__2996 (
            .O(N__19126),
            .I(N__19122));
    InMux I__2995 (
            .O(N__19125),
            .I(N__19119));
    LocalMux I__2994 (
            .O(N__19122),
            .I(N__19115));
    LocalMux I__2993 (
            .O(N__19119),
            .I(N__19112));
    InMux I__2992 (
            .O(N__19118),
            .I(N__19109));
    Odrv4 I__2991 (
            .O(N__19115),
            .I(\POWERLED.countZ0Z_15 ));
    Odrv12 I__2990 (
            .O(N__19112),
            .I(\POWERLED.countZ0Z_15 ));
    LocalMux I__2989 (
            .O(N__19109),
            .I(\POWERLED.countZ0Z_15 ));
    CascadeMux I__2988 (
            .O(N__19102),
            .I(N__19099));
    InMux I__2987 (
            .O(N__19099),
            .I(N__19096));
    LocalMux I__2986 (
            .O(N__19096),
            .I(N__19093));
    Odrv4 I__2985 (
            .O(N__19093),
            .I(\POWERLED.N_4712_i ));
    InMux I__2984 (
            .O(N__19090),
            .I(bfn_6_5_0_));
    CascadeMux I__2983 (
            .O(N__19087),
            .I(N__19084));
    InMux I__2982 (
            .O(N__19084),
            .I(N__19081));
    LocalMux I__2981 (
            .O(N__19081),
            .I(\POWERLED.un85_clk_100khz_2 ));
    InMux I__2980 (
            .O(N__19078),
            .I(N__19073));
    InMux I__2979 (
            .O(N__19077),
            .I(N__19070));
    InMux I__2978 (
            .O(N__19076),
            .I(N__19067));
    LocalMux I__2977 (
            .O(N__19073),
            .I(\POWERLED.countZ0Z_2 ));
    LocalMux I__2976 (
            .O(N__19070),
            .I(\POWERLED.countZ0Z_2 ));
    LocalMux I__2975 (
            .O(N__19067),
            .I(\POWERLED.countZ0Z_2 ));
    InMux I__2974 (
            .O(N__19060),
            .I(N__19057));
    LocalMux I__2973 (
            .O(N__19057),
            .I(\POWERLED.N_4699_i ));
    InMux I__2972 (
            .O(N__19054),
            .I(N__19051));
    LocalMux I__2971 (
            .O(N__19051),
            .I(N__19047));
    InMux I__2970 (
            .O(N__19050),
            .I(N__19044));
    Span4Mux_v I__2969 (
            .O(N__19047),
            .I(N__19040));
    LocalMux I__2968 (
            .O(N__19044),
            .I(N__19037));
    InMux I__2967 (
            .O(N__19043),
            .I(N__19034));
    Odrv4 I__2966 (
            .O(N__19040),
            .I(\POWERLED.countZ0Z_3 ));
    Odrv12 I__2965 (
            .O(N__19037),
            .I(\POWERLED.countZ0Z_3 ));
    LocalMux I__2964 (
            .O(N__19034),
            .I(\POWERLED.countZ0Z_3 ));
    InMux I__2963 (
            .O(N__19027),
            .I(N__19024));
    LocalMux I__2962 (
            .O(N__19024),
            .I(\POWERLED.un85_clk_100khz_3 ));
    CascadeMux I__2961 (
            .O(N__19021),
            .I(N__19018));
    InMux I__2960 (
            .O(N__19018),
            .I(N__19015));
    LocalMux I__2959 (
            .O(N__19015),
            .I(\POWERLED.N_4700_i ));
    CascadeMux I__2958 (
            .O(N__19012),
            .I(N__19007));
    InMux I__2957 (
            .O(N__19011),
            .I(N__19004));
    InMux I__2956 (
            .O(N__19010),
            .I(N__19001));
    InMux I__2955 (
            .O(N__19007),
            .I(N__18998));
    LocalMux I__2954 (
            .O(N__19004),
            .I(N__18995));
    LocalMux I__2953 (
            .O(N__19001),
            .I(N__18990));
    LocalMux I__2952 (
            .O(N__18998),
            .I(N__18990));
    Odrv12 I__2951 (
            .O(N__18995),
            .I(\POWERLED.countZ0Z_4 ));
    Odrv4 I__2950 (
            .O(N__18990),
            .I(\POWERLED.countZ0Z_4 ));
    InMux I__2949 (
            .O(N__18985),
            .I(N__18982));
    LocalMux I__2948 (
            .O(N__18982),
            .I(\POWERLED.un85_clk_100khz_4 ));
    CascadeMux I__2947 (
            .O(N__18979),
            .I(N__18976));
    InMux I__2946 (
            .O(N__18976),
            .I(N__18973));
    LocalMux I__2945 (
            .O(N__18973),
            .I(\POWERLED.N_4701_i ));
    InMux I__2944 (
            .O(N__18970),
            .I(N__18967));
    LocalMux I__2943 (
            .O(N__18967),
            .I(\POWERLED.un85_clk_100khz_5 ));
    InMux I__2942 (
            .O(N__18964),
            .I(N__18961));
    LocalMux I__2941 (
            .O(N__18961),
            .I(N__18956));
    InMux I__2940 (
            .O(N__18960),
            .I(N__18953));
    InMux I__2939 (
            .O(N__18959),
            .I(N__18950));
    Span4Mux_s2_v I__2938 (
            .O(N__18956),
            .I(N__18947));
    LocalMux I__2937 (
            .O(N__18953),
            .I(N__18944));
    LocalMux I__2936 (
            .O(N__18950),
            .I(\POWERLED.countZ0Z_5 ));
    Odrv4 I__2935 (
            .O(N__18947),
            .I(\POWERLED.countZ0Z_5 ));
    Odrv4 I__2934 (
            .O(N__18944),
            .I(\POWERLED.countZ0Z_5 ));
    CascadeMux I__2933 (
            .O(N__18937),
            .I(N__18934));
    InMux I__2932 (
            .O(N__18934),
            .I(N__18931));
    LocalMux I__2931 (
            .O(N__18931),
            .I(\POWERLED.N_4702_i ));
    CascadeMux I__2930 (
            .O(N__18928),
            .I(N__18925));
    InMux I__2929 (
            .O(N__18925),
            .I(N__18922));
    LocalMux I__2928 (
            .O(N__18922),
            .I(\POWERLED.un85_clk_100khz_6 ));
    InMux I__2927 (
            .O(N__18919),
            .I(N__18915));
    InMux I__2926 (
            .O(N__18918),
            .I(N__18911));
    LocalMux I__2925 (
            .O(N__18915),
            .I(N__18908));
    InMux I__2924 (
            .O(N__18914),
            .I(N__18905));
    LocalMux I__2923 (
            .O(N__18911),
            .I(\POWERLED.countZ0Z_6 ));
    Odrv4 I__2922 (
            .O(N__18908),
            .I(\POWERLED.countZ0Z_6 ));
    LocalMux I__2921 (
            .O(N__18905),
            .I(\POWERLED.countZ0Z_6 ));
    InMux I__2920 (
            .O(N__18898),
            .I(N__18895));
    LocalMux I__2919 (
            .O(N__18895),
            .I(\POWERLED.N_4703_i ));
    InMux I__2918 (
            .O(N__18892),
            .I(N__18889));
    LocalMux I__2917 (
            .O(N__18889),
            .I(N__18884));
    InMux I__2916 (
            .O(N__18888),
            .I(N__18881));
    InMux I__2915 (
            .O(N__18887),
            .I(N__18878));
    Span4Mux_h I__2914 (
            .O(N__18884),
            .I(N__18873));
    LocalMux I__2913 (
            .O(N__18881),
            .I(N__18873));
    LocalMux I__2912 (
            .O(N__18878),
            .I(\POWERLED.countZ0Z_7 ));
    Odrv4 I__2911 (
            .O(N__18873),
            .I(\POWERLED.countZ0Z_7 ));
    CascadeMux I__2910 (
            .O(N__18868),
            .I(N__18865));
    InMux I__2909 (
            .O(N__18865),
            .I(N__18862));
    LocalMux I__2908 (
            .O(N__18862),
            .I(\POWERLED.N_4704_i ));
    InMux I__2907 (
            .O(N__18859),
            .I(N__18856));
    LocalMux I__2906 (
            .O(N__18856),
            .I(N__18853));
    Sp12to4 I__2905 (
            .O(N__18853),
            .I(N__18848));
    InMux I__2904 (
            .O(N__18852),
            .I(N__18845));
    InMux I__2903 (
            .O(N__18851),
            .I(N__18842));
    Odrv12 I__2902 (
            .O(N__18848),
            .I(\POWERLED.countZ0Z_8 ));
    LocalMux I__2901 (
            .O(N__18845),
            .I(\POWERLED.countZ0Z_8 ));
    LocalMux I__2900 (
            .O(N__18842),
            .I(\POWERLED.countZ0Z_8 ));
    CascadeMux I__2899 (
            .O(N__18835),
            .I(N__18832));
    InMux I__2898 (
            .O(N__18832),
            .I(N__18829));
    LocalMux I__2897 (
            .O(N__18829),
            .I(\POWERLED.N_4705_i ));
    CascadeMux I__2896 (
            .O(N__18826),
            .I(N__18823));
    InMux I__2895 (
            .O(N__18823),
            .I(N__18817));
    InMux I__2894 (
            .O(N__18822),
            .I(N__18817));
    LocalMux I__2893 (
            .O(N__18817),
            .I(\POWERLED.un1_count_cry_8_c_RNIIGZ0Z79 ));
    InMux I__2892 (
            .O(N__18814),
            .I(N__18811));
    LocalMux I__2891 (
            .O(N__18811),
            .I(\POWERLED.count_0_9 ));
    InMux I__2890 (
            .O(N__18808),
            .I(N__18804));
    InMux I__2889 (
            .O(N__18807),
            .I(N__18801));
    LocalMux I__2888 (
            .O(N__18804),
            .I(\POWERLED.un1_count_cry_9_c_RNIJIZ0Z89 ));
    LocalMux I__2887 (
            .O(N__18801),
            .I(\POWERLED.un1_count_cry_9_c_RNIJIZ0Z89 ));
    InMux I__2886 (
            .O(N__18796),
            .I(N__18793));
    LocalMux I__2885 (
            .O(N__18793),
            .I(\POWERLED.count_0_10 ));
    CascadeMux I__2884 (
            .O(N__18790),
            .I(N__18786));
    InMux I__2883 (
            .O(N__18789),
            .I(N__18781));
    InMux I__2882 (
            .O(N__18786),
            .I(N__18781));
    LocalMux I__2881 (
            .O(N__18781),
            .I(\POWERLED.un1_count_cry_1_c_RNIBZ0Z209 ));
    InMux I__2880 (
            .O(N__18778),
            .I(N__18775));
    LocalMux I__2879 (
            .O(N__18775),
            .I(\POWERLED.count_0_2 ));
    InMux I__2878 (
            .O(N__18772),
            .I(N__18768));
    InMux I__2877 (
            .O(N__18771),
            .I(N__18765));
    LocalMux I__2876 (
            .O(N__18768),
            .I(\POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7 ));
    LocalMux I__2875 (
            .O(N__18765),
            .I(\POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7 ));
    InMux I__2874 (
            .O(N__18760),
            .I(N__18757));
    LocalMux I__2873 (
            .O(N__18757),
            .I(\POWERLED.count_0_11 ));
    InMux I__2872 (
            .O(N__18754),
            .I(N__18751));
    LocalMux I__2871 (
            .O(N__18751),
            .I(N__18747));
    CascadeMux I__2870 (
            .O(N__18750),
            .I(N__18740));
    Span4Mux_v I__2869 (
            .O(N__18747),
            .I(N__18737));
    InMux I__2868 (
            .O(N__18746),
            .I(N__18734));
    InMux I__2867 (
            .O(N__18745),
            .I(N__18727));
    InMux I__2866 (
            .O(N__18744),
            .I(N__18727));
    InMux I__2865 (
            .O(N__18743),
            .I(N__18727));
    InMux I__2864 (
            .O(N__18740),
            .I(N__18724));
    Odrv4 I__2863 (
            .O(N__18737),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__2862 (
            .O(N__18734),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__2861 (
            .O(N__18727),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__2860 (
            .O(N__18724),
            .I(\POWERLED.countZ0Z_0 ));
    InMux I__2859 (
            .O(N__18715),
            .I(N__18712));
    LocalMux I__2858 (
            .O(N__18712),
            .I(\POWERLED.un1_count_cry_0_i ));
    InMux I__2857 (
            .O(N__18709),
            .I(N__18706));
    LocalMux I__2856 (
            .O(N__18706),
            .I(N__18703));
    Span4Mux_v I__2855 (
            .O(N__18703),
            .I(N__18698));
    InMux I__2854 (
            .O(N__18702),
            .I(N__18695));
    InMux I__2853 (
            .O(N__18701),
            .I(N__18692));
    Odrv4 I__2852 (
            .O(N__18698),
            .I(\POWERLED.countZ0Z_1 ));
    LocalMux I__2851 (
            .O(N__18695),
            .I(\POWERLED.countZ0Z_1 ));
    LocalMux I__2850 (
            .O(N__18692),
            .I(\POWERLED.countZ0Z_1 ));
    InMux I__2849 (
            .O(N__18685),
            .I(N__18682));
    LocalMux I__2848 (
            .O(N__18682),
            .I(\POWERLED.N_4698_i ));
    CascadeMux I__2847 (
            .O(N__18679),
            .I(N__18675));
    InMux I__2846 (
            .O(N__18678),
            .I(N__18670));
    InMux I__2845 (
            .O(N__18675),
            .I(N__18670));
    LocalMux I__2844 (
            .O(N__18670),
            .I(\POWERLED.un1_count_cry_5_c_RNIFAZ0Z49 ));
    InMux I__2843 (
            .O(N__18667),
            .I(N__18664));
    LocalMux I__2842 (
            .O(N__18664),
            .I(\POWERLED.count_0_6 ));
    CascadeMux I__2841 (
            .O(N__18661),
            .I(N__18658));
    InMux I__2840 (
            .O(N__18658),
            .I(N__18652));
    InMux I__2839 (
            .O(N__18657),
            .I(N__18652));
    LocalMux I__2838 (
            .O(N__18652),
            .I(N__18649));
    Odrv4 I__2837 (
            .O(N__18649),
            .I(\POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ));
    InMux I__2836 (
            .O(N__18646),
            .I(N__18643));
    LocalMux I__2835 (
            .O(N__18643),
            .I(\POWERLED.count_0_15 ));
    CascadeMux I__2834 (
            .O(N__18640),
            .I(N__18637));
    InMux I__2833 (
            .O(N__18637),
            .I(N__18631));
    InMux I__2832 (
            .O(N__18636),
            .I(N__18631));
    LocalMux I__2831 (
            .O(N__18631),
            .I(\POWERLED.un1_count_cry_6_c_RNIGCZ0Z59 ));
    InMux I__2830 (
            .O(N__18628),
            .I(N__18625));
    LocalMux I__2829 (
            .O(N__18625),
            .I(\POWERLED.count_0_7 ));
    CascadeMux I__2828 (
            .O(N__18622),
            .I(N__18619));
    InMux I__2827 (
            .O(N__18619),
            .I(N__18613));
    InMux I__2826 (
            .O(N__18618),
            .I(N__18613));
    LocalMux I__2825 (
            .O(N__18613),
            .I(\POWERLED.un1_count_cry_7_c_RNIHEZ0Z69 ));
    InMux I__2824 (
            .O(N__18610),
            .I(N__18607));
    LocalMux I__2823 (
            .O(N__18607),
            .I(\POWERLED.count_0_8 ));
    InMux I__2822 (
            .O(N__18604),
            .I(N__18601));
    LocalMux I__2821 (
            .O(N__18601),
            .I(N__18598));
    Span4Mux_h I__2820 (
            .O(N__18598),
            .I(N__18595));
    Odrv4 I__2819 (
            .O(N__18595),
            .I(\COUNTER.counter_1_cry_1_THRU_CO ));
    InMux I__2818 (
            .O(N__18592),
            .I(N__18587));
    CascadeMux I__2817 (
            .O(N__18591),
            .I(N__18584));
    InMux I__2816 (
            .O(N__18590),
            .I(N__18581));
    LocalMux I__2815 (
            .O(N__18587),
            .I(N__18578));
    InMux I__2814 (
            .O(N__18584),
            .I(N__18575));
    LocalMux I__2813 (
            .O(N__18581),
            .I(\COUNTER.counterZ0Z_2 ));
    Odrv12 I__2812 (
            .O(N__18578),
            .I(\COUNTER.counterZ0Z_2 ));
    LocalMux I__2811 (
            .O(N__18575),
            .I(\COUNTER.counterZ0Z_2 ));
    InMux I__2810 (
            .O(N__18568),
            .I(N__18565));
    LocalMux I__2809 (
            .O(N__18565),
            .I(\POWERLED.count_off_0_13 ));
    InMux I__2808 (
            .O(N__18562),
            .I(N__18559));
    LocalMux I__2807 (
            .O(N__18559),
            .I(\POWERLED.count_off_0_5 ));
    InMux I__2806 (
            .O(N__18556),
            .I(N__18553));
    LocalMux I__2805 (
            .O(N__18553),
            .I(\POWERLED.count_off_0_14 ));
    InMux I__2804 (
            .O(N__18550),
            .I(N__18547));
    LocalMux I__2803 (
            .O(N__18547),
            .I(\POWERLED.count_off_0_6 ));
    CascadeMux I__2802 (
            .O(N__18544),
            .I(N__18541));
    InMux I__2801 (
            .O(N__18541),
            .I(N__18538));
    LocalMux I__2800 (
            .O(N__18538),
            .I(\POWERLED.count_off_0_3 ));
    InMux I__2799 (
            .O(N__18535),
            .I(N__18532));
    LocalMux I__2798 (
            .O(N__18532),
            .I(\POWERLED.count_off_1_0 ));
    CascadeMux I__2797 (
            .O(N__18529),
            .I(\POWERLED.count_offZ0Z_0_cascade_ ));
    InMux I__2796 (
            .O(N__18526),
            .I(N__18523));
    LocalMux I__2795 (
            .O(N__18523),
            .I(\POWERLED.count_off_0_0 ));
    InMux I__2794 (
            .O(N__18520),
            .I(N__18516));
    CascadeMux I__2793 (
            .O(N__18519),
            .I(N__18513));
    LocalMux I__2792 (
            .O(N__18516),
            .I(N__18510));
    InMux I__2791 (
            .O(N__18513),
            .I(N__18507));
    Span4Mux_h I__2790 (
            .O(N__18510),
            .I(N__18502));
    LocalMux I__2789 (
            .O(N__18507),
            .I(N__18502));
    Span4Mux_s2_h I__2788 (
            .O(N__18502),
            .I(N__18497));
    InMux I__2787 (
            .O(N__18501),
            .I(N__18492));
    InMux I__2786 (
            .O(N__18500),
            .I(N__18492));
    Odrv4 I__2785 (
            .O(N__18497),
            .I(\COUNTER.counterZ0Z_0 ));
    LocalMux I__2784 (
            .O(N__18492),
            .I(\COUNTER.counterZ0Z_0 ));
    InMux I__2783 (
            .O(N__18487),
            .I(N__18484));
    LocalMux I__2782 (
            .O(N__18484),
            .I(\POWERLED.count_off_RNIZ0Z_1 ));
    InMux I__2781 (
            .O(N__18481),
            .I(N__18478));
    LocalMux I__2780 (
            .O(N__18478),
            .I(\POWERLED.count_off_0_1 ));
    CascadeMux I__2779 (
            .O(N__18475),
            .I(\POWERLED.count_off_RNIZ0Z_1_cascade_ ));
    InMux I__2778 (
            .O(N__18472),
            .I(N__18469));
    LocalMux I__2777 (
            .O(N__18469),
            .I(N__18466));
    Odrv4 I__2776 (
            .O(N__18466),
            .I(\POWERLED.un34_clk_100khz_10 ));
    CascadeMux I__2775 (
            .O(N__18463),
            .I(\POWERLED.func_state_1_m0_0_cascade_ ));
    InMux I__2774 (
            .O(N__18460),
            .I(N__18457));
    LocalMux I__2773 (
            .O(N__18457),
            .I(N__18453));
    InMux I__2772 (
            .O(N__18456),
            .I(N__18450));
    Span4Mux_v I__2771 (
            .O(N__18453),
            .I(N__18444));
    LocalMux I__2770 (
            .O(N__18450),
            .I(N__18444));
    InMux I__2769 (
            .O(N__18449),
            .I(N__18441));
    Odrv4 I__2768 (
            .O(N__18444),
            .I(\POWERLED.count_clk_RNIZ0Z_7 ));
    LocalMux I__2767 (
            .O(N__18441),
            .I(\POWERLED.count_clk_RNIZ0Z_7 ));
    CascadeMux I__2766 (
            .O(N__18436),
            .I(\POWERLED.un34_clk_100khz_11_cascade_ ));
    InMux I__2765 (
            .O(N__18433),
            .I(N__18430));
    LocalMux I__2764 (
            .O(N__18430),
            .I(\POWERLED.un34_clk_100khz_8 ));
    CascadeMux I__2763 (
            .O(N__18427),
            .I(N__18424));
    InMux I__2762 (
            .O(N__18424),
            .I(N__18421));
    LocalMux I__2761 (
            .O(N__18421),
            .I(N__18416));
    InMux I__2760 (
            .O(N__18420),
            .I(N__18413));
    InMux I__2759 (
            .O(N__18419),
            .I(N__18410));
    Span4Mux_h I__2758 (
            .O(N__18416),
            .I(N__18407));
    LocalMux I__2757 (
            .O(N__18413),
            .I(\POWERLED.N_322 ));
    LocalMux I__2756 (
            .O(N__18410),
            .I(\POWERLED.N_322 ));
    Odrv4 I__2755 (
            .O(N__18407),
            .I(\POWERLED.N_322 ));
    InMux I__2754 (
            .O(N__18400),
            .I(N__18397));
    LocalMux I__2753 (
            .O(N__18397),
            .I(\POWERLED.un34_clk_100khz_9 ));
    InMux I__2752 (
            .O(N__18394),
            .I(N__18391));
    LocalMux I__2751 (
            .O(N__18391),
            .I(N__18388));
    Odrv12 I__2750 (
            .O(N__18388),
            .I(\POWERLED.mult1_un145_sum_cry_5_s ));
    InMux I__2749 (
            .O(N__18385),
            .I(N__18382));
    LocalMux I__2748 (
            .O(N__18382),
            .I(\POWERLED.mult1_un152_sum_cry_6_s ));
    InMux I__2747 (
            .O(N__18379),
            .I(\POWERLED.mult1_un152_sum_cry_5 ));
    InMux I__2746 (
            .O(N__18376),
            .I(N__18373));
    LocalMux I__2745 (
            .O(N__18373),
            .I(N__18370));
    Odrv12 I__2744 (
            .O(N__18370),
            .I(\POWERLED.mult1_un145_sum_cry_6_s ));
    CascadeMux I__2743 (
            .O(N__18367),
            .I(N__18364));
    InMux I__2742 (
            .O(N__18364),
            .I(N__18361));
    LocalMux I__2741 (
            .O(N__18361),
            .I(\POWERLED.mult1_un159_sum_axb_7 ));
    InMux I__2740 (
            .O(N__18358),
            .I(\POWERLED.mult1_un152_sum_cry_6 ));
    InMux I__2739 (
            .O(N__18355),
            .I(N__18352));
    LocalMux I__2738 (
            .O(N__18352),
            .I(N__18349));
    Odrv12 I__2737 (
            .O(N__18349),
            .I(\POWERLED.mult1_un152_sum_axb_8 ));
    InMux I__2736 (
            .O(N__18346),
            .I(\POWERLED.mult1_un152_sum_cry_7 ));
    InMux I__2735 (
            .O(N__18343),
            .I(N__18339));
    CascadeMux I__2734 (
            .O(N__18342),
            .I(N__18335));
    LocalMux I__2733 (
            .O(N__18339),
            .I(N__18330));
    InMux I__2732 (
            .O(N__18338),
            .I(N__18327));
    InMux I__2731 (
            .O(N__18335),
            .I(N__18320));
    InMux I__2730 (
            .O(N__18334),
            .I(N__18320));
    InMux I__2729 (
            .O(N__18333),
            .I(N__18320));
    Odrv12 I__2728 (
            .O(N__18330),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__2727 (
            .O(N__18327),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__2726 (
            .O(N__18320),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    CascadeMux I__2725 (
            .O(N__18313),
            .I(N__18310));
    InMux I__2724 (
            .O(N__18310),
            .I(N__18299));
    InMux I__2723 (
            .O(N__18309),
            .I(N__18299));
    InMux I__2722 (
            .O(N__18308),
            .I(N__18299));
    InMux I__2721 (
            .O(N__18307),
            .I(N__18296));
    InMux I__2720 (
            .O(N__18306),
            .I(N__18293));
    LocalMux I__2719 (
            .O(N__18299),
            .I(N__18290));
    LocalMux I__2718 (
            .O(N__18296),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__2717 (
            .O(N__18293),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    Odrv12 I__2716 (
            .O(N__18290),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    CascadeMux I__2715 (
            .O(N__18283),
            .I(N__18279));
    CascadeMux I__2714 (
            .O(N__18282),
            .I(N__18275));
    InMux I__2713 (
            .O(N__18279),
            .I(N__18268));
    InMux I__2712 (
            .O(N__18278),
            .I(N__18268));
    InMux I__2711 (
            .O(N__18275),
            .I(N__18268));
    LocalMux I__2710 (
            .O(N__18268),
            .I(\POWERLED.mult1_un145_sum_i_0_8 ));
    CascadeMux I__2709 (
            .O(N__18265),
            .I(N__18262));
    InMux I__2708 (
            .O(N__18262),
            .I(N__18259));
    LocalMux I__2707 (
            .O(N__18259),
            .I(N__18255));
    InMux I__2706 (
            .O(N__18258),
            .I(N__18252));
    Span4Mux_v I__2705 (
            .O(N__18255),
            .I(N__18246));
    LocalMux I__2704 (
            .O(N__18252),
            .I(N__18246));
    InMux I__2703 (
            .O(N__18251),
            .I(N__18243));
    Odrv4 I__2702 (
            .O(N__18246),
            .I(\POWERLED.count_clk_RNIZ0Z_9 ));
    LocalMux I__2701 (
            .O(N__18243),
            .I(\POWERLED.count_clk_RNIZ0Z_9 ));
    CascadeMux I__2700 (
            .O(N__18238),
            .I(\POWERLED.un1_func_state25_6_0_o_N_423_N_cascade_ ));
    InMux I__2699 (
            .O(N__18235),
            .I(N__18231));
    InMux I__2698 (
            .O(N__18234),
            .I(N__18228));
    LocalMux I__2697 (
            .O(N__18231),
            .I(N__18225));
    LocalMux I__2696 (
            .O(N__18228),
            .I(\POWERLED.N_348 ));
    Odrv4 I__2695 (
            .O(N__18225),
            .I(\POWERLED.N_348 ));
    InMux I__2694 (
            .O(N__18220),
            .I(N__18217));
    LocalMux I__2693 (
            .O(N__18217),
            .I(\POWERLED.func_state_1_m0_0_0_0 ));
    CascadeMux I__2692 (
            .O(N__18214),
            .I(\POWERLED.func_state_RNI5DLR_0Z0Z_0_cascade_ ));
    InMux I__2691 (
            .O(N__18211),
            .I(\POWERLED.mult1_un159_sum_cry_4 ));
    InMux I__2690 (
            .O(N__18208),
            .I(\POWERLED.mult1_un159_sum_cry_5 ));
    InMux I__2689 (
            .O(N__18205),
            .I(\POWERLED.mult1_un159_sum_cry_6 ));
    CascadeMux I__2688 (
            .O(N__18202),
            .I(N__18198));
    CascadeMux I__2687 (
            .O(N__18201),
            .I(N__18194));
    InMux I__2686 (
            .O(N__18198),
            .I(N__18187));
    InMux I__2685 (
            .O(N__18197),
            .I(N__18187));
    InMux I__2684 (
            .O(N__18194),
            .I(N__18187));
    LocalMux I__2683 (
            .O(N__18187),
            .I(\POWERLED.mult1_un152_sum_i_0_8 ));
    InMux I__2682 (
            .O(N__18184),
            .I(N__18181));
    LocalMux I__2681 (
            .O(N__18181),
            .I(N__18178));
    Odrv4 I__2680 (
            .O(N__18178),
            .I(\POWERLED.mult1_un145_sum_i ));
    CascadeMux I__2679 (
            .O(N__18175),
            .I(N__18172));
    InMux I__2678 (
            .O(N__18172),
            .I(N__18169));
    LocalMux I__2677 (
            .O(N__18169),
            .I(\POWERLED.mult1_un152_sum_cry_3_s ));
    InMux I__2676 (
            .O(N__18166),
            .I(\POWERLED.mult1_un152_sum_cry_2 ));
    CascadeMux I__2675 (
            .O(N__18163),
            .I(N__18160));
    InMux I__2674 (
            .O(N__18160),
            .I(N__18157));
    LocalMux I__2673 (
            .O(N__18157),
            .I(N__18154));
    Odrv12 I__2672 (
            .O(N__18154),
            .I(\POWERLED.mult1_un145_sum_cry_3_s ));
    CascadeMux I__2671 (
            .O(N__18151),
            .I(N__18148));
    InMux I__2670 (
            .O(N__18148),
            .I(N__18145));
    LocalMux I__2669 (
            .O(N__18145),
            .I(\POWERLED.mult1_un152_sum_cry_4_s ));
    InMux I__2668 (
            .O(N__18142),
            .I(\POWERLED.mult1_un152_sum_cry_3 ));
    CascadeMux I__2667 (
            .O(N__18139),
            .I(N__18136));
    InMux I__2666 (
            .O(N__18136),
            .I(N__18133));
    LocalMux I__2665 (
            .O(N__18133),
            .I(N__18130));
    Span4Mux_v I__2664 (
            .O(N__18130),
            .I(N__18127));
    Odrv4 I__2663 (
            .O(N__18127),
            .I(\POWERLED.mult1_un145_sum_cry_4_s ));
    InMux I__2662 (
            .O(N__18124),
            .I(N__18121));
    LocalMux I__2661 (
            .O(N__18121),
            .I(\POWERLED.mult1_un152_sum_cry_5_s ));
    InMux I__2660 (
            .O(N__18118),
            .I(\POWERLED.mult1_un152_sum_cry_4 ));
    InMux I__2659 (
            .O(N__18115),
            .I(N__18112));
    LocalMux I__2658 (
            .O(N__18112),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    InMux I__2657 (
            .O(N__18109),
            .I(\POWERLED.mult1_un124_sum_cry_5 ));
    CascadeMux I__2656 (
            .O(N__18106),
            .I(N__18103));
    InMux I__2655 (
            .O(N__18103),
            .I(N__18100));
    LocalMux I__2654 (
            .O(N__18100),
            .I(\POWERLED.mult1_un131_sum_axb_8 ));
    InMux I__2653 (
            .O(N__18097),
            .I(\POWERLED.mult1_un124_sum_cry_6 ));
    InMux I__2652 (
            .O(N__18094),
            .I(\POWERLED.mult1_un124_sum_cry_7 ));
    InMux I__2651 (
            .O(N__18091),
            .I(N__18087));
    CascadeMux I__2650 (
            .O(N__18090),
            .I(N__18083));
    LocalMux I__2649 (
            .O(N__18087),
            .I(N__18078));
    InMux I__2648 (
            .O(N__18086),
            .I(N__18073));
    InMux I__2647 (
            .O(N__18083),
            .I(N__18073));
    InMux I__2646 (
            .O(N__18082),
            .I(N__18070));
    InMux I__2645 (
            .O(N__18081),
            .I(N__18067));
    Odrv4 I__2644 (
            .O(N__18078),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__2643 (
            .O(N__18073),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__2642 (
            .O(N__18070),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__2641 (
            .O(N__18067),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    CascadeMux I__2640 (
            .O(N__18058),
            .I(N__18055));
    InMux I__2639 (
            .O(N__18055),
            .I(N__18052));
    LocalMux I__2638 (
            .O(N__18052),
            .I(\POWERLED.mult1_un124_sum_axb_7_l_fx ));
    InMux I__2637 (
            .O(N__18049),
            .I(\POWERLED.mult1_un159_sum_cry_1 ));
    InMux I__2636 (
            .O(N__18046),
            .I(\POWERLED.mult1_un159_sum_cry_2 ));
    InMux I__2635 (
            .O(N__18043),
            .I(\POWERLED.mult1_un159_sum_cry_3 ));
    CascadeMux I__2634 (
            .O(N__18040),
            .I(N__18037));
    InMux I__2633 (
            .O(N__18037),
            .I(N__18034));
    LocalMux I__2632 (
            .O(N__18034),
            .I(\POWERLED.mult1_un138_sum_cry_4_s ));
    InMux I__2631 (
            .O(N__18031),
            .I(\POWERLED.mult1_un145_sum_cry_4 ));
    InMux I__2630 (
            .O(N__18028),
            .I(N__18025));
    LocalMux I__2629 (
            .O(N__18025),
            .I(\POWERLED.mult1_un138_sum_cry_5_s ));
    InMux I__2628 (
            .O(N__18022),
            .I(\POWERLED.mult1_un145_sum_cry_5 ));
    InMux I__2627 (
            .O(N__18019),
            .I(N__18016));
    LocalMux I__2626 (
            .O(N__18016),
            .I(\POWERLED.mult1_un138_sum_cry_6_s ));
    InMux I__2625 (
            .O(N__18013),
            .I(\POWERLED.mult1_un145_sum_cry_6 ));
    CascadeMux I__2624 (
            .O(N__18010),
            .I(N__18007));
    InMux I__2623 (
            .O(N__18007),
            .I(N__18004));
    LocalMux I__2622 (
            .O(N__18004),
            .I(\POWERLED.mult1_un145_sum_axb_8 ));
    InMux I__2621 (
            .O(N__18001),
            .I(\POWERLED.mult1_un145_sum_cry_7 ));
    CascadeMux I__2620 (
            .O(N__17998),
            .I(N__17993));
    InMux I__2619 (
            .O(N__17997),
            .I(N__17988));
    InMux I__2618 (
            .O(N__17996),
            .I(N__17985));
    InMux I__2617 (
            .O(N__17993),
            .I(N__17978));
    InMux I__2616 (
            .O(N__17992),
            .I(N__17978));
    InMux I__2615 (
            .O(N__17991),
            .I(N__17978));
    LocalMux I__2614 (
            .O(N__17988),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__2613 (
            .O(N__17985),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__2612 (
            .O(N__17978),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    CascadeMux I__2611 (
            .O(N__17971),
            .I(N__17967));
    CascadeMux I__2610 (
            .O(N__17970),
            .I(N__17963));
    InMux I__2609 (
            .O(N__17967),
            .I(N__17956));
    InMux I__2608 (
            .O(N__17966),
            .I(N__17956));
    InMux I__2607 (
            .O(N__17963),
            .I(N__17956));
    LocalMux I__2606 (
            .O(N__17956),
            .I(\POWERLED.mult1_un138_sum_i_0_8 ));
    CascadeMux I__2605 (
            .O(N__17953),
            .I(N__17950));
    InMux I__2604 (
            .O(N__17950),
            .I(N__17947));
    LocalMux I__2603 (
            .O(N__17947),
            .I(\POWERLED.mult1_un124_sum_cry_3_s ));
    InMux I__2602 (
            .O(N__17944),
            .I(\POWERLED.mult1_un124_sum_cry_2 ));
    InMux I__2601 (
            .O(N__17941),
            .I(N__17938));
    LocalMux I__2600 (
            .O(N__17938),
            .I(\POWERLED.mult1_un124_sum_cry_4_s ));
    InMux I__2599 (
            .O(N__17935),
            .I(\POWERLED.mult1_un124_sum_cry_3 ));
    CascadeMux I__2598 (
            .O(N__17932),
            .I(N__17929));
    InMux I__2597 (
            .O(N__17929),
            .I(N__17926));
    LocalMux I__2596 (
            .O(N__17926),
            .I(\POWERLED.mult1_un124_sum_cry_5_s ));
    InMux I__2595 (
            .O(N__17923),
            .I(\POWERLED.mult1_un124_sum_cry_4 ));
    InMux I__2594 (
            .O(N__17920),
            .I(N__17916));
    CascadeMux I__2593 (
            .O(N__17919),
            .I(N__17912));
    LocalMux I__2592 (
            .O(N__17916),
            .I(N__17908));
    InMux I__2591 (
            .O(N__17915),
            .I(N__17903));
    InMux I__2590 (
            .O(N__17912),
            .I(N__17903));
    InMux I__2589 (
            .O(N__17911),
            .I(N__17900));
    Odrv4 I__2588 (
            .O(N__17908),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__2587 (
            .O(N__17903),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__2586 (
            .O(N__17900),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    IoInMux I__2585 (
            .O(N__17893),
            .I(N__17890));
    LocalMux I__2584 (
            .O(N__17890),
            .I(N__17887));
    Span4Mux_s2_v I__2583 (
            .O(N__17887),
            .I(N__17884));
    Odrv4 I__2582 (
            .O(N__17884),
            .I(vccst_pwrgd));
    InMux I__2581 (
            .O(N__17881),
            .I(\POWERLED.mult1_un145_sum_cry_2 ));
    CascadeMux I__2580 (
            .O(N__17878),
            .I(N__17875));
    InMux I__2579 (
            .O(N__17875),
            .I(N__17872));
    LocalMux I__2578 (
            .O(N__17872),
            .I(\POWERLED.mult1_un138_sum_cry_3_s ));
    InMux I__2577 (
            .O(N__17869),
            .I(\POWERLED.mult1_un145_sum_cry_3 ));
    InMux I__2576 (
            .O(N__17866),
            .I(\POWERLED.un1_count_cry_7 ));
    InMux I__2575 (
            .O(N__17863),
            .I(bfn_5_3_0_));
    InMux I__2574 (
            .O(N__17860),
            .I(\POWERLED.un1_count_cry_9 ));
    InMux I__2573 (
            .O(N__17857),
            .I(\POWERLED.un1_count_cry_10 ));
    InMux I__2572 (
            .O(N__17854),
            .I(N__17848));
    InMux I__2571 (
            .O(N__17853),
            .I(N__17848));
    LocalMux I__2570 (
            .O(N__17848),
            .I(\POWERLED.un1_count_cry_11_c_RNISEHZ0Z7 ));
    InMux I__2569 (
            .O(N__17845),
            .I(\POWERLED.un1_count_cry_11 ));
    InMux I__2568 (
            .O(N__17842),
            .I(N__17838));
    InMux I__2567 (
            .O(N__17841),
            .I(N__17835));
    LocalMux I__2566 (
            .O(N__17838),
            .I(\POWERLED.un1_count_cry_12_c_RNITGIZ0Z7 ));
    LocalMux I__2565 (
            .O(N__17835),
            .I(\POWERLED.un1_count_cry_12_c_RNITGIZ0Z7 ));
    InMux I__2564 (
            .O(N__17830),
            .I(\POWERLED.un1_count_cry_12 ));
    InMux I__2563 (
            .O(N__17827),
            .I(\POWERLED.un1_count_cry_13 ));
    CascadeMux I__2562 (
            .O(N__17824),
            .I(N__17813));
    InMux I__2561 (
            .O(N__17823),
            .I(N__17803));
    InMux I__2560 (
            .O(N__17822),
            .I(N__17803));
    InMux I__2559 (
            .O(N__17821),
            .I(N__17803));
    InMux I__2558 (
            .O(N__17820),
            .I(N__17803));
    InMux I__2557 (
            .O(N__17819),
            .I(N__17796));
    InMux I__2556 (
            .O(N__17818),
            .I(N__17796));
    InMux I__2555 (
            .O(N__17817),
            .I(N__17796));
    InMux I__2554 (
            .O(N__17816),
            .I(N__17782));
    InMux I__2553 (
            .O(N__17813),
            .I(N__17782));
    InMux I__2552 (
            .O(N__17812),
            .I(N__17782));
    LocalMux I__2551 (
            .O(N__17803),
            .I(N__17777));
    LocalMux I__2550 (
            .O(N__17796),
            .I(N__17777));
    InMux I__2549 (
            .O(N__17795),
            .I(N__17770));
    InMux I__2548 (
            .O(N__17794),
            .I(N__17770));
    InMux I__2547 (
            .O(N__17793),
            .I(N__17770));
    InMux I__2546 (
            .O(N__17792),
            .I(N__17761));
    InMux I__2545 (
            .O(N__17791),
            .I(N__17761));
    InMux I__2544 (
            .O(N__17790),
            .I(N__17761));
    InMux I__2543 (
            .O(N__17789),
            .I(N__17761));
    LocalMux I__2542 (
            .O(N__17782),
            .I(\POWERLED.count_0_sqmuxa_i ));
    Odrv4 I__2541 (
            .O(N__17777),
            .I(\POWERLED.count_0_sqmuxa_i ));
    LocalMux I__2540 (
            .O(N__17770),
            .I(\POWERLED.count_0_sqmuxa_i ));
    LocalMux I__2539 (
            .O(N__17761),
            .I(\POWERLED.count_0_sqmuxa_i ));
    InMux I__2538 (
            .O(N__17752),
            .I(\POWERLED.un1_count_cry_14 ));
    InMux I__2537 (
            .O(N__17749),
            .I(N__17745));
    InMux I__2536 (
            .O(N__17748),
            .I(N__17742));
    LocalMux I__2535 (
            .O(N__17745),
            .I(\POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7 ));
    LocalMux I__2534 (
            .O(N__17742),
            .I(\POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7 ));
    InMux I__2533 (
            .O(N__17737),
            .I(N__17734));
    LocalMux I__2532 (
            .O(N__17734),
            .I(\POWERLED.count_0_14 ));
    CascadeMux I__2531 (
            .O(N__17731),
            .I(\POWERLED.count_RNIZ0Z_8_cascade_ ));
    SRMux I__2530 (
            .O(N__17728),
            .I(N__17725));
    LocalMux I__2529 (
            .O(N__17725),
            .I(\POWERLED.pwm_out_1_sqmuxa ));
    InMux I__2528 (
            .O(N__17722),
            .I(N__17716));
    InMux I__2527 (
            .O(N__17721),
            .I(N__17716));
    LocalMux I__2526 (
            .O(N__17716),
            .I(\POWERLED.N_8 ));
    InMux I__2525 (
            .O(N__17713),
            .I(\POWERLED.un1_count_cry_1 ));
    CascadeMux I__2524 (
            .O(N__17710),
            .I(N__17707));
    InMux I__2523 (
            .O(N__17707),
            .I(N__17701));
    InMux I__2522 (
            .O(N__17706),
            .I(N__17701));
    LocalMux I__2521 (
            .O(N__17701),
            .I(\POWERLED.un1_count_cry_2_c_RNICZ0Z419 ));
    InMux I__2520 (
            .O(N__17698),
            .I(\POWERLED.un1_count_cry_2 ));
    InMux I__2519 (
            .O(N__17695),
            .I(N__17692));
    LocalMux I__2518 (
            .O(N__17692),
            .I(N__17688));
    InMux I__2517 (
            .O(N__17691),
            .I(N__17685));
    Odrv4 I__2516 (
            .O(N__17688),
            .I(\POWERLED.un1_count_cry_3_c_RNIDZ0Z629 ));
    LocalMux I__2515 (
            .O(N__17685),
            .I(\POWERLED.un1_count_cry_3_c_RNIDZ0Z629 ));
    InMux I__2514 (
            .O(N__17680),
            .I(\POWERLED.un1_count_cry_3 ));
    InMux I__2513 (
            .O(N__17677),
            .I(N__17674));
    LocalMux I__2512 (
            .O(N__17674),
            .I(N__17670));
    InMux I__2511 (
            .O(N__17673),
            .I(N__17667));
    Odrv4 I__2510 (
            .O(N__17670),
            .I(\POWERLED.un1_count_cry_4_c_RNIEZ0Z839 ));
    LocalMux I__2509 (
            .O(N__17667),
            .I(\POWERLED.un1_count_cry_4_c_RNIEZ0Z839 ));
    InMux I__2508 (
            .O(N__17662),
            .I(\POWERLED.un1_count_cry_4 ));
    InMux I__2507 (
            .O(N__17659),
            .I(\POWERLED.un1_count_cry_5 ));
    InMux I__2506 (
            .O(N__17656),
            .I(\POWERLED.un1_count_cry_6 ));
    CascadeMux I__2505 (
            .O(N__17653),
            .I(N__17650));
    InMux I__2504 (
            .O(N__17650),
            .I(N__17647));
    LocalMux I__2503 (
            .O(N__17647),
            .I(N__17643));
    InMux I__2502 (
            .O(N__17646),
            .I(N__17640));
    Span4Mux_s1_v I__2501 (
            .O(N__17643),
            .I(N__17637));
    LocalMux I__2500 (
            .O(N__17640),
            .I(\DSW_PWRGD.countZ0Z_13 ));
    Odrv4 I__2499 (
            .O(N__17637),
            .I(\DSW_PWRGD.countZ0Z_13 ));
    InMux I__2498 (
            .O(N__17632),
            .I(\DSW_PWRGD.un1_count_1_cry_12 ));
    InMux I__2497 (
            .O(N__17629),
            .I(N__17625));
    InMux I__2496 (
            .O(N__17628),
            .I(N__17622));
    LocalMux I__2495 (
            .O(N__17625),
            .I(N__17619));
    LocalMux I__2494 (
            .O(N__17622),
            .I(N__17614));
    Span4Mux_s1_v I__2493 (
            .O(N__17619),
            .I(N__17614));
    Odrv4 I__2492 (
            .O(N__17614),
            .I(\DSW_PWRGD.countZ0Z_14 ));
    InMux I__2491 (
            .O(N__17611),
            .I(\DSW_PWRGD.un1_count_1_cry_13 ));
    InMux I__2490 (
            .O(N__17608),
            .I(bfn_4_16_0_));
    InMux I__2489 (
            .O(N__17605),
            .I(N__17602));
    LocalMux I__2488 (
            .O(N__17602),
            .I(N__17598));
    InMux I__2487 (
            .O(N__17601),
            .I(N__17595));
    Span4Mux_s2_h I__2486 (
            .O(N__17598),
            .I(N__17592));
    LocalMux I__2485 (
            .O(N__17595),
            .I(\DSW_PWRGD.countZ0Z_15 ));
    Odrv4 I__2484 (
            .O(N__17592),
            .I(\DSW_PWRGD.countZ0Z_15 ));
    CEMux I__2483 (
            .O(N__17587),
            .I(N__17584));
    LocalMux I__2482 (
            .O(N__17584),
            .I(N__17581));
    Span4Mux_s1_v I__2481 (
            .O(N__17581),
            .I(N__17578));
    Odrv4 I__2480 (
            .O(N__17578),
            .I(\DSW_PWRGD.N_42_1 ));
    SRMux I__2479 (
            .O(N__17575),
            .I(N__17571));
    SRMux I__2478 (
            .O(N__17574),
            .I(N__17568));
    LocalMux I__2477 (
            .O(N__17571),
            .I(N__17564));
    LocalMux I__2476 (
            .O(N__17568),
            .I(N__17561));
    SRMux I__2475 (
            .O(N__17567),
            .I(N__17558));
    Span4Mux_s1_v I__2474 (
            .O(N__17564),
            .I(N__17551));
    Span4Mux_v I__2473 (
            .O(N__17561),
            .I(N__17551));
    LocalMux I__2472 (
            .O(N__17558),
            .I(N__17551));
    Odrv4 I__2471 (
            .O(N__17551),
            .I(G_28));
    CascadeMux I__2470 (
            .O(N__17548),
            .I(\POWERLED.un79_clk_100khzlt6_cascade_ ));
    CascadeMux I__2469 (
            .O(N__17545),
            .I(\POWERLED.un79_clk_100khzlto15_5_cascade_ ));
    CascadeMux I__2468 (
            .O(N__17542),
            .I(\POWERLED.un79_clk_100khzlto15_7_cascade_ ));
    InMux I__2467 (
            .O(N__17539),
            .I(N__17536));
    LocalMux I__2466 (
            .O(N__17536),
            .I(\POWERLED.un79_clk_100khzlto15_3 ));
    InMux I__2465 (
            .O(N__17533),
            .I(N__17529));
    InMux I__2464 (
            .O(N__17532),
            .I(N__17526));
    LocalMux I__2463 (
            .O(N__17529),
            .I(N__17523));
    LocalMux I__2462 (
            .O(N__17526),
            .I(\DSW_PWRGD.countZ0Z_5 ));
    Odrv4 I__2461 (
            .O(N__17523),
            .I(\DSW_PWRGD.countZ0Z_5 ));
    InMux I__2460 (
            .O(N__17518),
            .I(\DSW_PWRGD.un1_count_1_cry_4 ));
    InMux I__2459 (
            .O(N__17515),
            .I(N__17511));
    InMux I__2458 (
            .O(N__17514),
            .I(N__17508));
    LocalMux I__2457 (
            .O(N__17511),
            .I(N__17505));
    LocalMux I__2456 (
            .O(N__17508),
            .I(\DSW_PWRGD.countZ0Z_6 ));
    Odrv4 I__2455 (
            .O(N__17505),
            .I(\DSW_PWRGD.countZ0Z_6 ));
    InMux I__2454 (
            .O(N__17500),
            .I(\DSW_PWRGD.un1_count_1_cry_5 ));
    InMux I__2453 (
            .O(N__17497),
            .I(N__17493));
    InMux I__2452 (
            .O(N__17496),
            .I(N__17490));
    LocalMux I__2451 (
            .O(N__17493),
            .I(N__17487));
    LocalMux I__2450 (
            .O(N__17490),
            .I(N__17482));
    Span4Mux_s2_h I__2449 (
            .O(N__17487),
            .I(N__17482));
    Odrv4 I__2448 (
            .O(N__17482),
            .I(\DSW_PWRGD.countZ0Z_7 ));
    InMux I__2447 (
            .O(N__17479),
            .I(\DSW_PWRGD.un1_count_1_cry_6 ));
    InMux I__2446 (
            .O(N__17476),
            .I(N__17472));
    InMux I__2445 (
            .O(N__17475),
            .I(N__17469));
    LocalMux I__2444 (
            .O(N__17472),
            .I(N__17466));
    LocalMux I__2443 (
            .O(N__17469),
            .I(\DSW_PWRGD.countZ0Z_8 ));
    Odrv4 I__2442 (
            .O(N__17466),
            .I(\DSW_PWRGD.countZ0Z_8 ));
    InMux I__2441 (
            .O(N__17461),
            .I(bfn_4_15_0_));
    InMux I__2440 (
            .O(N__17458),
            .I(N__17454));
    InMux I__2439 (
            .O(N__17457),
            .I(N__17451));
    LocalMux I__2438 (
            .O(N__17454),
            .I(N__17448));
    LocalMux I__2437 (
            .O(N__17451),
            .I(N__17443));
    Span4Mux_v I__2436 (
            .O(N__17448),
            .I(N__17443));
    Odrv4 I__2435 (
            .O(N__17443),
            .I(\DSW_PWRGD.countZ0Z_9 ));
    InMux I__2434 (
            .O(N__17440),
            .I(\DSW_PWRGD.un1_count_1_cry_8 ));
    InMux I__2433 (
            .O(N__17437),
            .I(N__17433));
    InMux I__2432 (
            .O(N__17436),
            .I(N__17430));
    LocalMux I__2431 (
            .O(N__17433),
            .I(N__17427));
    LocalMux I__2430 (
            .O(N__17430),
            .I(\DSW_PWRGD.countZ0Z_10 ));
    Odrv12 I__2429 (
            .O(N__17427),
            .I(\DSW_PWRGD.countZ0Z_10 ));
    InMux I__2428 (
            .O(N__17422),
            .I(\DSW_PWRGD.un1_count_1_cry_9 ));
    InMux I__2427 (
            .O(N__17419),
            .I(N__17415));
    InMux I__2426 (
            .O(N__17418),
            .I(N__17412));
    LocalMux I__2425 (
            .O(N__17415),
            .I(N__17409));
    LocalMux I__2424 (
            .O(N__17412),
            .I(\DSW_PWRGD.countZ0Z_11 ));
    Odrv4 I__2423 (
            .O(N__17409),
            .I(\DSW_PWRGD.countZ0Z_11 ));
    InMux I__2422 (
            .O(N__17404),
            .I(\DSW_PWRGD.un1_count_1_cry_10 ));
    InMux I__2421 (
            .O(N__17401),
            .I(N__17398));
    LocalMux I__2420 (
            .O(N__17398),
            .I(N__17394));
    InMux I__2419 (
            .O(N__17397),
            .I(N__17391));
    Span4Mux_s1_v I__2418 (
            .O(N__17394),
            .I(N__17388));
    LocalMux I__2417 (
            .O(N__17391),
            .I(\DSW_PWRGD.countZ0Z_12 ));
    Odrv4 I__2416 (
            .O(N__17388),
            .I(\DSW_PWRGD.countZ0Z_12 ));
    InMux I__2415 (
            .O(N__17383),
            .I(\DSW_PWRGD.un1_count_1_cry_11 ));
    InMux I__2414 (
            .O(N__17380),
            .I(N__17376));
    InMux I__2413 (
            .O(N__17379),
            .I(N__17372));
    LocalMux I__2412 (
            .O(N__17376),
            .I(N__17369));
    InMux I__2411 (
            .O(N__17375),
            .I(N__17366));
    LocalMux I__2410 (
            .O(N__17372),
            .I(\COUNTER.counterZ0Z_1 ));
    Odrv12 I__2409 (
            .O(N__17369),
            .I(\COUNTER.counterZ0Z_1 ));
    LocalMux I__2408 (
            .O(N__17366),
            .I(\COUNTER.counterZ0Z_1 ));
    InMux I__2407 (
            .O(N__17359),
            .I(N__17356));
    LocalMux I__2406 (
            .O(N__17356),
            .I(N__17351));
    InMux I__2405 (
            .O(N__17355),
            .I(N__17346));
    InMux I__2404 (
            .O(N__17354),
            .I(N__17346));
    Odrv12 I__2403 (
            .O(N__17351),
            .I(\COUNTER.counterZ0Z_5 ));
    LocalMux I__2402 (
            .O(N__17346),
            .I(\COUNTER.counterZ0Z_5 ));
    InMux I__2401 (
            .O(N__17341),
            .I(N__17337));
    InMux I__2400 (
            .O(N__17340),
            .I(N__17334));
    LocalMux I__2399 (
            .O(N__17337),
            .I(N__17331));
    LocalMux I__2398 (
            .O(N__17334),
            .I(\COUNTER.counterZ0Z_7 ));
    Odrv12 I__2397 (
            .O(N__17331),
            .I(\COUNTER.counterZ0Z_7 ));
    CascadeMux I__2396 (
            .O(N__17326),
            .I(N__17323));
    InMux I__2395 (
            .O(N__17323),
            .I(N__17320));
    LocalMux I__2394 (
            .O(N__17320),
            .I(\COUNTER.un4_counter_1_and ));
    InMux I__2393 (
            .O(N__17317),
            .I(N__17314));
    LocalMux I__2392 (
            .O(N__17314),
            .I(N__17311));
    Odrv4 I__2391 (
            .O(N__17311),
            .I(\COUNTER.counter_1_cry_3_THRU_CO ));
    InMux I__2390 (
            .O(N__17308),
            .I(N__17304));
    CascadeMux I__2389 (
            .O(N__17307),
            .I(N__17301));
    LocalMux I__2388 (
            .O(N__17304),
            .I(N__17297));
    InMux I__2387 (
            .O(N__17301),
            .I(N__17292));
    InMux I__2386 (
            .O(N__17300),
            .I(N__17292));
    Odrv4 I__2385 (
            .O(N__17297),
            .I(\COUNTER.counterZ0Z_4 ));
    LocalMux I__2384 (
            .O(N__17292),
            .I(\COUNTER.counterZ0Z_4 ));
    InMux I__2383 (
            .O(N__17287),
            .I(N__17284));
    LocalMux I__2382 (
            .O(N__17284),
            .I(N__17281));
    Odrv12 I__2381 (
            .O(N__17281),
            .I(\COUNTER.counter_1_cry_5_THRU_CO ));
    InMux I__2380 (
            .O(N__17278),
            .I(N__17273));
    CascadeMux I__2379 (
            .O(N__17277),
            .I(N__17270));
    InMux I__2378 (
            .O(N__17276),
            .I(N__17267));
    LocalMux I__2377 (
            .O(N__17273),
            .I(N__17264));
    InMux I__2376 (
            .O(N__17270),
            .I(N__17261));
    LocalMux I__2375 (
            .O(N__17267),
            .I(\COUNTER.counterZ0Z_6 ));
    Odrv4 I__2374 (
            .O(N__17264),
            .I(\COUNTER.counterZ0Z_6 ));
    LocalMux I__2373 (
            .O(N__17261),
            .I(\COUNTER.counterZ0Z_6 ));
    CascadeMux I__2372 (
            .O(N__17254),
            .I(N__17250));
    InMux I__2371 (
            .O(N__17253),
            .I(N__17247));
    InMux I__2370 (
            .O(N__17250),
            .I(N__17244));
    LocalMux I__2369 (
            .O(N__17247),
            .I(N__17239));
    LocalMux I__2368 (
            .O(N__17244),
            .I(N__17239));
    Span4Mux_h I__2367 (
            .O(N__17239),
            .I(N__17236));
    Odrv4 I__2366 (
            .O(N__17236),
            .I(\DSW_PWRGD.un1_curr_state10_0 ));
    CascadeMux I__2365 (
            .O(N__17233),
            .I(N__17230));
    InMux I__2364 (
            .O(N__17230),
            .I(N__17227));
    LocalMux I__2363 (
            .O(N__17227),
            .I(N__17223));
    InMux I__2362 (
            .O(N__17226),
            .I(N__17220));
    Span4Mux_s3_h I__2361 (
            .O(N__17223),
            .I(N__17217));
    LocalMux I__2360 (
            .O(N__17220),
            .I(\DSW_PWRGD.countZ0Z_0 ));
    Odrv4 I__2359 (
            .O(N__17217),
            .I(\DSW_PWRGD.countZ0Z_0 ));
    InMux I__2358 (
            .O(N__17212),
            .I(N__17209));
    LocalMux I__2357 (
            .O(N__17209),
            .I(N__17205));
    InMux I__2356 (
            .O(N__17208),
            .I(N__17202));
    Span4Mux_s2_h I__2355 (
            .O(N__17205),
            .I(N__17199));
    LocalMux I__2354 (
            .O(N__17202),
            .I(\DSW_PWRGD.countZ0Z_1 ));
    Odrv4 I__2353 (
            .O(N__17199),
            .I(\DSW_PWRGD.countZ0Z_1 ));
    InMux I__2352 (
            .O(N__17194),
            .I(\DSW_PWRGD.un1_count_1_cry_0 ));
    InMux I__2351 (
            .O(N__17191),
            .I(N__17187));
    InMux I__2350 (
            .O(N__17190),
            .I(N__17184));
    LocalMux I__2349 (
            .O(N__17187),
            .I(N__17181));
    LocalMux I__2348 (
            .O(N__17184),
            .I(\DSW_PWRGD.countZ0Z_2 ));
    Odrv12 I__2347 (
            .O(N__17181),
            .I(\DSW_PWRGD.countZ0Z_2 ));
    InMux I__2346 (
            .O(N__17176),
            .I(\DSW_PWRGD.un1_count_1_cry_1 ));
    CascadeMux I__2345 (
            .O(N__17173),
            .I(N__17170));
    InMux I__2344 (
            .O(N__17170),
            .I(N__17167));
    LocalMux I__2343 (
            .O(N__17167),
            .I(N__17163));
    InMux I__2342 (
            .O(N__17166),
            .I(N__17160));
    Span4Mux_s2_h I__2341 (
            .O(N__17163),
            .I(N__17157));
    LocalMux I__2340 (
            .O(N__17160),
            .I(\DSW_PWRGD.countZ0Z_3 ));
    Odrv4 I__2339 (
            .O(N__17157),
            .I(\DSW_PWRGD.countZ0Z_3 ));
    InMux I__2338 (
            .O(N__17152),
            .I(\DSW_PWRGD.un1_count_1_cry_2 ));
    CascadeMux I__2337 (
            .O(N__17149),
            .I(N__17146));
    InMux I__2336 (
            .O(N__17146),
            .I(N__17143));
    LocalMux I__2335 (
            .O(N__17143),
            .I(N__17139));
    InMux I__2334 (
            .O(N__17142),
            .I(N__17136));
    Span4Mux_s3_h I__2333 (
            .O(N__17139),
            .I(N__17133));
    LocalMux I__2332 (
            .O(N__17136),
            .I(\DSW_PWRGD.countZ0Z_4 ));
    Odrv4 I__2331 (
            .O(N__17133),
            .I(\DSW_PWRGD.countZ0Z_4 ));
    InMux I__2330 (
            .O(N__17128),
            .I(\DSW_PWRGD.un1_count_1_cry_3 ));
    CascadeMux I__2329 (
            .O(N__17125),
            .I(N__17122));
    InMux I__2328 (
            .O(N__17122),
            .I(N__17119));
    LocalMux I__2327 (
            .O(N__17119),
            .I(N__17116));
    Span4Mux_v I__2326 (
            .O(N__17116),
            .I(N__17113));
    Odrv4 I__2325 (
            .O(N__17113),
            .I(\COUNTER.un4_counter_4_and ));
    CascadeMux I__2324 (
            .O(N__17110),
            .I(N__17107));
    InMux I__2323 (
            .O(N__17107),
            .I(N__17104));
    LocalMux I__2322 (
            .O(N__17104),
            .I(N__17101));
    Span4Mux_h I__2321 (
            .O(N__17101),
            .I(N__17098));
    Odrv4 I__2320 (
            .O(N__17098),
            .I(\COUNTER.un4_counter_5_and ));
    CascadeMux I__2319 (
            .O(N__17095),
            .I(N__17092));
    InMux I__2318 (
            .O(N__17092),
            .I(N__17089));
    LocalMux I__2317 (
            .O(N__17089),
            .I(N__17086));
    Span4Mux_h I__2316 (
            .O(N__17086),
            .I(N__17083));
    Odrv4 I__2315 (
            .O(N__17083),
            .I(\COUNTER.un4_counter_6_and ));
    CascadeMux I__2314 (
            .O(N__17080),
            .I(N__17077));
    InMux I__2313 (
            .O(N__17077),
            .I(N__17074));
    LocalMux I__2312 (
            .O(N__17074),
            .I(N__17071));
    Span4Mux_h I__2311 (
            .O(N__17071),
            .I(N__17068));
    Odrv4 I__2310 (
            .O(N__17068),
            .I(\COUNTER.un4_counter_7_and ));
    InMux I__2309 (
            .O(N__17065),
            .I(bfn_4_13_0_));
    InMux I__2308 (
            .O(N__17062),
            .I(N__17059));
    LocalMux I__2307 (
            .O(N__17059),
            .I(N__17056));
    Odrv12 I__2306 (
            .O(N__17056),
            .I(\COUNTER.counter_1_cry_4_THRU_CO ));
    InMux I__2305 (
            .O(N__17053),
            .I(N__17050));
    LocalMux I__2304 (
            .O(N__17050),
            .I(N__17047));
    Span4Mux_h I__2303 (
            .O(N__17047),
            .I(N__17044));
    Odrv4 I__2302 (
            .O(N__17044),
            .I(\COUNTER.counter_1_cry_2_THRU_CO ));
    InMux I__2301 (
            .O(N__17041),
            .I(N__17037));
    CascadeMux I__2300 (
            .O(N__17040),
            .I(N__17034));
    LocalMux I__2299 (
            .O(N__17037),
            .I(N__17030));
    InMux I__2298 (
            .O(N__17034),
            .I(N__17025));
    InMux I__2297 (
            .O(N__17033),
            .I(N__17025));
    Odrv4 I__2296 (
            .O(N__17030),
            .I(\COUNTER.counterZ0Z_3 ));
    LocalMux I__2295 (
            .O(N__17025),
            .I(\COUNTER.counterZ0Z_3 ));
    CascadeMux I__2294 (
            .O(N__17020),
            .I(N__17017));
    InMux I__2293 (
            .O(N__17017),
            .I(N__17014));
    LocalMux I__2292 (
            .O(N__17014),
            .I(\COUNTER.un4_counter_0_and ));
    CascadeMux I__2291 (
            .O(N__17011),
            .I(\POWERLED.N_321_cascade_ ));
    InMux I__2290 (
            .O(N__17008),
            .I(N__17005));
    LocalMux I__2289 (
            .O(N__17005),
            .I(\POWERLED.func_state_1_ss0_i_0_o3_0 ));
    IoInMux I__2288 (
            .O(N__17002),
            .I(N__16999));
    LocalMux I__2287 (
            .O(N__16999),
            .I(N__16996));
    Odrv12 I__2286 (
            .O(N__16996),
            .I(vccst_en));
    InMux I__2285 (
            .O(N__16993),
            .I(N__16989));
    InMux I__2284 (
            .O(N__16992),
            .I(N__16986));
    LocalMux I__2283 (
            .O(N__16989),
            .I(N__16983));
    LocalMux I__2282 (
            .O(N__16986),
            .I(\POWERLED.N_516 ));
    Odrv4 I__2281 (
            .O(N__16983),
            .I(\POWERLED.N_516 ));
    CascadeMux I__2280 (
            .O(N__16978),
            .I(\POWERLED.N_516_cascade_ ));
    InMux I__2279 (
            .O(N__16975),
            .I(N__16972));
    LocalMux I__2278 (
            .O(N__16972),
            .I(\POWERLED.N_403 ));
    CascadeMux I__2277 (
            .O(N__16969),
            .I(N__16966));
    InMux I__2276 (
            .O(N__16966),
            .I(N__16963));
    LocalMux I__2275 (
            .O(N__16963),
            .I(N__16960));
    Span4Mux_h I__2274 (
            .O(N__16960),
            .I(N__16957));
    Odrv4 I__2273 (
            .O(N__16957),
            .I(\COUNTER.un4_counter_2_and ));
    CascadeMux I__2272 (
            .O(N__16954),
            .I(N__16951));
    InMux I__2271 (
            .O(N__16951),
            .I(N__16948));
    LocalMux I__2270 (
            .O(N__16948),
            .I(N__16945));
    Span4Mux_h I__2269 (
            .O(N__16945),
            .I(N__16942));
    Odrv4 I__2268 (
            .O(N__16942),
            .I(\COUNTER.un4_counter_3_and ));
    CascadeMux I__2267 (
            .O(N__16939),
            .I(\POWERLED.count_clk_en_0_cascade_ ));
    CEMux I__2266 (
            .O(N__16936),
            .I(N__16913));
    CEMux I__2265 (
            .O(N__16935),
            .I(N__16910));
    CEMux I__2264 (
            .O(N__16934),
            .I(N__16907));
    CEMux I__2263 (
            .O(N__16933),
            .I(N__16904));
    InMux I__2262 (
            .O(N__16932),
            .I(N__16897));
    InMux I__2261 (
            .O(N__16931),
            .I(N__16897));
    InMux I__2260 (
            .O(N__16930),
            .I(N__16897));
    CEMux I__2259 (
            .O(N__16929),
            .I(N__16893));
    InMux I__2258 (
            .O(N__16928),
            .I(N__16886));
    InMux I__2257 (
            .O(N__16927),
            .I(N__16886));
    InMux I__2256 (
            .O(N__16926),
            .I(N__16886));
    CEMux I__2255 (
            .O(N__16925),
            .I(N__16883));
    InMux I__2254 (
            .O(N__16924),
            .I(N__16876));
    InMux I__2253 (
            .O(N__16923),
            .I(N__16876));
    InMux I__2252 (
            .O(N__16922),
            .I(N__16876));
    InMux I__2251 (
            .O(N__16921),
            .I(N__16873));
    InMux I__2250 (
            .O(N__16920),
            .I(N__16870));
    InMux I__2249 (
            .O(N__16919),
            .I(N__16861));
    InMux I__2248 (
            .O(N__16918),
            .I(N__16861));
    InMux I__2247 (
            .O(N__16917),
            .I(N__16861));
    InMux I__2246 (
            .O(N__16916),
            .I(N__16861));
    LocalMux I__2245 (
            .O(N__16913),
            .I(N__16856));
    LocalMux I__2244 (
            .O(N__16910),
            .I(N__16856));
    LocalMux I__2243 (
            .O(N__16907),
            .I(N__16853));
    LocalMux I__2242 (
            .O(N__16904),
            .I(N__16850));
    LocalMux I__2241 (
            .O(N__16897),
            .I(N__16847));
    InMux I__2240 (
            .O(N__16896),
            .I(N__16844));
    LocalMux I__2239 (
            .O(N__16893),
            .I(N__16841));
    LocalMux I__2238 (
            .O(N__16886),
            .I(N__16838));
    LocalMux I__2237 (
            .O(N__16883),
            .I(N__16831));
    LocalMux I__2236 (
            .O(N__16876),
            .I(N__16831));
    LocalMux I__2235 (
            .O(N__16873),
            .I(N__16831));
    LocalMux I__2234 (
            .O(N__16870),
            .I(N__16826));
    LocalMux I__2233 (
            .O(N__16861),
            .I(N__16826));
    Span4Mux_v I__2232 (
            .O(N__16856),
            .I(N__16815));
    Span4Mux_s1_h I__2231 (
            .O(N__16853),
            .I(N__16815));
    Span4Mux_v I__2230 (
            .O(N__16850),
            .I(N__16815));
    Span4Mux_s1_h I__2229 (
            .O(N__16847),
            .I(N__16815));
    LocalMux I__2228 (
            .O(N__16844),
            .I(N__16815));
    Span4Mux_s3_h I__2227 (
            .O(N__16841),
            .I(N__16810));
    Span4Mux_s3_h I__2226 (
            .O(N__16838),
            .I(N__16810));
    Span4Mux_s3_h I__2225 (
            .O(N__16831),
            .I(N__16807));
    Span4Mux_s3_h I__2224 (
            .O(N__16826),
            .I(N__16804));
    Odrv4 I__2223 (
            .O(N__16815),
            .I(\POWERLED.func_state_RNI81TV4Z0Z_1 ));
    Odrv4 I__2222 (
            .O(N__16810),
            .I(\POWERLED.func_state_RNI81TV4Z0Z_1 ));
    Odrv4 I__2221 (
            .O(N__16807),
            .I(\POWERLED.func_state_RNI81TV4Z0Z_1 ));
    Odrv4 I__2220 (
            .O(N__16804),
            .I(\POWERLED.func_state_RNI81TV4Z0Z_1 ));
    InMux I__2219 (
            .O(N__16795),
            .I(N__16792));
    LocalMux I__2218 (
            .O(N__16792),
            .I(\POWERLED.N_480 ));
    CascadeMux I__2217 (
            .O(N__16789),
            .I(\POWERLED.func_state_1_ss0_i_0_o3_1_cascade_ ));
    InMux I__2216 (
            .O(N__16786),
            .I(N__16783));
    LocalMux I__2215 (
            .O(N__16783),
            .I(N__16780));
    Odrv4 I__2214 (
            .O(N__16780),
            .I(\POWERLED.N_217 ));
    CascadeMux I__2213 (
            .O(N__16777),
            .I(\POWERLED.N_217_cascade_ ));
    CascadeMux I__2212 (
            .O(N__16774),
            .I(N__16771));
    InMux I__2211 (
            .O(N__16771),
            .I(N__16768));
    LocalMux I__2210 (
            .O(N__16768),
            .I(\POWERLED.mult1_un138_sum_axb_8 ));
    InMux I__2209 (
            .O(N__16765),
            .I(\POWERLED.mult1_un131_sum_cry_6 ));
    InMux I__2208 (
            .O(N__16762),
            .I(\POWERLED.mult1_un131_sum_cry_7 ));
    CascadeMux I__2207 (
            .O(N__16759),
            .I(\POWERLED.mult1_un131_sum_s_8_cascade_ ));
    CascadeMux I__2206 (
            .O(N__16756),
            .I(N__16752));
    CascadeMux I__2205 (
            .O(N__16755),
            .I(N__16748));
    InMux I__2204 (
            .O(N__16752),
            .I(N__16741));
    InMux I__2203 (
            .O(N__16751),
            .I(N__16741));
    InMux I__2202 (
            .O(N__16748),
            .I(N__16741));
    LocalMux I__2201 (
            .O(N__16741),
            .I(\POWERLED.mult1_un131_sum_i_0_8 ));
    CascadeMux I__2200 (
            .O(N__16738),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_0_a3_0_0_cascade_ ));
    CascadeMux I__2199 (
            .O(N__16735),
            .I(\POWERLED.N_96_cascade_ ));
    CascadeMux I__2198 (
            .O(N__16732),
            .I(N__16729));
    InMux I__2197 (
            .O(N__16729),
            .I(N__16726));
    LocalMux I__2196 (
            .O(N__16726),
            .I(N__16723));
    Odrv4 I__2195 (
            .O(N__16723),
            .I(\POWERLED.count_off_0_4 ));
    InMux I__2194 (
            .O(N__16720),
            .I(N__16717));
    LocalMux I__2193 (
            .O(N__16717),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_0_a3_1 ));
    CascadeMux I__2192 (
            .O(N__16714),
            .I(\POWERLED.N_455_cascade_ ));
    InMux I__2191 (
            .O(N__16711),
            .I(\POWERLED.mult1_un138_sum_cry_6 ));
    InMux I__2190 (
            .O(N__16708),
            .I(\POWERLED.mult1_un138_sum_cry_7 ));
    CascadeMux I__2189 (
            .O(N__16705),
            .I(N__16702));
    InMux I__2188 (
            .O(N__16702),
            .I(N__16699));
    LocalMux I__2187 (
            .O(N__16699),
            .I(\POWERLED.mult1_un131_sum_cry_3_s ));
    InMux I__2186 (
            .O(N__16696),
            .I(\POWERLED.mult1_un131_sum_cry_2 ));
    InMux I__2185 (
            .O(N__16693),
            .I(N__16690));
    LocalMux I__2184 (
            .O(N__16690),
            .I(\POWERLED.mult1_un131_sum_cry_4_s ));
    InMux I__2183 (
            .O(N__16687),
            .I(\POWERLED.mult1_un131_sum_cry_3 ));
    CascadeMux I__2182 (
            .O(N__16684),
            .I(N__16681));
    InMux I__2181 (
            .O(N__16681),
            .I(N__16678));
    LocalMux I__2180 (
            .O(N__16678),
            .I(\POWERLED.mult1_un131_sum_cry_5_s ));
    InMux I__2179 (
            .O(N__16675),
            .I(\POWERLED.mult1_un131_sum_cry_4 ));
    InMux I__2178 (
            .O(N__16672),
            .I(N__16669));
    LocalMux I__2177 (
            .O(N__16669),
            .I(\POWERLED.mult1_un131_sum_cry_6_s ));
    InMux I__2176 (
            .O(N__16666),
            .I(\POWERLED.mult1_un131_sum_cry_5 ));
    CascadeMux I__2175 (
            .O(N__16663),
            .I(N__16659));
    CascadeMux I__2174 (
            .O(N__16662),
            .I(N__16655));
    InMux I__2173 (
            .O(N__16659),
            .I(N__16648));
    InMux I__2172 (
            .O(N__16658),
            .I(N__16648));
    InMux I__2171 (
            .O(N__16655),
            .I(N__16648));
    LocalMux I__2170 (
            .O(N__16648),
            .I(\POWERLED.mult1_un124_sum_i_0_8 ));
    InMux I__2169 (
            .O(N__16645),
            .I(N__16642));
    LocalMux I__2168 (
            .O(N__16642),
            .I(N__16639));
    Odrv4 I__2167 (
            .O(N__16639),
            .I(\POWERLED.count_0_13 ));
    InMux I__2166 (
            .O(N__16636),
            .I(N__16633));
    LocalMux I__2165 (
            .O(N__16633),
            .I(N__16630));
    Odrv4 I__2164 (
            .O(N__16630),
            .I(\POWERLED.count_0_4 ));
    InMux I__2163 (
            .O(N__16627),
            .I(N__16624));
    LocalMux I__2162 (
            .O(N__16624),
            .I(\POWERLED.count_0_5 ));
    InMux I__2161 (
            .O(N__16621),
            .I(\POWERLED.mult1_un138_sum_cry_2 ));
    InMux I__2160 (
            .O(N__16618),
            .I(\POWERLED.mult1_un138_sum_cry_3 ));
    InMux I__2159 (
            .O(N__16615),
            .I(\POWERLED.mult1_un138_sum_cry_4 ));
    InMux I__2158 (
            .O(N__16612),
            .I(\POWERLED.mult1_un138_sum_cry_5 ));
    InMux I__2157 (
            .O(N__16609),
            .I(N__16606));
    LocalMux I__2156 (
            .O(N__16606),
            .I(\POWERLED.count_0_3 ));
    InMux I__2155 (
            .O(N__16603),
            .I(N__16600));
    LocalMux I__2154 (
            .O(N__16600),
            .I(\POWERLED.count_0_12 ));
    InMux I__2153 (
            .O(N__16597),
            .I(N__16594));
    LocalMux I__2152 (
            .O(N__16594),
            .I(N__16590));
    InMux I__2151 (
            .O(N__16593),
            .I(N__16587));
    Span4Mux_s2_v I__2150 (
            .O(N__16590),
            .I(N__16584));
    LocalMux I__2149 (
            .O(N__16587),
            .I(N__16581));
    Odrv4 I__2148 (
            .O(N__16584),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    Odrv12 I__2147 (
            .O(N__16581),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    CascadeMux I__2146 (
            .O(N__16576),
            .I(N__16573));
    InMux I__2145 (
            .O(N__16573),
            .I(N__16567));
    InMux I__2144 (
            .O(N__16572),
            .I(N__16567));
    LocalMux I__2143 (
            .O(N__16567),
            .I(N__16564));
    Odrv12 I__2142 (
            .O(N__16564),
            .I(\PCH_PWRGD.count_rst ));
    InMux I__2141 (
            .O(N__16561),
            .I(N__16558));
    LocalMux I__2140 (
            .O(N__16558),
            .I(\PCH_PWRGD.count_0_15 ));
    InMux I__2139 (
            .O(N__16555),
            .I(N__16552));
    LocalMux I__2138 (
            .O(N__16552),
            .I(N__16549));
    Span4Mux_v I__2137 (
            .O(N__16549),
            .I(N__16545));
    InMux I__2136 (
            .O(N__16548),
            .I(N__16542));
    Odrv4 I__2135 (
            .O(N__16545),
            .I(\PCH_PWRGD.N_2110_i ));
    LocalMux I__2134 (
            .O(N__16542),
            .I(\PCH_PWRGD.N_2110_i ));
    InMux I__2133 (
            .O(N__16537),
            .I(N__16532));
    InMux I__2132 (
            .O(N__16536),
            .I(N__16529));
    InMux I__2131 (
            .O(N__16535),
            .I(N__16526));
    LocalMux I__2130 (
            .O(N__16532),
            .I(N__16523));
    LocalMux I__2129 (
            .O(N__16529),
            .I(N__16516));
    LocalMux I__2128 (
            .O(N__16526),
            .I(N__16516));
    Span4Mux_h I__2127 (
            .O(N__16523),
            .I(N__16516));
    Span4Mux_v I__2126 (
            .O(N__16516),
            .I(N__16513));
    Odrv4 I__2125 (
            .O(N__16513),
            .I(\PCH_PWRGD.N_314 ));
    InMux I__2124 (
            .O(N__16510),
            .I(N__16503));
    InMux I__2123 (
            .O(N__16509),
            .I(N__16503));
    CascadeMux I__2122 (
            .O(N__16508),
            .I(N__16500));
    LocalMux I__2121 (
            .O(N__16503),
            .I(N__16497));
    InMux I__2120 (
            .O(N__16500),
            .I(N__16494));
    Span4Mux_v I__2119 (
            .O(N__16497),
            .I(N__16491));
    LocalMux I__2118 (
            .O(N__16494),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    Odrv4 I__2117 (
            .O(N__16491),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    InMux I__2116 (
            .O(N__16486),
            .I(N__16480));
    InMux I__2115 (
            .O(N__16485),
            .I(N__16473));
    InMux I__2114 (
            .O(N__16484),
            .I(N__16473));
    InMux I__2113 (
            .O(N__16483),
            .I(N__16473));
    LocalMux I__2112 (
            .O(N__16480),
            .I(N__16468));
    LocalMux I__2111 (
            .O(N__16473),
            .I(N__16468));
    Span4Mux_v I__2110 (
            .O(N__16468),
            .I(N__16465));
    Odrv4 I__2109 (
            .O(N__16465),
            .I(\PCH_PWRGD.N_2091_i ));
    CascadeMux I__2108 (
            .O(N__16462),
            .I(\POWERLED.curr_state_3_0_cascade_ ));
    CascadeMux I__2107 (
            .O(N__16459),
            .I(\POWERLED.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__2106 (
            .O(N__16456),
            .I(\POWERLED.count_0_sqmuxa_i_cascade_ ));
    CascadeMux I__2105 (
            .O(N__16453),
            .I(\POWERLED.count_RNIZ0Z_0_cascade_ ));
    CascadeMux I__2104 (
            .O(N__16450),
            .I(\POWERLED.count_RNIZ0Z_1_cascade_ ));
    CascadeMux I__2103 (
            .O(N__16447),
            .I(\POWERLED.countZ0Z_1_cascade_ ));
    InMux I__2102 (
            .O(N__16444),
            .I(N__16441));
    LocalMux I__2101 (
            .O(N__16441),
            .I(\POWERLED.count_0_1 ));
    InMux I__2100 (
            .O(N__16438),
            .I(N__16435));
    LocalMux I__2099 (
            .O(N__16435),
            .I(\POWERLED.count_0_0 ));
    InMux I__2098 (
            .O(N__16432),
            .I(N__16429));
    LocalMux I__2097 (
            .O(N__16429),
            .I(\DSW_PWRGD.un4_count_11 ));
    InMux I__2096 (
            .O(N__16426),
            .I(N__16423));
    LocalMux I__2095 (
            .O(N__16423),
            .I(N__16420));
    Odrv12 I__2094 (
            .O(N__16420),
            .I(\DSW_PWRGD.un4_count_10 ));
    CascadeMux I__2093 (
            .O(N__16417),
            .I(\DSW_PWRGD.un4_count_9_cascade_ ));
    InMux I__2092 (
            .O(N__16414),
            .I(N__16411));
    LocalMux I__2091 (
            .O(N__16411),
            .I(N__16408));
    Odrv4 I__2090 (
            .O(N__16408),
            .I(\DSW_PWRGD.un4_count_8 ));
    CascadeMux I__2089 (
            .O(N__16405),
            .I(N__16401));
    CascadeMux I__2088 (
            .O(N__16404),
            .I(N__16398));
    InMux I__2087 (
            .O(N__16401),
            .I(N__16394));
    InMux I__2086 (
            .O(N__16398),
            .I(N__16389));
    InMux I__2085 (
            .O(N__16397),
            .I(N__16389));
    LocalMux I__2084 (
            .O(N__16394),
            .I(\DSW_PWRGD.N_1_i ));
    LocalMux I__2083 (
            .O(N__16389),
            .I(\DSW_PWRGD.N_1_i ));
    InMux I__2082 (
            .O(N__16384),
            .I(N__16380));
    InMux I__2081 (
            .O(N__16383),
            .I(N__16377));
    LocalMux I__2080 (
            .O(N__16380),
            .I(\COUNTER.counterZ0Z_22 ));
    LocalMux I__2079 (
            .O(N__16377),
            .I(\COUNTER.counterZ0Z_22 ));
    InMux I__2078 (
            .O(N__16372),
            .I(N__16368));
    InMux I__2077 (
            .O(N__16371),
            .I(N__16365));
    LocalMux I__2076 (
            .O(N__16368),
            .I(\COUNTER.counterZ0Z_20 ));
    LocalMux I__2075 (
            .O(N__16365),
            .I(\COUNTER.counterZ0Z_20 ));
    CascadeMux I__2074 (
            .O(N__16360),
            .I(N__16356));
    InMux I__2073 (
            .O(N__16359),
            .I(N__16353));
    InMux I__2072 (
            .O(N__16356),
            .I(N__16350));
    LocalMux I__2071 (
            .O(N__16353),
            .I(\COUNTER.counterZ0Z_23 ));
    LocalMux I__2070 (
            .O(N__16350),
            .I(\COUNTER.counterZ0Z_23 ));
    InMux I__2069 (
            .O(N__16345),
            .I(N__16341));
    InMux I__2068 (
            .O(N__16344),
            .I(N__16338));
    LocalMux I__2067 (
            .O(N__16341),
            .I(\COUNTER.counterZ0Z_21 ));
    LocalMux I__2066 (
            .O(N__16338),
            .I(\COUNTER.counterZ0Z_21 ));
    InMux I__2065 (
            .O(N__16333),
            .I(N__16329));
    InMux I__2064 (
            .O(N__16332),
            .I(N__16326));
    LocalMux I__2063 (
            .O(N__16329),
            .I(\COUNTER.counterZ0Z_28 ));
    LocalMux I__2062 (
            .O(N__16326),
            .I(\COUNTER.counterZ0Z_28 ));
    InMux I__2061 (
            .O(N__16321),
            .I(N__16317));
    InMux I__2060 (
            .O(N__16320),
            .I(N__16314));
    LocalMux I__2059 (
            .O(N__16317),
            .I(\COUNTER.counterZ0Z_30 ));
    LocalMux I__2058 (
            .O(N__16314),
            .I(\COUNTER.counterZ0Z_30 ));
    CascadeMux I__2057 (
            .O(N__16309),
            .I(N__16305));
    InMux I__2056 (
            .O(N__16308),
            .I(N__16302));
    InMux I__2055 (
            .O(N__16305),
            .I(N__16299));
    LocalMux I__2054 (
            .O(N__16302),
            .I(\COUNTER.counterZ0Z_29 ));
    LocalMux I__2053 (
            .O(N__16299),
            .I(\COUNTER.counterZ0Z_29 ));
    InMux I__2052 (
            .O(N__16294),
            .I(N__16290));
    InMux I__2051 (
            .O(N__16293),
            .I(N__16287));
    LocalMux I__2050 (
            .O(N__16290),
            .I(\COUNTER.counterZ0Z_31 ));
    LocalMux I__2049 (
            .O(N__16287),
            .I(\COUNTER.counterZ0Z_31 ));
    InMux I__2048 (
            .O(N__16282),
            .I(N__16278));
    InMux I__2047 (
            .O(N__16281),
            .I(N__16275));
    LocalMux I__2046 (
            .O(N__16278),
            .I(\COUNTER.counterZ0Z_25 ));
    LocalMux I__2045 (
            .O(N__16275),
            .I(\COUNTER.counterZ0Z_25 ));
    InMux I__2044 (
            .O(N__16270),
            .I(N__16266));
    InMux I__2043 (
            .O(N__16269),
            .I(N__16263));
    LocalMux I__2042 (
            .O(N__16266),
            .I(\COUNTER.counterZ0Z_24 ));
    LocalMux I__2041 (
            .O(N__16263),
            .I(\COUNTER.counterZ0Z_24 ));
    CascadeMux I__2040 (
            .O(N__16258),
            .I(N__16254));
    InMux I__2039 (
            .O(N__16257),
            .I(N__16251));
    InMux I__2038 (
            .O(N__16254),
            .I(N__16248));
    LocalMux I__2037 (
            .O(N__16251),
            .I(\COUNTER.counterZ0Z_26 ));
    LocalMux I__2036 (
            .O(N__16248),
            .I(\COUNTER.counterZ0Z_26 ));
    InMux I__2035 (
            .O(N__16243),
            .I(N__16239));
    InMux I__2034 (
            .O(N__16242),
            .I(N__16236));
    LocalMux I__2033 (
            .O(N__16239),
            .I(\COUNTER.counterZ0Z_27 ));
    LocalMux I__2032 (
            .O(N__16236),
            .I(\COUNTER.counterZ0Z_27 ));
    CascadeMux I__2031 (
            .O(N__16231),
            .I(\POWERLED.g0_i_o3_0_cascade_ ));
    InMux I__2030 (
            .O(N__16228),
            .I(N__16222));
    InMux I__2029 (
            .O(N__16227),
            .I(N__16222));
    LocalMux I__2028 (
            .O(N__16222),
            .I(\POWERLED.pwm_outZ0 ));
    InMux I__2027 (
            .O(N__16219),
            .I(N__16216));
    LocalMux I__2026 (
            .O(N__16216),
            .I(\POWERLED.g0_i_o3_0 ));
    IoInMux I__2025 (
            .O(N__16213),
            .I(N__16210));
    LocalMux I__2024 (
            .O(N__16210),
            .I(N__16207));
    IoSpan4Mux I__2023 (
            .O(N__16207),
            .I(N__16204));
    Span4Mux_s3_h I__2022 (
            .O(N__16204),
            .I(N__16201));
    Sp12to4 I__2021 (
            .O(N__16201),
            .I(N__16198));
    Span12Mux_v I__2020 (
            .O(N__16198),
            .I(N__16195));
    Odrv12 I__2019 (
            .O(N__16195),
            .I(pwrbtn_led));
    InMux I__2018 (
            .O(N__16192),
            .I(N__16181));
    InMux I__2017 (
            .O(N__16191),
            .I(N__16181));
    InMux I__2016 (
            .O(N__16190),
            .I(N__16181));
    InMux I__2015 (
            .O(N__16189),
            .I(N__16176));
    InMux I__2014 (
            .O(N__16188),
            .I(N__16176));
    LocalMux I__2013 (
            .O(N__16181),
            .I(N__16171));
    LocalMux I__2012 (
            .O(N__16176),
            .I(N__16171));
    Span4Mux_s3_v I__2011 (
            .O(N__16171),
            .I(N__16168));
    Odrv4 I__2010 (
            .O(N__16168),
            .I(v33dsw_ok));
    InMux I__2009 (
            .O(N__16165),
            .I(N__16150));
    InMux I__2008 (
            .O(N__16164),
            .I(N__16150));
    InMux I__2007 (
            .O(N__16163),
            .I(N__16150));
    InMux I__2006 (
            .O(N__16162),
            .I(N__16150));
    InMux I__2005 (
            .O(N__16161),
            .I(N__16150));
    LocalMux I__2004 (
            .O(N__16150),
            .I(\DSW_PWRGD.curr_stateZ0Z_0 ));
    CascadeMux I__2003 (
            .O(N__16147),
            .I(N__16141));
    InMux I__2002 (
            .O(N__16146),
            .I(N__16129));
    InMux I__2001 (
            .O(N__16145),
            .I(N__16129));
    InMux I__2000 (
            .O(N__16144),
            .I(N__16129));
    InMux I__1999 (
            .O(N__16141),
            .I(N__16129));
    InMux I__1998 (
            .O(N__16140),
            .I(N__16129));
    LocalMux I__1997 (
            .O(N__16129),
            .I(\DSW_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__1996 (
            .O(N__16126),
            .I(DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_));
    CascadeMux I__1995 (
            .O(N__16123),
            .I(G_28_cascade_));
    InMux I__1994 (
            .O(N__16120),
            .I(N__16110));
    InMux I__1993 (
            .O(N__16119),
            .I(N__16110));
    InMux I__1992 (
            .O(N__16118),
            .I(N__16110));
    InMux I__1991 (
            .O(N__16117),
            .I(N__16107));
    LocalMux I__1990 (
            .O(N__16110),
            .I(N__16104));
    LocalMux I__1989 (
            .O(N__16107),
            .I(\POWERLED.count_clkZ0Z_7 ));
    Odrv12 I__1988 (
            .O(N__16104),
            .I(\POWERLED.count_clkZ0Z_7 ));
    CascadeMux I__1987 (
            .O(N__16099),
            .I(N__16096));
    InMux I__1986 (
            .O(N__16096),
            .I(N__16090));
    InMux I__1985 (
            .O(N__16095),
            .I(N__16090));
    LocalMux I__1984 (
            .O(N__16090),
            .I(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ));
    InMux I__1983 (
            .O(N__16087),
            .I(N__16084));
    LocalMux I__1982 (
            .O(N__16084),
            .I(\POWERLED.count_clk_0_7 ));
    InMux I__1981 (
            .O(N__16081),
            .I(N__16078));
    LocalMux I__1980 (
            .O(N__16078),
            .I(N__16075));
    Odrv4 I__1979 (
            .O(N__16075),
            .I(vpp_ok));
    IoInMux I__1978 (
            .O(N__16072),
            .I(N__16069));
    LocalMux I__1977 (
            .O(N__16069),
            .I(N__16066));
    Span4Mux_s3_v I__1976 (
            .O(N__16066),
            .I(N__16063));
    Odrv4 I__1975 (
            .O(N__16063),
            .I(vddq_en));
    InMux I__1974 (
            .O(N__16060),
            .I(N__16056));
    InMux I__1973 (
            .O(N__16059),
            .I(N__16053));
    LocalMux I__1972 (
            .O(N__16056),
            .I(\COUNTER.counterZ0Z_8 ));
    LocalMux I__1971 (
            .O(N__16053),
            .I(\COUNTER.counterZ0Z_8 ));
    InMux I__1970 (
            .O(N__16048),
            .I(N__16044));
    InMux I__1969 (
            .O(N__16047),
            .I(N__16041));
    LocalMux I__1968 (
            .O(N__16044),
            .I(\COUNTER.counterZ0Z_11 ));
    LocalMux I__1967 (
            .O(N__16041),
            .I(\COUNTER.counterZ0Z_11 ));
    CascadeMux I__1966 (
            .O(N__16036),
            .I(N__16032));
    InMux I__1965 (
            .O(N__16035),
            .I(N__16029));
    InMux I__1964 (
            .O(N__16032),
            .I(N__16026));
    LocalMux I__1963 (
            .O(N__16029),
            .I(\COUNTER.counterZ0Z_10 ));
    LocalMux I__1962 (
            .O(N__16026),
            .I(\COUNTER.counterZ0Z_10 ));
    InMux I__1961 (
            .O(N__16021),
            .I(N__16017));
    InMux I__1960 (
            .O(N__16020),
            .I(N__16014));
    LocalMux I__1959 (
            .O(N__16017),
            .I(\COUNTER.counterZ0Z_9 ));
    LocalMux I__1958 (
            .O(N__16014),
            .I(\COUNTER.counterZ0Z_9 ));
    InMux I__1957 (
            .O(N__16009),
            .I(N__16005));
    InMux I__1956 (
            .O(N__16008),
            .I(N__16002));
    LocalMux I__1955 (
            .O(N__16005),
            .I(\COUNTER.counterZ0Z_14 ));
    LocalMux I__1954 (
            .O(N__16002),
            .I(\COUNTER.counterZ0Z_14 ));
    InMux I__1953 (
            .O(N__15997),
            .I(N__15993));
    InMux I__1952 (
            .O(N__15996),
            .I(N__15990));
    LocalMux I__1951 (
            .O(N__15993),
            .I(\COUNTER.counterZ0Z_13 ));
    LocalMux I__1950 (
            .O(N__15990),
            .I(\COUNTER.counterZ0Z_13 ));
    CascadeMux I__1949 (
            .O(N__15985),
            .I(N__15981));
    InMux I__1948 (
            .O(N__15984),
            .I(N__15978));
    InMux I__1947 (
            .O(N__15981),
            .I(N__15975));
    LocalMux I__1946 (
            .O(N__15978),
            .I(\COUNTER.counterZ0Z_15 ));
    LocalMux I__1945 (
            .O(N__15975),
            .I(\COUNTER.counterZ0Z_15 ));
    InMux I__1944 (
            .O(N__15970),
            .I(N__15966));
    InMux I__1943 (
            .O(N__15969),
            .I(N__15963));
    LocalMux I__1942 (
            .O(N__15966),
            .I(\COUNTER.counterZ0Z_12 ));
    LocalMux I__1941 (
            .O(N__15963),
            .I(\COUNTER.counterZ0Z_12 ));
    InMux I__1940 (
            .O(N__15958),
            .I(N__15954));
    InMux I__1939 (
            .O(N__15957),
            .I(N__15951));
    LocalMux I__1938 (
            .O(N__15954),
            .I(\COUNTER.counterZ0Z_18 ));
    LocalMux I__1937 (
            .O(N__15951),
            .I(\COUNTER.counterZ0Z_18 ));
    InMux I__1936 (
            .O(N__15946),
            .I(N__15942));
    InMux I__1935 (
            .O(N__15945),
            .I(N__15939));
    LocalMux I__1934 (
            .O(N__15942),
            .I(\COUNTER.counterZ0Z_17 ));
    LocalMux I__1933 (
            .O(N__15939),
            .I(\COUNTER.counterZ0Z_17 ));
    CascadeMux I__1932 (
            .O(N__15934),
            .I(N__15930));
    InMux I__1931 (
            .O(N__15933),
            .I(N__15927));
    InMux I__1930 (
            .O(N__15930),
            .I(N__15924));
    LocalMux I__1929 (
            .O(N__15927),
            .I(\COUNTER.counterZ0Z_19 ));
    LocalMux I__1928 (
            .O(N__15924),
            .I(\COUNTER.counterZ0Z_19 ));
    InMux I__1927 (
            .O(N__15919),
            .I(N__15915));
    InMux I__1926 (
            .O(N__15918),
            .I(N__15912));
    LocalMux I__1925 (
            .O(N__15915),
            .I(\COUNTER.counterZ0Z_16 ));
    LocalMux I__1924 (
            .O(N__15912),
            .I(\COUNTER.counterZ0Z_16 ));
    InMux I__1923 (
            .O(N__15907),
            .I(N__15892));
    InMux I__1922 (
            .O(N__15906),
            .I(N__15892));
    InMux I__1921 (
            .O(N__15905),
            .I(N__15892));
    InMux I__1920 (
            .O(N__15904),
            .I(N__15892));
    InMux I__1919 (
            .O(N__15903),
            .I(N__15885));
    InMux I__1918 (
            .O(N__15902),
            .I(N__15885));
    InMux I__1917 (
            .O(N__15901),
            .I(N__15885));
    LocalMux I__1916 (
            .O(N__15892),
            .I(N__15879));
    LocalMux I__1915 (
            .O(N__15885),
            .I(N__15876));
    InMux I__1914 (
            .O(N__15884),
            .I(N__15866));
    InMux I__1913 (
            .O(N__15883),
            .I(N__15863));
    InMux I__1912 (
            .O(N__15882),
            .I(N__15860));
    Span4Mux_s2_h I__1911 (
            .O(N__15879),
            .I(N__15855));
    Span4Mux_s2_h I__1910 (
            .O(N__15876),
            .I(N__15855));
    InMux I__1909 (
            .O(N__15875),
            .I(N__15848));
    InMux I__1908 (
            .O(N__15874),
            .I(N__15848));
    InMux I__1907 (
            .O(N__15873),
            .I(N__15848));
    InMux I__1906 (
            .O(N__15872),
            .I(N__15839));
    InMux I__1905 (
            .O(N__15871),
            .I(N__15839));
    InMux I__1904 (
            .O(N__15870),
            .I(N__15839));
    InMux I__1903 (
            .O(N__15869),
            .I(N__15839));
    LocalMux I__1902 (
            .O(N__15866),
            .I(\POWERLED.N_47_i ));
    LocalMux I__1901 (
            .O(N__15863),
            .I(\POWERLED.N_47_i ));
    LocalMux I__1900 (
            .O(N__15860),
            .I(\POWERLED.N_47_i ));
    Odrv4 I__1899 (
            .O(N__15855),
            .I(\POWERLED.N_47_i ));
    LocalMux I__1898 (
            .O(N__15848),
            .I(\POWERLED.N_47_i ));
    LocalMux I__1897 (
            .O(N__15839),
            .I(\POWERLED.N_47_i ));
    InMux I__1896 (
            .O(N__15826),
            .I(N__15819));
    InMux I__1895 (
            .O(N__15825),
            .I(N__15814));
    InMux I__1894 (
            .O(N__15824),
            .I(N__15814));
    InMux I__1893 (
            .O(N__15823),
            .I(N__15811));
    InMux I__1892 (
            .O(N__15822),
            .I(N__15808));
    LocalMux I__1891 (
            .O(N__15819),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__1890 (
            .O(N__15814),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__1889 (
            .O(N__15811),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__1888 (
            .O(N__15808),
            .I(\POWERLED.count_clkZ0Z_0 ));
    InMux I__1887 (
            .O(N__15799),
            .I(N__15796));
    LocalMux I__1886 (
            .O(N__15796),
            .I(\POWERLED.count_clk_0_1 ));
    CascadeMux I__1885 (
            .O(N__15793),
            .I(\POWERLED.count_clk_RNIZ0Z_0_cascade_ ));
    CascadeMux I__1884 (
            .O(N__15790),
            .I(N__15786));
    InMux I__1883 (
            .O(N__15789),
            .I(N__15780));
    InMux I__1882 (
            .O(N__15786),
            .I(N__15777));
    InMux I__1881 (
            .O(N__15785),
            .I(N__15770));
    InMux I__1880 (
            .O(N__15784),
            .I(N__15770));
    InMux I__1879 (
            .O(N__15783),
            .I(N__15770));
    LocalMux I__1878 (
            .O(N__15780),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__1877 (
            .O(N__15777),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__1876 (
            .O(N__15770),
            .I(\POWERLED.count_clkZ0Z_1 ));
    InMux I__1875 (
            .O(N__15763),
            .I(N__15757));
    InMux I__1874 (
            .O(N__15762),
            .I(N__15757));
    LocalMux I__1873 (
            .O(N__15757),
            .I(\POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ));
    CascadeMux I__1872 (
            .O(N__15754),
            .I(N__15751));
    InMux I__1871 (
            .O(N__15751),
            .I(N__15748));
    LocalMux I__1870 (
            .O(N__15748),
            .I(\POWERLED.count_clk_0_9 ));
    InMux I__1869 (
            .O(N__15745),
            .I(N__15739));
    InMux I__1868 (
            .O(N__15744),
            .I(N__15739));
    LocalMux I__1867 (
            .O(N__15739),
            .I(N__15735));
    InMux I__1866 (
            .O(N__15738),
            .I(N__15732));
    Odrv12 I__1865 (
            .O(N__15735),
            .I(\POWERLED.count_clkZ0Z_6 ));
    LocalMux I__1864 (
            .O(N__15732),
            .I(\POWERLED.count_clkZ0Z_6 ));
    InMux I__1863 (
            .O(N__15727),
            .I(N__15721));
    InMux I__1862 (
            .O(N__15726),
            .I(N__15721));
    LocalMux I__1861 (
            .O(N__15721),
            .I(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ));
    CascadeMux I__1860 (
            .O(N__15718),
            .I(N__15715));
    InMux I__1859 (
            .O(N__15715),
            .I(N__15712));
    LocalMux I__1858 (
            .O(N__15712),
            .I(\POWERLED.count_clk_0_6 ));
    CascadeMux I__1857 (
            .O(N__15709),
            .I(N__15705));
    InMux I__1856 (
            .O(N__15708),
            .I(N__15700));
    InMux I__1855 (
            .O(N__15705),
            .I(N__15700));
    LocalMux I__1854 (
            .O(N__15700),
            .I(N__15696));
    InMux I__1853 (
            .O(N__15699),
            .I(N__15693));
    Odrv4 I__1852 (
            .O(N__15696),
            .I(\POWERLED.count_clkZ0Z_8 ));
    LocalMux I__1851 (
            .O(N__15693),
            .I(\POWERLED.count_clkZ0Z_8 ));
    InMux I__1850 (
            .O(N__15688),
            .I(N__15682));
    InMux I__1849 (
            .O(N__15687),
            .I(N__15682));
    LocalMux I__1848 (
            .O(N__15682),
            .I(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ));
    CascadeMux I__1847 (
            .O(N__15679),
            .I(N__15676));
    InMux I__1846 (
            .O(N__15676),
            .I(N__15673));
    LocalMux I__1845 (
            .O(N__15673),
            .I(\POWERLED.count_clk_0_8 ));
    InMux I__1844 (
            .O(N__15670),
            .I(N__15664));
    InMux I__1843 (
            .O(N__15669),
            .I(N__15664));
    LocalMux I__1842 (
            .O(N__15664),
            .I(N__15660));
    InMux I__1841 (
            .O(N__15663),
            .I(N__15657));
    Odrv4 I__1840 (
            .O(N__15660),
            .I(\POWERLED.count_clkZ0Z_2 ));
    LocalMux I__1839 (
            .O(N__15657),
            .I(\POWERLED.count_clkZ0Z_2 ));
    InMux I__1838 (
            .O(N__15652),
            .I(N__15646));
    InMux I__1837 (
            .O(N__15651),
            .I(N__15646));
    LocalMux I__1836 (
            .O(N__15646),
            .I(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ));
    CascadeMux I__1835 (
            .O(N__15643),
            .I(N__15640));
    InMux I__1834 (
            .O(N__15640),
            .I(N__15637));
    LocalMux I__1833 (
            .O(N__15637),
            .I(\POWERLED.count_clk_0_2 ));
    InMux I__1832 (
            .O(N__15634),
            .I(N__15631));
    LocalMux I__1831 (
            .O(N__15631),
            .I(\POWERLED.count_clk_0_0 ));
    InMux I__1830 (
            .O(N__15628),
            .I(N__15625));
    LocalMux I__1829 (
            .O(N__15625),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_i_i_0 ));
    InMux I__1828 (
            .O(N__15622),
            .I(N__15619));
    LocalMux I__1827 (
            .O(N__15619),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_i_i_1 ));
    InMux I__1826 (
            .O(N__15616),
            .I(N__15613));
    LocalMux I__1825 (
            .O(N__15613),
            .I(\POWERLED.N_415 ));
    InMux I__1824 (
            .O(N__15610),
            .I(N__15607));
    LocalMux I__1823 (
            .O(N__15607),
            .I(N__15603));
    InMux I__1822 (
            .O(N__15606),
            .I(N__15600));
    Odrv4 I__1821 (
            .O(N__15603),
            .I(\POWERLED.count_clkZ0Z_9 ));
    LocalMux I__1820 (
            .O(N__15600),
            .I(\POWERLED.count_clkZ0Z_9 ));
    CascadeMux I__1819 (
            .O(N__15595),
            .I(\POWERLED.count_clkZ0Z_9_cascade_ ));
    InMux I__1818 (
            .O(N__15592),
            .I(N__15586));
    InMux I__1817 (
            .O(N__15591),
            .I(N__15586));
    LocalMux I__1816 (
            .O(N__15586),
            .I(N__15583));
    Odrv4 I__1815 (
            .O(N__15583),
            .I(\POWERLED.N_320 ));
    InMux I__1814 (
            .O(N__15580),
            .I(N__15576));
    InMux I__1813 (
            .O(N__15579),
            .I(N__15573));
    LocalMux I__1812 (
            .O(N__15576),
            .I(\POWERLED.count_clkZ0Z_5 ));
    LocalMux I__1811 (
            .O(N__15573),
            .I(\POWERLED.count_clkZ0Z_5 ));
    InMux I__1810 (
            .O(N__15568),
            .I(N__15562));
    InMux I__1809 (
            .O(N__15567),
            .I(N__15562));
    LocalMux I__1808 (
            .O(N__15562),
            .I(\POWERLED.N_289 ));
    CascadeMux I__1807 (
            .O(N__15559),
            .I(\POWERLED.count_clkZ0Z_5_cascade_ ));
    InMux I__1806 (
            .O(N__15556),
            .I(N__15553));
    LocalMux I__1805 (
            .O(N__15553),
            .I(N__15550));
    Odrv4 I__1804 (
            .O(N__15550),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_i_i_a2_1_2 ));
    InMux I__1803 (
            .O(N__15547),
            .I(N__15541));
    InMux I__1802 (
            .O(N__15546),
            .I(N__15541));
    LocalMux I__1801 (
            .O(N__15541),
            .I(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ));
    CascadeMux I__1800 (
            .O(N__15538),
            .I(N__15535));
    InMux I__1799 (
            .O(N__15535),
            .I(N__15532));
    LocalMux I__1798 (
            .O(N__15532),
            .I(\POWERLED.count_clk_0_5 ));
    InMux I__1797 (
            .O(N__15529),
            .I(N__15523));
    InMux I__1796 (
            .O(N__15528),
            .I(N__15523));
    LocalMux I__1795 (
            .O(N__15523),
            .I(N__15520));
    Odrv4 I__1794 (
            .O(N__15520),
            .I(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ));
    CascadeMux I__1793 (
            .O(N__15517),
            .I(N__15514));
    InMux I__1792 (
            .O(N__15514),
            .I(N__15511));
    LocalMux I__1791 (
            .O(N__15511),
            .I(\POWERLED.count_clk_0_3 ));
    InMux I__1790 (
            .O(N__15508),
            .I(N__15504));
    InMux I__1789 (
            .O(N__15507),
            .I(N__15501));
    LocalMux I__1788 (
            .O(N__15504),
            .I(N__15498));
    LocalMux I__1787 (
            .O(N__15501),
            .I(N__15495));
    Span4Mux_v I__1786 (
            .O(N__15498),
            .I(N__15492));
    Odrv4 I__1785 (
            .O(N__15495),
            .I(\POWERLED.count_clkZ0Z_3 ));
    Odrv4 I__1784 (
            .O(N__15492),
            .I(\POWERLED.count_clkZ0Z_3 ));
    CascadeMux I__1783 (
            .O(N__15487),
            .I(\POWERLED.count_clkZ0Z_3_cascade_ ));
    CascadeMux I__1782 (
            .O(N__15484),
            .I(N__15481));
    InMux I__1781 (
            .O(N__15481),
            .I(N__15476));
    InMux I__1780 (
            .O(N__15480),
            .I(N__15471));
    InMux I__1779 (
            .O(N__15479),
            .I(N__15471));
    LocalMux I__1778 (
            .O(N__15476),
            .I(N__15468));
    LocalMux I__1777 (
            .O(N__15471),
            .I(\POWERLED.count_clkZ0Z_4 ));
    Odrv4 I__1776 (
            .O(N__15468),
            .I(\POWERLED.count_clkZ0Z_4 ));
    CascadeMux I__1775 (
            .O(N__15463),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_i_i_a2_5_0_cascade_ ));
    CascadeMux I__1774 (
            .O(N__15460),
            .I(\POWERLED.N_515_cascade_ ));
    CascadeMux I__1773 (
            .O(N__15457),
            .I(N__15454));
    InMux I__1772 (
            .O(N__15454),
            .I(N__15451));
    LocalMux I__1771 (
            .O(N__15451),
            .I(\POWERLED.N_515 ));
    CascadeMux I__1770 (
            .O(N__15448),
            .I(\POWERLED.N_47_i_cascade_ ));
    CascadeMux I__1769 (
            .O(N__15445),
            .I(\POWERLED.count_clk_RNI_0Z0Z_0_cascade_ ));
    CascadeMux I__1768 (
            .O(N__15442),
            .I(\POWERLED.count_clkZ0Z_0_cascade_ ));
    InMux I__1767 (
            .O(N__15439),
            .I(N__15436));
    LocalMux I__1766 (
            .O(N__15436),
            .I(N__15433));
    Odrv4 I__1765 (
            .O(N__15433),
            .I(\HDA_STRAP.un1_count_1_cry_7_THRU_CO ));
    InMux I__1764 (
            .O(N__15430),
            .I(N__15425));
    InMux I__1763 (
            .O(N__15429),
            .I(N__15420));
    InMux I__1762 (
            .O(N__15428),
            .I(N__15420));
    LocalMux I__1761 (
            .O(N__15425),
            .I(\HDA_STRAP.countZ0Z_8 ));
    LocalMux I__1760 (
            .O(N__15420),
            .I(\HDA_STRAP.countZ0Z_8 ));
    CascadeMux I__1759 (
            .O(N__15415),
            .I(N__15409));
    CascadeMux I__1758 (
            .O(N__15414),
            .I(N__15404));
    CascadeMux I__1757 (
            .O(N__15413),
            .I(N__15401));
    CascadeMux I__1756 (
            .O(N__15412),
            .I(N__15396));
    InMux I__1755 (
            .O(N__15409),
            .I(N__15392));
    InMux I__1754 (
            .O(N__15408),
            .I(N__15389));
    InMux I__1753 (
            .O(N__15407),
            .I(N__15380));
    InMux I__1752 (
            .O(N__15404),
            .I(N__15380));
    InMux I__1751 (
            .O(N__15401),
            .I(N__15380));
    InMux I__1750 (
            .O(N__15400),
            .I(N__15380));
    CascadeMux I__1749 (
            .O(N__15399),
            .I(N__15377));
    InMux I__1748 (
            .O(N__15396),
            .I(N__15373));
    InMux I__1747 (
            .O(N__15395),
            .I(N__15370));
    LocalMux I__1746 (
            .O(N__15392),
            .I(N__15367));
    LocalMux I__1745 (
            .O(N__15389),
            .I(N__15362));
    LocalMux I__1744 (
            .O(N__15380),
            .I(N__15362));
    InMux I__1743 (
            .O(N__15377),
            .I(N__15357));
    InMux I__1742 (
            .O(N__15376),
            .I(N__15357));
    LocalMux I__1741 (
            .O(N__15373),
            .I(N__15354));
    LocalMux I__1740 (
            .O(N__15370),
            .I(\HDA_STRAP.curr_state_RNIH91A_0Z0Z_0 ));
    Odrv4 I__1739 (
            .O(N__15367),
            .I(\HDA_STRAP.curr_state_RNIH91A_0Z0Z_0 ));
    Odrv4 I__1738 (
            .O(N__15362),
            .I(\HDA_STRAP.curr_state_RNIH91A_0Z0Z_0 ));
    LocalMux I__1737 (
            .O(N__15357),
            .I(\HDA_STRAP.curr_state_RNIH91A_0Z0Z_0 ));
    Odrv4 I__1736 (
            .O(N__15354),
            .I(\HDA_STRAP.curr_state_RNIH91A_0Z0Z_0 ));
    CascadeMux I__1735 (
            .O(N__15343),
            .I(\HDA_STRAP.N_9_cascade_ ));
    InMux I__1734 (
            .O(N__15340),
            .I(N__15334));
    InMux I__1733 (
            .O(N__15339),
            .I(N__15334));
    LocalMux I__1732 (
            .O(N__15334),
            .I(\HDA_STRAP.N_336 ));
    InMux I__1731 (
            .O(N__15331),
            .I(N__15325));
    InMux I__1730 (
            .O(N__15330),
            .I(N__15325));
    LocalMux I__1729 (
            .O(N__15325),
            .I(\HDA_STRAP.curr_stateZ0Z_2 ));
    IoInMux I__1728 (
            .O(N__15322),
            .I(N__15319));
    LocalMux I__1727 (
            .O(N__15319),
            .I(N__15316));
    Span4Mux_s1_h I__1726 (
            .O(N__15316),
            .I(N__15313));
    Odrv4 I__1725 (
            .O(N__15313),
            .I(hda_sdo_atp));
    CascadeMux I__1724 (
            .O(N__15310),
            .I(N__15306));
    CascadeMux I__1723 (
            .O(N__15309),
            .I(N__15297));
    InMux I__1722 (
            .O(N__15306),
            .I(N__15294));
    InMux I__1721 (
            .O(N__15305),
            .I(N__15284));
    InMux I__1720 (
            .O(N__15304),
            .I(N__15284));
    InMux I__1719 (
            .O(N__15303),
            .I(N__15284));
    InMux I__1718 (
            .O(N__15302),
            .I(N__15284));
    InMux I__1717 (
            .O(N__15301),
            .I(N__15277));
    InMux I__1716 (
            .O(N__15300),
            .I(N__15277));
    InMux I__1715 (
            .O(N__15297),
            .I(N__15277));
    LocalMux I__1714 (
            .O(N__15294),
            .I(N__15274));
    InMux I__1713 (
            .O(N__15293),
            .I(N__15271));
    LocalMux I__1712 (
            .O(N__15284),
            .I(N__15268));
    LocalMux I__1711 (
            .O(N__15277),
            .I(\HDA_STRAP.un4_count ));
    Odrv12 I__1710 (
            .O(N__15274),
            .I(\HDA_STRAP.un4_count ));
    LocalMux I__1709 (
            .O(N__15271),
            .I(\HDA_STRAP.un4_count ));
    Odrv4 I__1708 (
            .O(N__15268),
            .I(\HDA_STRAP.un4_count ));
    CascadeMux I__1707 (
            .O(N__15259),
            .I(N__15256));
    InMux I__1706 (
            .O(N__15256),
            .I(N__15251));
    CascadeMux I__1705 (
            .O(N__15255),
            .I(N__15247));
    CascadeMux I__1704 (
            .O(N__15254),
            .I(N__15244));
    LocalMux I__1703 (
            .O(N__15251),
            .I(N__15240));
    InMux I__1702 (
            .O(N__15250),
            .I(N__15237));
    InMux I__1701 (
            .O(N__15247),
            .I(N__15230));
    InMux I__1700 (
            .O(N__15244),
            .I(N__15230));
    InMux I__1699 (
            .O(N__15243),
            .I(N__15230));
    Odrv12 I__1698 (
            .O(N__15240),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__1697 (
            .O(N__15237),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__1696 (
            .O(N__15230),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    InMux I__1695 (
            .O(N__15223),
            .I(N__15216));
    InMux I__1694 (
            .O(N__15222),
            .I(N__15207));
    InMux I__1693 (
            .O(N__15221),
            .I(N__15207));
    InMux I__1692 (
            .O(N__15220),
            .I(N__15207));
    InMux I__1691 (
            .O(N__15219),
            .I(N__15207));
    LocalMux I__1690 (
            .O(N__15216),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    LocalMux I__1689 (
            .O(N__15207),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    InMux I__1688 (
            .O(N__15202),
            .I(N__15199));
    LocalMux I__1687 (
            .O(N__15199),
            .I(N__15196));
    Span4Mux_v I__1686 (
            .O(N__15196),
            .I(N__15193));
    Odrv4 I__1685 (
            .O(N__15193),
            .I(vr_ready_vccin));
    CascadeMux I__1684 (
            .O(N__15190),
            .I(\POWERLED.un1_dutycycle_168_0_0_o3_4_cascade_ ));
    CascadeMux I__1683 (
            .O(N__15187),
            .I(\PCH_PWRGD.N_38_f0_cascade_ ));
    InMux I__1682 (
            .O(N__15184),
            .I(N__15181));
    LocalMux I__1681 (
            .O(N__15181),
            .I(\PCH_PWRGD.delayed_vccin_okZ0 ));
    InMux I__1680 (
            .O(N__15178),
            .I(N__15175));
    LocalMux I__1679 (
            .O(N__15175),
            .I(N__15172));
    Span4Mux_h I__1678 (
            .O(N__15172),
            .I(N__15169));
    Span4Mux_h I__1677 (
            .O(N__15169),
            .I(N__15166));
    Span4Mux_v I__1676 (
            .O(N__15166),
            .I(N__15163));
    Odrv4 I__1675 (
            .O(N__15163),
            .I(gpio_fpga_soc_1));
    CascadeMux I__1674 (
            .O(N__15160),
            .I(\HDA_STRAP.m14_i_0_cascade_ ));
    InMux I__1673 (
            .O(N__15157),
            .I(N__15153));
    InMux I__1672 (
            .O(N__15156),
            .I(N__15150));
    LocalMux I__1671 (
            .O(N__15153),
            .I(\HDA_STRAP.countZ0Z_13 ));
    LocalMux I__1670 (
            .O(N__15150),
            .I(\HDA_STRAP.countZ0Z_13 ));
    InMux I__1669 (
            .O(N__15145),
            .I(N__15141));
    InMux I__1668 (
            .O(N__15144),
            .I(N__15138));
    LocalMux I__1667 (
            .O(N__15141),
            .I(\HDA_STRAP.countZ0Z_9 ));
    LocalMux I__1666 (
            .O(N__15138),
            .I(\HDA_STRAP.countZ0Z_9 ));
    CascadeMux I__1665 (
            .O(N__15133),
            .I(N__15129));
    InMux I__1664 (
            .O(N__15132),
            .I(N__15126));
    InMux I__1663 (
            .O(N__15129),
            .I(N__15123));
    LocalMux I__1662 (
            .O(N__15126),
            .I(\HDA_STRAP.countZ0Z_12 ));
    LocalMux I__1661 (
            .O(N__15123),
            .I(\HDA_STRAP.countZ0Z_12 ));
    InMux I__1660 (
            .O(N__15118),
            .I(N__15114));
    InMux I__1659 (
            .O(N__15117),
            .I(N__15111));
    LocalMux I__1658 (
            .O(N__15114),
            .I(\HDA_STRAP.countZ0Z_7 ));
    LocalMux I__1657 (
            .O(N__15111),
            .I(\HDA_STRAP.countZ0Z_7 ));
    InMux I__1656 (
            .O(N__15106),
            .I(N__15103));
    LocalMux I__1655 (
            .O(N__15103),
            .I(N__15100));
    Span4Mux_v I__1654 (
            .O(N__15100),
            .I(N__15097));
    Odrv4 I__1653 (
            .O(N__15097),
            .I(\HDA_STRAP.un4_count_11 ));
    InMux I__1652 (
            .O(N__15094),
            .I(N__15090));
    InMux I__1651 (
            .O(N__15093),
            .I(N__15087));
    LocalMux I__1650 (
            .O(N__15090),
            .I(\HDA_STRAP.countZ0Z_14 ));
    LocalMux I__1649 (
            .O(N__15087),
            .I(\HDA_STRAP.countZ0Z_14 ));
    InMux I__1648 (
            .O(N__15082),
            .I(N__15078));
    InMux I__1647 (
            .O(N__15081),
            .I(N__15075));
    LocalMux I__1646 (
            .O(N__15078),
            .I(\HDA_STRAP.countZ0Z_15 ));
    LocalMux I__1645 (
            .O(N__15075),
            .I(\HDA_STRAP.countZ0Z_15 ));
    InMux I__1644 (
            .O(N__15070),
            .I(N__15067));
    LocalMux I__1643 (
            .O(N__15067),
            .I(N__15064));
    Odrv4 I__1642 (
            .O(N__15064),
            .I(\HDA_STRAP.un4_count_12 ));
    InMux I__1641 (
            .O(N__15061),
            .I(N__15058));
    LocalMux I__1640 (
            .O(N__15058),
            .I(\HDA_STRAP.un1_count_1_cry_5_THRU_CO ));
    CascadeMux I__1639 (
            .O(N__15055),
            .I(N__15051));
    InMux I__1638 (
            .O(N__15054),
            .I(N__15045));
    InMux I__1637 (
            .O(N__15051),
            .I(N__15045));
    InMux I__1636 (
            .O(N__15050),
            .I(N__15042));
    LocalMux I__1635 (
            .O(N__15045),
            .I(\HDA_STRAP.countZ0Z_6 ));
    LocalMux I__1634 (
            .O(N__15042),
            .I(\HDA_STRAP.countZ0Z_6 ));
    InMux I__1633 (
            .O(N__15037),
            .I(N__15034));
    LocalMux I__1632 (
            .O(N__15034),
            .I(\PCH_PWRGD.curr_state_0_0 ));
    CascadeMux I__1631 (
            .O(N__15031),
            .I(\PCH_PWRGD.curr_state_7_0_cascade_ ));
    CascadeMux I__1630 (
            .O(N__15028),
            .I(\PCH_PWRGD.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__1629 (
            .O(N__15025),
            .I(N__15021));
    CascadeMux I__1628 (
            .O(N__15024),
            .I(N__15018));
    InMux I__1627 (
            .O(N__15021),
            .I(N__15012));
    InMux I__1626 (
            .O(N__15018),
            .I(N__15012));
    InMux I__1625 (
            .O(N__15017),
            .I(N__15000));
    LocalMux I__1624 (
            .O(N__15012),
            .I(N__14992));
    InMux I__1623 (
            .O(N__15011),
            .I(N__14983));
    InMux I__1622 (
            .O(N__15010),
            .I(N__14983));
    InMux I__1621 (
            .O(N__15009),
            .I(N__14983));
    InMux I__1620 (
            .O(N__15008),
            .I(N__14983));
    InMux I__1619 (
            .O(N__15007),
            .I(N__14974));
    InMux I__1618 (
            .O(N__15006),
            .I(N__14974));
    InMux I__1617 (
            .O(N__15005),
            .I(N__14974));
    InMux I__1616 (
            .O(N__15004),
            .I(N__14974));
    InMux I__1615 (
            .O(N__15003),
            .I(N__14971));
    LocalMux I__1614 (
            .O(N__15000),
            .I(N__14968));
    InMux I__1613 (
            .O(N__14999),
            .I(N__14957));
    InMux I__1612 (
            .O(N__14998),
            .I(N__14957));
    InMux I__1611 (
            .O(N__14997),
            .I(N__14957));
    InMux I__1610 (
            .O(N__14996),
            .I(N__14957));
    InMux I__1609 (
            .O(N__14995),
            .I(N__14957));
    Span4Mux_v I__1608 (
            .O(N__14992),
            .I(N__14950));
    LocalMux I__1607 (
            .O(N__14983),
            .I(N__14950));
    LocalMux I__1606 (
            .O(N__14974),
            .I(N__14950));
    LocalMux I__1605 (
            .O(N__14971),
            .I(\PCH_PWRGD.N_540 ));
    Odrv12 I__1604 (
            .O(N__14968),
            .I(\PCH_PWRGD.N_540 ));
    LocalMux I__1603 (
            .O(N__14957),
            .I(\PCH_PWRGD.N_540 ));
    Odrv4 I__1602 (
            .O(N__14950),
            .I(\PCH_PWRGD.N_540 ));
    InMux I__1601 (
            .O(N__14941),
            .I(N__14938));
    LocalMux I__1600 (
            .O(N__14938),
            .I(\PCH_PWRGD.N_205 ));
    InMux I__1599 (
            .O(N__14935),
            .I(N__14932));
    LocalMux I__1598 (
            .O(N__14932),
            .I(\PCH_PWRGD.curr_state_0_1 ));
    CascadeMux I__1597 (
            .O(N__14929),
            .I(\PCH_PWRGD.N_205_cascade_ ));
    InMux I__1596 (
            .O(N__14926),
            .I(N__14917));
    InMux I__1595 (
            .O(N__14925),
            .I(N__14917));
    InMux I__1594 (
            .O(N__14924),
            .I(N__14917));
    LocalMux I__1593 (
            .O(N__14917),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__1592 (
            .O(N__14914),
            .I(\PCH_PWRGD.curr_stateZ0Z_1_cascade_ ));
    CascadeMux I__1591 (
            .O(N__14911),
            .I(\PCH_PWRGD.N_2110_i_cascade_ ));
    InMux I__1590 (
            .O(N__14908),
            .I(N__14904));
    InMux I__1589 (
            .O(N__14907),
            .I(N__14901));
    LocalMux I__1588 (
            .O(N__14904),
            .I(N__14898));
    LocalMux I__1587 (
            .O(N__14901),
            .I(\PCH_PWRGD.N_562 ));
    Odrv4 I__1586 (
            .O(N__14898),
            .I(\PCH_PWRGD.N_562 ));
    CascadeMux I__1585 (
            .O(N__14893),
            .I(\PCH_PWRGD.N_562_cascade_ ));
    InMux I__1584 (
            .O(N__14890),
            .I(N__14887));
    LocalMux I__1583 (
            .O(N__14887),
            .I(\PCH_PWRGD.count_0_2 ));
    InMux I__1582 (
            .O(N__14884),
            .I(N__14878));
    InMux I__1581 (
            .O(N__14883),
            .I(N__14878));
    LocalMux I__1580 (
            .O(N__14878),
            .I(N__14875));
    Span4Mux_h I__1579 (
            .O(N__14875),
            .I(N__14872));
    Odrv4 I__1578 (
            .O(N__14872),
            .I(\PCH_PWRGD.count_rst_12 ));
    InMux I__1577 (
            .O(N__14869),
            .I(N__14866));
    LocalMux I__1576 (
            .O(N__14866),
            .I(\PCH_PWRGD.count_0_10 ));
    CascadeMux I__1575 (
            .O(N__14863),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0_cascade_ ));
    InMux I__1574 (
            .O(N__14860),
            .I(N__14854));
    InMux I__1573 (
            .O(N__14859),
            .I(N__14854));
    LocalMux I__1572 (
            .O(N__14854),
            .I(\PCH_PWRGD.count_rst_4 ));
    InMux I__1571 (
            .O(N__14851),
            .I(N__14848));
    LocalMux I__1570 (
            .O(N__14848),
            .I(\PCH_PWRGD.countZ0Z_10 ));
    InMux I__1569 (
            .O(N__14845),
            .I(N__14841));
    InMux I__1568 (
            .O(N__14844),
            .I(N__14838));
    LocalMux I__1567 (
            .O(N__14841),
            .I(N__14835));
    LocalMux I__1566 (
            .O(N__14838),
            .I(\PCH_PWRGD.countZ0Z_2 ));
    Odrv4 I__1565 (
            .O(N__14835),
            .I(\PCH_PWRGD.countZ0Z_2 ));
    InMux I__1564 (
            .O(N__14830),
            .I(N__14826));
    InMux I__1563 (
            .O(N__14829),
            .I(N__14823));
    LocalMux I__1562 (
            .O(N__14826),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    LocalMux I__1561 (
            .O(N__14823),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    CascadeMux I__1560 (
            .O(N__14818),
            .I(\PCH_PWRGD.countZ0Z_10_cascade_ ));
    InMux I__1559 (
            .O(N__14815),
            .I(N__14811));
    InMux I__1558 (
            .O(N__14814),
            .I(N__14808));
    LocalMux I__1557 (
            .O(N__14811),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    LocalMux I__1556 (
            .O(N__14808),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    InMux I__1555 (
            .O(N__14803),
            .I(N__14798));
    InMux I__1554 (
            .O(N__14802),
            .I(N__14794));
    InMux I__1553 (
            .O(N__14801),
            .I(N__14791));
    LocalMux I__1552 (
            .O(N__14798),
            .I(N__14788));
    InMux I__1551 (
            .O(N__14797),
            .I(N__14785));
    LocalMux I__1550 (
            .O(N__14794),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    LocalMux I__1549 (
            .O(N__14791),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    Odrv4 I__1548 (
            .O(N__14788),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    LocalMux I__1547 (
            .O(N__14785),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    InMux I__1546 (
            .O(N__14776),
            .I(N__14772));
    InMux I__1545 (
            .O(N__14775),
            .I(N__14768));
    LocalMux I__1544 (
            .O(N__14772),
            .I(N__14765));
    InMux I__1543 (
            .O(N__14771),
            .I(N__14762));
    LocalMux I__1542 (
            .O(N__14768),
            .I(N__14759));
    Odrv4 I__1541 (
            .O(N__14765),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    LocalMux I__1540 (
            .O(N__14762),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    Odrv4 I__1539 (
            .O(N__14759),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    CascadeMux I__1538 (
            .O(N__14752),
            .I(\PCH_PWRGD.count_1_i_a2_8_0_cascade_ ));
    CascadeMux I__1537 (
            .O(N__14749),
            .I(N__14744));
    InMux I__1536 (
            .O(N__14748),
            .I(N__14741));
    InMux I__1535 (
            .O(N__14747),
            .I(N__14738));
    InMux I__1534 (
            .O(N__14744),
            .I(N__14735));
    LocalMux I__1533 (
            .O(N__14741),
            .I(N__14732));
    LocalMux I__1532 (
            .O(N__14738),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    LocalMux I__1531 (
            .O(N__14735),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    Odrv4 I__1530 (
            .O(N__14732),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    InMux I__1529 (
            .O(N__14725),
            .I(N__14716));
    InMux I__1528 (
            .O(N__14724),
            .I(N__14716));
    InMux I__1527 (
            .O(N__14723),
            .I(N__14716));
    LocalMux I__1526 (
            .O(N__14716),
            .I(N__14713));
    Odrv12 I__1525 (
            .O(N__14713),
            .I(\PCH_PWRGD.count_1_i_a2_11_0 ));
    InMux I__1524 (
            .O(N__14710),
            .I(N__14706));
    InMux I__1523 (
            .O(N__14709),
            .I(N__14703));
    LocalMux I__1522 (
            .O(N__14706),
            .I(\PCH_PWRGD.count_rst_2 ));
    LocalMux I__1521 (
            .O(N__14703),
            .I(\PCH_PWRGD.count_rst_2 ));
    CascadeMux I__1520 (
            .O(N__14698),
            .I(N__14695));
    InMux I__1519 (
            .O(N__14695),
            .I(N__14692));
    LocalMux I__1518 (
            .O(N__14692),
            .I(\PCH_PWRGD.count_0_12 ));
    InMux I__1517 (
            .O(N__14689),
            .I(N__14685));
    InMux I__1516 (
            .O(N__14688),
            .I(N__14682));
    LocalMux I__1515 (
            .O(N__14685),
            .I(\PCH_PWRGD.un2_count_1_axb_11 ));
    LocalMux I__1514 (
            .O(N__14682),
            .I(\PCH_PWRGD.un2_count_1_axb_11 ));
    InMux I__1513 (
            .O(N__14677),
            .I(N__14673));
    InMux I__1512 (
            .O(N__14676),
            .I(N__14670));
    LocalMux I__1511 (
            .O(N__14673),
            .I(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ));
    LocalMux I__1510 (
            .O(N__14670),
            .I(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ));
    CascadeMux I__1509 (
            .O(N__14665),
            .I(N__14662));
    InMux I__1508 (
            .O(N__14662),
            .I(N__14656));
    InMux I__1507 (
            .O(N__14661),
            .I(N__14656));
    LocalMux I__1506 (
            .O(N__14656),
            .I(\PCH_PWRGD.count_rst_3 ));
    CascadeMux I__1505 (
            .O(N__14653),
            .I(N__14650));
    InMux I__1504 (
            .O(N__14650),
            .I(N__14646));
    InMux I__1503 (
            .O(N__14649),
            .I(N__14643));
    LocalMux I__1502 (
            .O(N__14646),
            .I(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ));
    LocalMux I__1501 (
            .O(N__14643),
            .I(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ));
    CascadeMux I__1500 (
            .O(N__14638),
            .I(\PCH_PWRGD.count_rst_9_cascade_ ));
    InMux I__1499 (
            .O(N__14635),
            .I(N__14632));
    LocalMux I__1498 (
            .O(N__14632),
            .I(N__14629));
    Odrv4 I__1497 (
            .O(N__14629),
            .I(\PCH_PWRGD.count_0_5 ));
    CascadeMux I__1496 (
            .O(N__14626),
            .I(\PCH_PWRGD.count_rst_5_cascade_ ));
    CascadeMux I__1495 (
            .O(N__14623),
            .I(N__14620));
    InMux I__1494 (
            .O(N__14620),
            .I(N__14615));
    InMux I__1493 (
            .O(N__14619),
            .I(N__14612));
    InMux I__1492 (
            .O(N__14618),
            .I(N__14609));
    LocalMux I__1491 (
            .O(N__14615),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    LocalMux I__1490 (
            .O(N__14612),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    LocalMux I__1489 (
            .O(N__14609),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    InMux I__1488 (
            .O(N__14602),
            .I(N__14596));
    InMux I__1487 (
            .O(N__14601),
            .I(N__14596));
    LocalMux I__1486 (
            .O(N__14596),
            .I(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ));
    CascadeMux I__1485 (
            .O(N__14593),
            .I(\PCH_PWRGD.countZ0Z_9_cascade_ ));
    InMux I__1484 (
            .O(N__14590),
            .I(N__14587));
    LocalMux I__1483 (
            .O(N__14587),
            .I(\PCH_PWRGD.count_0_9 ));
    CascadeMux I__1482 (
            .O(N__14584),
            .I(\PCH_PWRGD.N_2093_i_cascade_ ));
    InMux I__1481 (
            .O(N__14581),
            .I(N__14578));
    LocalMux I__1480 (
            .O(N__14578),
            .I(N__14574));
    InMux I__1479 (
            .O(N__14577),
            .I(N__14571));
    Odrv4 I__1478 (
            .O(N__14574),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    LocalMux I__1477 (
            .O(N__14571),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    InMux I__1476 (
            .O(N__14566),
            .I(N__14562));
    InMux I__1475 (
            .O(N__14565),
            .I(N__14559));
    LocalMux I__1474 (
            .O(N__14562),
            .I(\PCH_PWRGD.count_0_1 ));
    LocalMux I__1473 (
            .O(N__14559),
            .I(\PCH_PWRGD.count_0_1 ));
    CascadeMux I__1472 (
            .O(N__14554),
            .I(N__14551));
    InMux I__1471 (
            .O(N__14551),
            .I(N__14548));
    LocalMux I__1470 (
            .O(N__14548),
            .I(\PCH_PWRGD.count_rst_13 ));
    InMux I__1469 (
            .O(N__14545),
            .I(N__14542));
    LocalMux I__1468 (
            .O(N__14542),
            .I(\PCH_PWRGD.count_1_i_a2_3_0 ));
    InMux I__1467 (
            .O(N__14539),
            .I(N__14536));
    LocalMux I__1466 (
            .O(N__14536),
            .I(\PCH_PWRGD.count_1_i_a2_6_0 ));
    CascadeMux I__1465 (
            .O(N__14533),
            .I(\PCH_PWRGD.count_1_i_a2_4_0_cascade_ ));
    InMux I__1464 (
            .O(N__14530),
            .I(N__14521));
    InMux I__1463 (
            .O(N__14529),
            .I(N__14521));
    InMux I__1462 (
            .O(N__14528),
            .I(N__14521));
    LocalMux I__1461 (
            .O(N__14521),
            .I(\PCH_PWRGD.count_1_i_a2_12_0 ));
    CascadeMux I__1460 (
            .O(N__14518),
            .I(N__14515));
    InMux I__1459 (
            .O(N__14515),
            .I(N__14508));
    InMux I__1458 (
            .O(N__14514),
            .I(N__14508));
    InMux I__1457 (
            .O(N__14513),
            .I(N__14505));
    LocalMux I__1456 (
            .O(N__14508),
            .I(\PCH_PWRGD.count_rst_0 ));
    LocalMux I__1455 (
            .O(N__14505),
            .I(\PCH_PWRGD.count_rst_0 ));
    InMux I__1454 (
            .O(N__14500),
            .I(N__14496));
    InMux I__1453 (
            .O(N__14499),
            .I(N__14493));
    LocalMux I__1452 (
            .O(N__14496),
            .I(\PCH_PWRGD.count_0_14 ));
    LocalMux I__1451 (
            .O(N__14493),
            .I(\PCH_PWRGD.count_0_14 ));
    InMux I__1450 (
            .O(N__14488),
            .I(N__14485));
    LocalMux I__1449 (
            .O(N__14485),
            .I(\PCH_PWRGD.count_1_i_a2_5_0 ));
    CascadeMux I__1448 (
            .O(N__14482),
            .I(\PCH_PWRGD.un2_count_1_axb_11_cascade_ ));
    InMux I__1447 (
            .O(N__14479),
            .I(N__14473));
    InMux I__1446 (
            .O(N__14478),
            .I(N__14473));
    LocalMux I__1445 (
            .O(N__14473),
            .I(\PCH_PWRGD.count_0_11 ));
    InMux I__1444 (
            .O(N__14470),
            .I(\COUNTER.counter_1_cry_29 ));
    InMux I__1443 (
            .O(N__14467),
            .I(\COUNTER.counter_1_cry_30 ));
    CascadeMux I__1442 (
            .O(N__14464),
            .I(\PCH_PWRGD.count_rst_13_cascade_ ));
    InMux I__1441 (
            .O(N__14461),
            .I(N__14457));
    InMux I__1440 (
            .O(N__14460),
            .I(N__14454));
    LocalMux I__1439 (
            .O(N__14457),
            .I(\PCH_PWRGD.un2_count_1_axb_1 ));
    LocalMux I__1438 (
            .O(N__14454),
            .I(\PCH_PWRGD.un2_count_1_axb_1 ));
    CascadeMux I__1437 (
            .O(N__14449),
            .I(\PCH_PWRGD.un2_count_1_axb_1_cascade_ ));
    CascadeMux I__1436 (
            .O(N__14446),
            .I(\PCH_PWRGD.count_RNI6HKKGZ0Z_1_cascade_ ));
    InMux I__1435 (
            .O(N__14443),
            .I(N__14440));
    LocalMux I__1434 (
            .O(N__14440),
            .I(\PCH_PWRGD.count_0_0 ));
    CascadeMux I__1433 (
            .O(N__14437),
            .I(N__14434));
    InMux I__1432 (
            .O(N__14434),
            .I(N__14429));
    InMux I__1431 (
            .O(N__14433),
            .I(N__14424));
    InMux I__1430 (
            .O(N__14432),
            .I(N__14424));
    LocalMux I__1429 (
            .O(N__14429),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    LocalMux I__1428 (
            .O(N__14424),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    CascadeMux I__1427 (
            .O(N__14419),
            .I(\PCH_PWRGD.countZ0Z_0_cascade_ ));
    CascadeMux I__1426 (
            .O(N__14416),
            .I(N__14412));
    CascadeMux I__1425 (
            .O(N__14415),
            .I(N__14409));
    InMux I__1424 (
            .O(N__14412),
            .I(N__14404));
    InMux I__1423 (
            .O(N__14409),
            .I(N__14404));
    LocalMux I__1422 (
            .O(N__14404),
            .I(\PCH_PWRGD.N_2093_i ));
    InMux I__1421 (
            .O(N__14401),
            .I(\COUNTER.counter_1_cry_19 ));
    InMux I__1420 (
            .O(N__14398),
            .I(\COUNTER.counter_1_cry_20 ));
    InMux I__1419 (
            .O(N__14395),
            .I(\COUNTER.counter_1_cry_21 ));
    InMux I__1418 (
            .O(N__14392),
            .I(\COUNTER.counter_1_cry_22 ));
    InMux I__1417 (
            .O(N__14389),
            .I(\COUNTER.counter_1_cry_23 ));
    InMux I__1416 (
            .O(N__14386),
            .I(bfn_1_16_0_));
    InMux I__1415 (
            .O(N__14383),
            .I(\COUNTER.counter_1_cry_25 ));
    InMux I__1414 (
            .O(N__14380),
            .I(\COUNTER.counter_1_cry_26 ));
    InMux I__1413 (
            .O(N__14377),
            .I(\COUNTER.counter_1_cry_27 ));
    InMux I__1412 (
            .O(N__14374),
            .I(\COUNTER.counter_1_cry_28 ));
    InMux I__1411 (
            .O(N__14371),
            .I(\COUNTER.counter_1_cry_10 ));
    InMux I__1410 (
            .O(N__14368),
            .I(\COUNTER.counter_1_cry_11 ));
    InMux I__1409 (
            .O(N__14365),
            .I(\COUNTER.counter_1_cry_12 ));
    InMux I__1408 (
            .O(N__14362),
            .I(\COUNTER.counter_1_cry_13 ));
    InMux I__1407 (
            .O(N__14359),
            .I(\COUNTER.counter_1_cry_14 ));
    InMux I__1406 (
            .O(N__14356),
            .I(\COUNTER.counter_1_cry_15 ));
    InMux I__1405 (
            .O(N__14353),
            .I(bfn_1_15_0_));
    InMux I__1404 (
            .O(N__14350),
            .I(\COUNTER.counter_1_cry_17 ));
    InMux I__1403 (
            .O(N__14347),
            .I(\COUNTER.counter_1_cry_18 ));
    InMux I__1402 (
            .O(N__14344),
            .I(\COUNTER.counter_1_cry_1 ));
    InMux I__1401 (
            .O(N__14341),
            .I(\COUNTER.counter_1_cry_2 ));
    InMux I__1400 (
            .O(N__14338),
            .I(\COUNTER.counter_1_cry_3 ));
    InMux I__1399 (
            .O(N__14335),
            .I(\COUNTER.counter_1_cry_4 ));
    InMux I__1398 (
            .O(N__14332),
            .I(\COUNTER.counter_1_cry_5 ));
    InMux I__1397 (
            .O(N__14329),
            .I(\COUNTER.counter_1_cry_6 ));
    InMux I__1396 (
            .O(N__14326),
            .I(\COUNTER.counter_1_cry_7 ));
    InMux I__1395 (
            .O(N__14323),
            .I(bfn_1_14_0_));
    InMux I__1394 (
            .O(N__14320),
            .I(\COUNTER.counter_1_cry_9 ));
    CascadeMux I__1393 (
            .O(N__14317),
            .I(N__14314));
    InMux I__1392 (
            .O(N__14314),
            .I(N__14310));
    InMux I__1391 (
            .O(N__14313),
            .I(N__14307));
    LocalMux I__1390 (
            .O(N__14310),
            .I(N__14304));
    LocalMux I__1389 (
            .O(N__14307),
            .I(\POWERLED.count_clkZ0Z_10 ));
    Odrv4 I__1388 (
            .O(N__14304),
            .I(\POWERLED.count_clkZ0Z_10 ));
    InMux I__1387 (
            .O(N__14299),
            .I(N__14293));
    InMux I__1386 (
            .O(N__14298),
            .I(N__14293));
    LocalMux I__1385 (
            .O(N__14293),
            .I(N__14290));
    Odrv4 I__1384 (
            .O(N__14290),
            .I(\POWERLED.count_clk_1_10 ));
    InMux I__1383 (
            .O(N__14287),
            .I(\POWERLED.un1_count_clk_2_cry_9_cZ0 ));
    InMux I__1382 (
            .O(N__14284),
            .I(N__14280));
    InMux I__1381 (
            .O(N__14283),
            .I(N__14277));
    LocalMux I__1380 (
            .O(N__14280),
            .I(N__14274));
    LocalMux I__1379 (
            .O(N__14277),
            .I(\POWERLED.count_clkZ0Z_11 ));
    Odrv4 I__1378 (
            .O(N__14274),
            .I(\POWERLED.count_clkZ0Z_11 ));
    InMux I__1377 (
            .O(N__14269),
            .I(N__14263));
    InMux I__1376 (
            .O(N__14268),
            .I(N__14263));
    LocalMux I__1375 (
            .O(N__14263),
            .I(N__14260));
    Odrv4 I__1374 (
            .O(N__14260),
            .I(\POWERLED.count_clk_1_11 ));
    InMux I__1373 (
            .O(N__14257),
            .I(\POWERLED.un1_count_clk_2_cry_10 ));
    InMux I__1372 (
            .O(N__14254),
            .I(N__14250));
    InMux I__1371 (
            .O(N__14253),
            .I(N__14247));
    LocalMux I__1370 (
            .O(N__14250),
            .I(N__14244));
    LocalMux I__1369 (
            .O(N__14247),
            .I(\POWERLED.count_clkZ0Z_12 ));
    Odrv4 I__1368 (
            .O(N__14244),
            .I(\POWERLED.count_clkZ0Z_12 ));
    InMux I__1367 (
            .O(N__14239),
            .I(N__14233));
    InMux I__1366 (
            .O(N__14238),
            .I(N__14233));
    LocalMux I__1365 (
            .O(N__14233),
            .I(N__14230));
    Odrv4 I__1364 (
            .O(N__14230),
            .I(\POWERLED.count_clk_1_12 ));
    InMux I__1363 (
            .O(N__14227),
            .I(\POWERLED.un1_count_clk_2_cry_11 ));
    InMux I__1362 (
            .O(N__14224),
            .I(\POWERLED.un1_count_clk_2_cry_12 ));
    InMux I__1361 (
            .O(N__14221),
            .I(N__14217));
    InMux I__1360 (
            .O(N__14220),
            .I(N__14214));
    LocalMux I__1359 (
            .O(N__14217),
            .I(N__14211));
    LocalMux I__1358 (
            .O(N__14214),
            .I(\POWERLED.count_clkZ0Z_14 ));
    Odrv4 I__1357 (
            .O(N__14211),
            .I(\POWERLED.count_clkZ0Z_14 ));
    CascadeMux I__1356 (
            .O(N__14206),
            .I(N__14202));
    InMux I__1355 (
            .O(N__14205),
            .I(N__14197));
    InMux I__1354 (
            .O(N__14202),
            .I(N__14197));
    LocalMux I__1353 (
            .O(N__14197),
            .I(N__14194));
    Odrv12 I__1352 (
            .O(N__14194),
            .I(\POWERLED.count_clk_1_14 ));
    InMux I__1351 (
            .O(N__14191),
            .I(\POWERLED.un1_count_clk_2_cry_13 ));
    InMux I__1350 (
            .O(N__14188),
            .I(N__14185));
    LocalMux I__1349 (
            .O(N__14185),
            .I(N__14181));
    InMux I__1348 (
            .O(N__14184),
            .I(N__14178));
    Odrv4 I__1347 (
            .O(N__14181),
            .I(\POWERLED.count_clkZ0Z_15 ));
    LocalMux I__1346 (
            .O(N__14178),
            .I(\POWERLED.count_clkZ0Z_15 ));
    InMux I__1345 (
            .O(N__14173),
            .I(\POWERLED.un1_count_clk_2_cry_14 ));
    CascadeMux I__1344 (
            .O(N__14170),
            .I(N__14167));
    InMux I__1343 (
            .O(N__14167),
            .I(N__14161));
    InMux I__1342 (
            .O(N__14166),
            .I(N__14161));
    LocalMux I__1341 (
            .O(N__14161),
            .I(N__14158));
    Span4Mux_s1_h I__1340 (
            .O(N__14158),
            .I(N__14155));
    Odrv4 I__1339 (
            .O(N__14155),
            .I(\POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ));
    InMux I__1338 (
            .O(N__14152),
            .I(N__14149));
    LocalMux I__1337 (
            .O(N__14149),
            .I(N__14146));
    Odrv4 I__1336 (
            .O(N__14146),
            .I(\POWERLED.count_clk_0_13 ));
    InMux I__1335 (
            .O(N__14143),
            .I(N__14140));
    LocalMux I__1334 (
            .O(N__14140),
            .I(N__14136));
    InMux I__1333 (
            .O(N__14139),
            .I(N__14133));
    Odrv12 I__1332 (
            .O(N__14136),
            .I(\POWERLED.count_clk_1_13 ));
    LocalMux I__1331 (
            .O(N__14133),
            .I(\POWERLED.count_clk_1_13 ));
    CascadeMux I__1330 (
            .O(N__14128),
            .I(N__14125));
    InMux I__1329 (
            .O(N__14125),
            .I(N__14122));
    LocalMux I__1328 (
            .O(N__14122),
            .I(N__14118));
    InMux I__1327 (
            .O(N__14121),
            .I(N__14115));
    Odrv4 I__1326 (
            .O(N__14118),
            .I(\POWERLED.count_clkZ0Z_13 ));
    LocalMux I__1325 (
            .O(N__14115),
            .I(\POWERLED.count_clkZ0Z_13 ));
    InMux I__1324 (
            .O(N__14110),
            .I(\POWERLED.un1_count_clk_2_cry_1 ));
    InMux I__1323 (
            .O(N__14107),
            .I(\POWERLED.un1_count_clk_2_cry_2 ));
    InMux I__1322 (
            .O(N__14104),
            .I(N__14098));
    InMux I__1321 (
            .O(N__14103),
            .I(N__14098));
    LocalMux I__1320 (
            .O(N__14098),
            .I(N__14095));
    Odrv4 I__1319 (
            .O(N__14095),
            .I(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ));
    InMux I__1318 (
            .O(N__14092),
            .I(\POWERLED.un1_count_clk_2_cry_3 ));
    InMux I__1317 (
            .O(N__14089),
            .I(\POWERLED.un1_count_clk_2_cry_4 ));
    InMux I__1316 (
            .O(N__14086),
            .I(\POWERLED.un1_count_clk_2_cry_5 ));
    InMux I__1315 (
            .O(N__14083),
            .I(\POWERLED.un1_count_clk_2_cry_6 ));
    InMux I__1314 (
            .O(N__14080),
            .I(\POWERLED.un1_count_clk_2_cry_7 ));
    InMux I__1313 (
            .O(N__14077),
            .I(bfn_1_12_0_));
    CascadeMux I__1312 (
            .O(N__14074),
            .I(N__14071));
    InMux I__1311 (
            .O(N__14071),
            .I(N__14068));
    LocalMux I__1310 (
            .O(N__14068),
            .I(\POWERLED.count_clk_0_10 ));
    CascadeMux I__1309 (
            .O(N__14065),
            .I(\POWERLED.un1_dutycycle_168_0_0_o2_1_4_cascade_ ));
    InMux I__1308 (
            .O(N__14062),
            .I(N__14059));
    LocalMux I__1307 (
            .O(N__14059),
            .I(\POWERLED.count_clk_0_14 ));
    CascadeMux I__1306 (
            .O(N__14056),
            .I(N__14053));
    InMux I__1305 (
            .O(N__14053),
            .I(N__14050));
    LocalMux I__1304 (
            .O(N__14050),
            .I(\POWERLED.count_clk_0_11 ));
    CascadeMux I__1303 (
            .O(N__14047),
            .I(N__14044));
    InMux I__1302 (
            .O(N__14044),
            .I(N__14041));
    LocalMux I__1301 (
            .O(N__14041),
            .I(\POWERLED.count_clk_0_12 ));
    InMux I__1300 (
            .O(N__14038),
            .I(\HDA_STRAP.un1_count_1_cry_13 ));
    InMux I__1299 (
            .O(N__14035),
            .I(\HDA_STRAP.un1_count_1_cry_14 ));
    InMux I__1298 (
            .O(N__14032),
            .I(N__14029));
    LocalMux I__1297 (
            .O(N__14029),
            .I(N__14024));
    InMux I__1296 (
            .O(N__14028),
            .I(N__14019));
    InMux I__1295 (
            .O(N__14027),
            .I(N__14019));
    Odrv12 I__1294 (
            .O(N__14024),
            .I(\HDA_STRAP.countZ0Z_16 ));
    LocalMux I__1293 (
            .O(N__14019),
            .I(\HDA_STRAP.countZ0Z_16 ));
    InMux I__1292 (
            .O(N__14014),
            .I(N__14011));
    LocalMux I__1291 (
            .O(N__14011),
            .I(N__14008));
    Odrv4 I__1290 (
            .O(N__14008),
            .I(\HDA_STRAP.un1_count_1_cry_15_THRU_CO ));
    InMux I__1289 (
            .O(N__14005),
            .I(bfn_1_8_0_));
    InMux I__1288 (
            .O(N__14002),
            .I(\HDA_STRAP.un1_count_1_cry_16 ));
    InMux I__1287 (
            .O(N__13999),
            .I(N__13995));
    InMux I__1286 (
            .O(N__13998),
            .I(N__13992));
    LocalMux I__1285 (
            .O(N__13995),
            .I(N__13989));
    LocalMux I__1284 (
            .O(N__13992),
            .I(\HDA_STRAP.countZ0Z_17 ));
    Odrv4 I__1283 (
            .O(N__13989),
            .I(\HDA_STRAP.countZ0Z_17 ));
    CascadeMux I__1282 (
            .O(N__13984),
            .I(N__13981));
    InMux I__1281 (
            .O(N__13981),
            .I(N__13978));
    LocalMux I__1280 (
            .O(N__13978),
            .I(\POWERLED.count_clk_0_4 ));
    InMux I__1279 (
            .O(N__13975),
            .I(N__13972));
    LocalMux I__1278 (
            .O(N__13972),
            .I(\POWERLED.count_clk_0_15 ));
    InMux I__1277 (
            .O(N__13969),
            .I(\HDA_STRAP.un1_count_1_cry_5 ));
    InMux I__1276 (
            .O(N__13966),
            .I(\HDA_STRAP.un1_count_1_cry_6 ));
    InMux I__1275 (
            .O(N__13963),
            .I(bfn_1_7_0_));
    InMux I__1274 (
            .O(N__13960),
            .I(\HDA_STRAP.un1_count_1_cry_8 ));
    InMux I__1273 (
            .O(N__13957),
            .I(N__13954));
    LocalMux I__1272 (
            .O(N__13954),
            .I(N__13949));
    InMux I__1271 (
            .O(N__13953),
            .I(N__13944));
    InMux I__1270 (
            .O(N__13952),
            .I(N__13944));
    Odrv4 I__1269 (
            .O(N__13949),
            .I(\HDA_STRAP.countZ0Z_10 ));
    LocalMux I__1268 (
            .O(N__13944),
            .I(\HDA_STRAP.countZ0Z_10 ));
    InMux I__1267 (
            .O(N__13939),
            .I(N__13936));
    LocalMux I__1266 (
            .O(N__13936),
            .I(N__13933));
    Odrv4 I__1265 (
            .O(N__13933),
            .I(\HDA_STRAP.un1_count_1_cry_9_THRU_CO ));
    InMux I__1264 (
            .O(N__13930),
            .I(\HDA_STRAP.un1_count_1_cry_9 ));
    InMux I__1263 (
            .O(N__13927),
            .I(N__13924));
    LocalMux I__1262 (
            .O(N__13924),
            .I(N__13919));
    InMux I__1261 (
            .O(N__13923),
            .I(N__13914));
    InMux I__1260 (
            .O(N__13922),
            .I(N__13914));
    Odrv4 I__1259 (
            .O(N__13919),
            .I(\HDA_STRAP.countZ0Z_11 ));
    LocalMux I__1258 (
            .O(N__13914),
            .I(\HDA_STRAP.countZ0Z_11 ));
    InMux I__1257 (
            .O(N__13909),
            .I(N__13906));
    LocalMux I__1256 (
            .O(N__13906),
            .I(N__13903));
    Odrv4 I__1255 (
            .O(N__13903),
            .I(\HDA_STRAP.un1_count_1_cry_10_THRU_CO ));
    InMux I__1254 (
            .O(N__13900),
            .I(\HDA_STRAP.un1_count_1_cry_10 ));
    InMux I__1253 (
            .O(N__13897),
            .I(\HDA_STRAP.un1_count_1_cry_11 ));
    InMux I__1252 (
            .O(N__13894),
            .I(\HDA_STRAP.un1_count_1_cry_12 ));
    CascadeMux I__1251 (
            .O(N__13891),
            .I(\HDA_STRAP.un4_count_10_cascade_ ));
    InMux I__1250 (
            .O(N__13888),
            .I(N__13885));
    LocalMux I__1249 (
            .O(N__13885),
            .I(\HDA_STRAP.un4_count_13 ));
    CascadeMux I__1248 (
            .O(N__13882),
            .I(\HDA_STRAP.un4_count_cascade_ ));
    CascadeMux I__1247 (
            .O(N__13879),
            .I(N__13875));
    InMux I__1246 (
            .O(N__13878),
            .I(N__13871));
    InMux I__1245 (
            .O(N__13875),
            .I(N__13868));
    InMux I__1244 (
            .O(N__13874),
            .I(N__13865));
    LocalMux I__1243 (
            .O(N__13871),
            .I(\HDA_STRAP.countZ0Z_0 ));
    LocalMux I__1242 (
            .O(N__13868),
            .I(\HDA_STRAP.countZ0Z_0 ));
    LocalMux I__1241 (
            .O(N__13865),
            .I(\HDA_STRAP.countZ0Z_0 ));
    InMux I__1240 (
            .O(N__13858),
            .I(N__13854));
    InMux I__1239 (
            .O(N__13857),
            .I(N__13851));
    LocalMux I__1238 (
            .O(N__13854),
            .I(\HDA_STRAP.countZ0Z_1 ));
    LocalMux I__1237 (
            .O(N__13851),
            .I(\HDA_STRAP.countZ0Z_1 ));
    InMux I__1236 (
            .O(N__13846),
            .I(\HDA_STRAP.un1_count_1_cry_0 ));
    InMux I__1235 (
            .O(N__13843),
            .I(N__13839));
    InMux I__1234 (
            .O(N__13842),
            .I(N__13836));
    LocalMux I__1233 (
            .O(N__13839),
            .I(\HDA_STRAP.countZ0Z_2 ));
    LocalMux I__1232 (
            .O(N__13836),
            .I(\HDA_STRAP.countZ0Z_2 ));
    InMux I__1231 (
            .O(N__13831),
            .I(\HDA_STRAP.un1_count_1_cry_1 ));
    CascadeMux I__1230 (
            .O(N__13828),
            .I(N__13825));
    InMux I__1229 (
            .O(N__13825),
            .I(N__13821));
    InMux I__1228 (
            .O(N__13824),
            .I(N__13818));
    LocalMux I__1227 (
            .O(N__13821),
            .I(\HDA_STRAP.countZ0Z_3 ));
    LocalMux I__1226 (
            .O(N__13818),
            .I(\HDA_STRAP.countZ0Z_3 ));
    InMux I__1225 (
            .O(N__13813),
            .I(\HDA_STRAP.un1_count_1_cry_2 ));
    InMux I__1224 (
            .O(N__13810),
            .I(N__13806));
    InMux I__1223 (
            .O(N__13809),
            .I(N__13803));
    LocalMux I__1222 (
            .O(N__13806),
            .I(\HDA_STRAP.countZ0Z_4 ));
    LocalMux I__1221 (
            .O(N__13803),
            .I(\HDA_STRAP.countZ0Z_4 ));
    InMux I__1220 (
            .O(N__13798),
            .I(\HDA_STRAP.un1_count_1_cry_3 ));
    InMux I__1219 (
            .O(N__13795),
            .I(N__13791));
    InMux I__1218 (
            .O(N__13794),
            .I(N__13788));
    LocalMux I__1217 (
            .O(N__13791),
            .I(\HDA_STRAP.countZ0Z_5 ));
    LocalMux I__1216 (
            .O(N__13788),
            .I(\HDA_STRAP.countZ0Z_5 ));
    InMux I__1215 (
            .O(N__13783),
            .I(\HDA_STRAP.un1_count_1_cry_4 ));
    InMux I__1214 (
            .O(N__13780),
            .I(N__13774));
    InMux I__1213 (
            .O(N__13779),
            .I(N__13774));
    LocalMux I__1212 (
            .O(N__13774),
            .I(N__13771));
    Odrv12 I__1211 (
            .O(N__13771),
            .I(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ));
    CascadeMux I__1210 (
            .O(N__13768),
            .I(\PCH_PWRGD.countZ0Z_3_cascade_ ));
    InMux I__1209 (
            .O(N__13765),
            .I(N__13762));
    LocalMux I__1208 (
            .O(N__13762),
            .I(\PCH_PWRGD.count_0_3 ));
    CascadeMux I__1207 (
            .O(N__13759),
            .I(\PCH_PWRGD.count_rst_10_cascade_ ));
    CascadeMux I__1206 (
            .O(N__13756),
            .I(\PCH_PWRGD.countZ0Z_4_cascade_ ));
    InMux I__1205 (
            .O(N__13753),
            .I(N__13747));
    InMux I__1204 (
            .O(N__13752),
            .I(N__13747));
    LocalMux I__1203 (
            .O(N__13747),
            .I(N__13744));
    Odrv4 I__1202 (
            .O(N__13744),
            .I(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ));
    InMux I__1201 (
            .O(N__13741),
            .I(N__13738));
    LocalMux I__1200 (
            .O(N__13738),
            .I(\PCH_PWRGD.count_0_4 ));
    CascadeMux I__1199 (
            .O(N__13735),
            .I(\HDA_STRAP.un4_count_9_cascade_ ));
    InMux I__1198 (
            .O(N__13732),
            .I(\PCH_PWRGD.un2_count_1_cry_11 ));
    InMux I__1197 (
            .O(N__13729),
            .I(\PCH_PWRGD.un2_count_1_cry_12 ));
    InMux I__1196 (
            .O(N__13726),
            .I(\PCH_PWRGD.un2_count_1_cry_13 ));
    InMux I__1195 (
            .O(N__13723),
            .I(\PCH_PWRGD.un2_count_1_cry_14 ));
    InMux I__1194 (
            .O(N__13720),
            .I(N__13717));
    LocalMux I__1193 (
            .O(N__13717),
            .I(\PCH_PWRGD.un2_count_1_axb_14 ));
    InMux I__1192 (
            .O(N__13714),
            .I(N__13708));
    InMux I__1191 (
            .O(N__13713),
            .I(N__13708));
    LocalMux I__1190 (
            .O(N__13708),
            .I(\PCH_PWRGD.un2_count_1_cry_12_c_RNIA8PZ0Z7 ));
    CascadeMux I__1189 (
            .O(N__13705),
            .I(N__13702));
    InMux I__1188 (
            .O(N__13702),
            .I(N__13699));
    LocalMux I__1187 (
            .O(N__13699),
            .I(\PCH_PWRGD.count_0_13 ));
    CascadeMux I__1186 (
            .O(N__13696),
            .I(\PCH_PWRGD.count_rst_11_cascade_ ));
    InMux I__1185 (
            .O(N__13693),
            .I(\PCH_PWRGD.un2_count_1_cry_2 ));
    InMux I__1184 (
            .O(N__13690),
            .I(\PCH_PWRGD.un2_count_1_cry_3 ));
    InMux I__1183 (
            .O(N__13687),
            .I(\PCH_PWRGD.un2_count_1_cry_4 ));
    InMux I__1182 (
            .O(N__13684),
            .I(\PCH_PWRGD.un2_count_1_cry_5 ));
    CascadeMux I__1181 (
            .O(N__13681),
            .I(N__13677));
    CascadeMux I__1180 (
            .O(N__13680),
            .I(N__13674));
    InMux I__1179 (
            .O(N__13677),
            .I(N__13668));
    InMux I__1178 (
            .O(N__13674),
            .I(N__13668));
    InMux I__1177 (
            .O(N__13673),
            .I(N__13665));
    LocalMux I__1176 (
            .O(N__13668),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    LocalMux I__1175 (
            .O(N__13665),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    InMux I__1174 (
            .O(N__13660),
            .I(N__13654));
    InMux I__1173 (
            .O(N__13659),
            .I(N__13654));
    LocalMux I__1172 (
            .O(N__13654),
            .I(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ));
    InMux I__1171 (
            .O(N__13651),
            .I(\PCH_PWRGD.un2_count_1_cry_6 ));
    CascadeMux I__1170 (
            .O(N__13648),
            .I(N__13645));
    InMux I__1169 (
            .O(N__13645),
            .I(N__13641));
    InMux I__1168 (
            .O(N__13644),
            .I(N__13638));
    LocalMux I__1167 (
            .O(N__13641),
            .I(\PCH_PWRGD.un2_count_1_axb_8 ));
    LocalMux I__1166 (
            .O(N__13638),
            .I(\PCH_PWRGD.un2_count_1_axb_8 ));
    InMux I__1165 (
            .O(N__13633),
            .I(N__13627));
    InMux I__1164 (
            .O(N__13632),
            .I(N__13627));
    LocalMux I__1163 (
            .O(N__13627),
            .I(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ));
    InMux I__1162 (
            .O(N__13624),
            .I(\PCH_PWRGD.un2_count_1_cry_7 ));
    InMux I__1161 (
            .O(N__13621),
            .I(bfn_1_3_0_));
    InMux I__1160 (
            .O(N__13618),
            .I(\PCH_PWRGD.un2_count_1_cry_9 ));
    InMux I__1159 (
            .O(N__13615),
            .I(\PCH_PWRGD.un2_count_1_cry_10 ));
    InMux I__1158 (
            .O(N__13612),
            .I(N__13609));
    LocalMux I__1157 (
            .O(N__13609),
            .I(\PCH_PWRGD.count_rst_6 ));
    CascadeMux I__1156 (
            .O(N__13606),
            .I(\PCH_PWRGD.count_rst_6_cascade_ ));
    CascadeMux I__1155 (
            .O(N__13603),
            .I(\PCH_PWRGD.un2_count_1_axb_8_cascade_ ));
    InMux I__1154 (
            .O(N__13600),
            .I(N__13594));
    InMux I__1153 (
            .O(N__13599),
            .I(N__13594));
    LocalMux I__1152 (
            .O(N__13594),
            .I(\PCH_PWRGD.count_0_8 ));
    CascadeMux I__1151 (
            .O(N__13591),
            .I(\PCH_PWRGD.count_rst_7_cascade_ ));
    CascadeMux I__1150 (
            .O(N__13588),
            .I(\PCH_PWRGD.countZ0Z_7_cascade_ ));
    InMux I__1149 (
            .O(N__13585),
            .I(N__13582));
    LocalMux I__1148 (
            .O(N__13582),
            .I(\PCH_PWRGD.count_0_7 ));
    InMux I__1147 (
            .O(N__13579),
            .I(\PCH_PWRGD.un2_count_1_cry_1 ));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_6_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_12_0_));
    defparam IN_MUX_bfv_6_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_13_0_ (
            .carryinitin(\POWERLED.un3_count_off_1_cry_8 ),
            .carryinitout(bfn_6_13_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_1_0_));
    defparam IN_MUX_bfv_9_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_1_0_));
    defparam IN_MUX_bfv_9_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_2_0_));
    defparam IN_MUX_bfv_11_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_2_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_9_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_3_0_));
    defparam IN_MUX_bfv_9_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_4_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_5_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_5_0_));
    defparam IN_MUX_bfv_4_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_5_0_));
    defparam IN_MUX_bfv_4_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_6_0_));
    defparam IN_MUX_bfv_5_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_6_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_7_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_4_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_5_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_2_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(\POWERLED.un1_count_cry_8 ),
            .carryinitout(bfn_5_3_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_2_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(\PCH_PWRGD.un2_count_1_cry_8 ),
            .carryinitout(bfn_1_3_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(\HDA_STRAP.un1_count_1_cry_7 ),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(\HDA_STRAP.un1_count_1_cry_15 ),
            .carryinitout(bfn_1_8_0_));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(COUNTER_un4_counter_7),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\COUNTER.counter_1_cry_8 ),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\COUNTER.counter_1_cry_16 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\COUNTER.counter_1_cry_24 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_7 ),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_7 ),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_6_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_8_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_94_cry_7_cZ0 ),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_7_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_5_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_7_cZ0 ),
            .carryinitout(bfn_7_6_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_15 ),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_4_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_15_0_ (
            .carryinitin(\DSW_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_4_15_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(\DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_4_16_0_));
    ICE_GB N_587_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__28176),
            .GLOBALBUFFEROUTPUT(N_587_g));
    ICE_GB N_42_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__20491),
            .GLOBALBUFFEROUTPUT(N_42_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIQOP84_0_8_LC_1_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQOP84_0_8_LC_1_1_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQOP84_0_8_LC_1_1_0 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \PCH_PWRGD.count_RNIQOP84_0_8_LC_1_1_0  (
            .in0(N__21156),
            .in1(N__13612),
            .in2(N__13680),
            .in3(N__13600),
            .lcout(\PCH_PWRGD.count_1_i_a2_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIPICU1_LC_1_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIPICU1_LC_1_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIPICU1_LC_1_1_1 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_c_RNIPICU1_LC_1_1_1  (
            .in0(N__14996),
            .in1(N__13632),
            .in2(N__13648),
            .in3(N__20967),
            .lcout(\PCH_PWRGD.count_rst_6 ),
            .ltout(\PCH_PWRGD.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIQOP84_8_LC_1_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQOP84_8_LC_1_1_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQOP84_8_LC_1_1_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNIQOP84_8_LC_1_1_2  (
            .in0(N__21145),
            .in1(_gnd_net_),
            .in2(N__13606),
            .in3(N__13599),
            .lcout(\PCH_PWRGD.un2_count_1_axb_8 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_8_LC_1_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_8_LC_1_1_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_8_LC_1_1_3 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \PCH_PWRGD.count_8_LC_1_1_3  (
            .in0(N__14998),
            .in1(N__20970),
            .in2(N__13603),
            .in3(N__13633),
            .lcout(\PCH_PWRGD.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32817),
            .ce(N__21155),
            .sr(N__21006));
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIOGBU1_LC_1_1_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIOGBU1_LC_1_1_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIOGBU1_LC_1_1_4 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_c_RNIOGBU1_LC_1_1_4  (
            .in0(N__20966),
            .in1(N__13659),
            .in2(N__13681),
            .in3(N__14995),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIOLO84_7_LC_1_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIOLO84_7_LC_1_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIOLO84_7_LC_1_1_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.count_RNIOLO84_7_LC_1_1_5  (
            .in0(_gnd_net_),
            .in1(N__13585),
            .in2(N__13591),
            .in3(N__21144),
            .lcout(\PCH_PWRGD.countZ0Z_7 ),
            .ltout(\PCH_PWRGD.countZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_7_LC_1_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_7_LC_1_1_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_7_LC_1_1_6 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.count_7_LC_1_1_6  (
            .in0(N__20968),
            .in1(N__13660),
            .in2(N__13588),
            .in3(N__14999),
            .lcout(\PCH_PWRGD.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32817),
            .ce(N__21155),
            .sr(N__21006));
    defparam \PCH_PWRGD.count_5_LC_1_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_5_LC_1_1_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_5_LC_1_1_7 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \PCH_PWRGD.count_5_LC_1_1_7  (
            .in0(N__14997),
            .in1(N__20969),
            .in2(N__14653),
            .in3(N__14803),
            .lcout(\PCH_PWRGD.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32817),
            .ce(N__21155),
            .sr(N__21006));
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_2_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_2_0  (
            .in0(_gnd_net_),
            .in1(N__14460),
            .in2(N__14437),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_2_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNIJ66U1_LC_1_2_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNIJ66U1_LC_1_2_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNIJ66U1_LC_1_2_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_1_c_RNIJ66U1_LC_1_2_1  (
            .in0(N__20948),
            .in1(N__14845),
            .in2(_gnd_net_),
            .in3(N__13579),
            .lcout(\PCH_PWRGD.count_rst_12 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_1 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_2_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_2_2  (
            .in0(_gnd_net_),
            .in1(N__14775),
            .in2(_gnd_net_),
            .in3(N__13693),
            .lcout(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_2 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_2_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_2_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_2_3  (
            .in0(_gnd_net_),
            .in1(N__14748),
            .in2(_gnd_net_),
            .in3(N__13690),
            .lcout(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_3 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_2_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_2_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_2_4  (
            .in0(_gnd_net_),
            .in1(N__14797),
            .in2(_gnd_net_),
            .in3(N__13687),
            .lcout(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_4 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNINEAU1_LC_1_2_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNINEAU1_LC_1_2_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNINEAU1_LC_1_2_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_5_c_RNINEAU1_LC_1_2_5  (
            .in0(N__20949),
            .in1(N__14829),
            .in2(_gnd_net_),
            .in3(N__13684),
            .lcout(\PCH_PWRGD.count_rst_8 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_5 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_2_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_2_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_2_6  (
            .in0(_gnd_net_),
            .in1(N__13673),
            .in2(_gnd_net_),
            .in3(N__13651),
            .lcout(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_6 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_2_7 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_2_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_2_7  (
            .in0(_gnd_net_),
            .in1(N__13644),
            .in2(_gnd_net_),
            .in3(N__13624),
            .lcout(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_7 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_3_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_3_0  (
            .in0(_gnd_net_),
            .in1(N__14619),
            .in2(_gnd_net_),
            .in3(N__13621),
            .lcout(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIRMEU1_LC_1_3_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIRMEU1_LC_1_3_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIRMEU1_LC_1_3_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_9_c_RNIRMEU1_LC_1_3_1  (
            .in0(N__20984),
            .in1(N__14851),
            .in2(_gnd_net_),
            .in3(N__13618),
            .lcout(\PCH_PWRGD.count_rst_4 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_9 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_3_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_3_2  (
            .in0(_gnd_net_),
            .in1(N__14688),
            .in2(_gnd_net_),
            .in3(N__13615),
            .lcout(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_10 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNI402P1_LC_1_3_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNI402P1_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNI402P1_LC_1_3_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_11_c_RNI402P1_LC_1_3_3  (
            .in0(N__20985),
            .in1(N__14814),
            .in2(_gnd_net_),
            .in3(N__13732),
            .lcout(\PCH_PWRGD.count_rst_2 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_11 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8P7_LC_1_3_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8P7_LC_1_3_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8P7_LC_1_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8P7_LC_1_3_4  (
            .in0(_gnd_net_),
            .in1(N__14577),
            .in2(_gnd_net_),
            .in3(N__13729),
            .lcout(\PCH_PWRGD.un2_count_1_cry_12_c_RNIA8PZ0Z7 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_12 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIKP0C4_LC_1_3_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIKP0C4_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIKP0C4_LC_1_3_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_13_c_RNIKP0C4_LC_1_3_5  (
            .in0(N__20986),
            .in1(N__13720),
            .in2(_gnd_net_),
            .in3(N__13726),
            .lcout(\PCH_PWRGD.count_rst_0 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_13 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNI765P1_LC_1_3_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNI765P1_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNI765P1_LC_1_3_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_14_c_RNI765P1_LC_1_3_6  (
            .in0(N__16593),
            .in1(N__20987),
            .in2(_gnd_net_),
            .in3(N__13723),
            .lcout(\PCH_PWRGD.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIELSI2_14_LC_1_3_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIELSI2_14_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIELSI2_14_LC_1_3_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \PCH_PWRGD.count_RNIELSI2_14_LC_1_3_7  (
            .in0(N__14499),
            .in1(N__21102),
            .in2(_gnd_net_),
            .in3(N__14513),
            .lcout(\PCH_PWRGD.un2_count_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIIMVB4_13_LC_1_4_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIIMVB4_13_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIIMVB4_13_LC_1_4_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \PCH_PWRGD.count_RNIIMVB4_13_LC_1_4_0  (
            .in0(N__21100),
            .in1(N__20875),
            .in2(N__13705),
            .in3(N__13713),
            .lcout(\PCH_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_13_LC_1_4_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_13_LC_1_4_1 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_13_LC_1_4_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \PCH_PWRGD.count_13_LC_1_4_1  (
            .in0(N__13714),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20874),
            .lcout(\PCH_PWRGD.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32903),
            .ce(N__21101),
            .sr(N__20977));
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNIK87U1_LC_1_4_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNIK87U1_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNIK87U1_LC_1_4_2 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_c_RNIK87U1_LC_1_4_2  (
            .in0(N__13779),
            .in1(N__14771),
            .in2(N__20931),
            .in3(N__15008),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIG9K84_3_LC_1_4_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIG9K84_3_LC_1_4_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIG9K84_3_LC_1_4_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.count_RNIG9K84_3_LC_1_4_3  (
            .in0(_gnd_net_),
            .in1(N__13765),
            .in2(N__13696),
            .in3(N__21098),
            .lcout(\PCH_PWRGD.countZ0Z_3 ),
            .ltout(\PCH_PWRGD.countZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_3_LC_1_4_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_3_LC_1_4_4 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_3_LC_1_4_4 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.count_3_LC_1_4_4  (
            .in0(N__13780),
            .in1(N__20876),
            .in2(N__13768),
            .in3(N__15011),
            .lcout(\PCH_PWRGD.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32903),
            .ce(N__21101),
            .sr(N__20977));
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNILA8U1_LC_1_4_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNILA8U1_LC_1_4_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNILA8U1_LC_1_4_5 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_c_RNILA8U1_LC_1_4_5  (
            .in0(N__15009),
            .in1(N__13752),
            .in2(N__14749),
            .in3(N__20872),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIICL84_4_LC_1_4_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIICL84_4_LC_1_4_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIICL84_4_LC_1_4_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNIICL84_4_LC_1_4_6  (
            .in0(N__21099),
            .in1(_gnd_net_),
            .in2(N__13759),
            .in3(N__13741),
            .lcout(\PCH_PWRGD.countZ0Z_4 ),
            .ltout(\PCH_PWRGD.countZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_4_LC_1_4_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_4_LC_1_4_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_4_LC_1_4_7 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \PCH_PWRGD.count_4_LC_1_4_7  (
            .in0(N__15010),
            .in1(N__20873),
            .in2(N__13756),
            .in3(N__13753),
            .lcout(\PCH_PWRGD.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32903),
            .ce(N__21101),
            .sr(N__20977));
    defparam \HDA_STRAP.count_0_LC_1_5_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_0_LC_1_5_0 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_0_LC_1_5_0 .LUT_INIT=16'b0000011001100110;
    LogicCell40 \HDA_STRAP.count_0_LC_1_5_0  (
            .in0(N__13878),
            .in1(N__15395),
            .in2(N__15414),
            .in3(N__15300),
            .lcout(\HDA_STRAP.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32901),
            .ce(N__27388),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_16_LC_1_5_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_16_LC_1_5_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_16_LC_1_5_1 .LUT_INIT=16'b0000011001100110;
    LogicCell40 \HDA_STRAP.count_16_LC_1_5_1  (
            .in0(N__14028),
            .in1(N__14014),
            .in2(N__15309),
            .in3(N__15407),
            .lcout(\HDA_STRAP.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32901),
            .ce(N__27388),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_10_LC_1_5_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_10_LC_1_5_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_10_LC_1_5_2 .LUT_INIT=16'b0000011001100110;
    LogicCell40 \HDA_STRAP.count_10_LC_1_5_2  (
            .in0(N__13939),
            .in1(N__13953),
            .in2(N__15413),
            .in3(N__15301),
            .lcout(\HDA_STRAP.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32901),
            .ce(N__27388),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_1_5_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_1_5_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \HDA_STRAP.count_RNI4CB61_17_LC_1_5_3  (
            .in0(N__14027),
            .in1(N__13857),
            .in2(N__13879),
            .in3(N__13999),
            .lcout(),
            .ltout(\HDA_STRAP.un4_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIH7IR1_10_LC_1_5_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIH7IR1_10_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIH7IR1_10_LC_1_5_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \HDA_STRAP.count_RNIH7IR1_10_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(N__13922),
            .in2(N__13735),
            .in3(N__13952),
            .lcout(\HDA_STRAP.un4_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI2L821_2_LC_1_5_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI2L821_2_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI2L821_2_LC_1_5_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \HDA_STRAP.count_RNI2L821_2_LC_1_5_5  (
            .in0(N__13794),
            .in1(N__13843),
            .in2(N__13828),
            .in3(N__13809),
            .lcout(),
            .ltout(\HDA_STRAP.un4_count_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_1_5_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_1_5_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \HDA_STRAP.count_RNIB5IA5_2_LC_1_5_6  (
            .in0(N__15106),
            .in1(N__15070),
            .in2(N__13891),
            .in3(N__13888),
            .lcout(\HDA_STRAP.un4_count ),
            .ltout(\HDA_STRAP.un4_count_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_11_LC_1_5_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_11_LC_1_5_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_11_LC_1_5_7 .LUT_INIT=16'b0001010100101010;
    LogicCell40 \HDA_STRAP.count_11_LC_1_5_7  (
            .in0(N__13923),
            .in1(N__15400),
            .in2(N__13882),
            .in3(N__13909),
            .lcout(\HDA_STRAP.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32901),
            .ce(N__27388),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_0_c_LC_1_6_0 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_0_c_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_0_c_LC_1_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_0_c_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__13874),
            .in2(N__15412),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_1_LC_1_6_1 .C_ON=1'b1;
    defparam \HDA_STRAP.count_1_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_1_LC_1_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_1_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__13858),
            .in2(_gnd_net_),
            .in3(N__13846),
            .lcout(\HDA_STRAP.countZ0Z_1 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_0 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_1 ),
            .clk(N__32964),
            .ce(N__27394),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_2_LC_1_6_2 .C_ON=1'b1;
    defparam \HDA_STRAP.count_2_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_2_LC_1_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_2_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(N__13842),
            .in2(_gnd_net_),
            .in3(N__13831),
            .lcout(\HDA_STRAP.countZ0Z_2 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_1 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_2 ),
            .clk(N__32964),
            .ce(N__27394),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_3_LC_1_6_3 .C_ON=1'b1;
    defparam \HDA_STRAP.count_3_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_3_LC_1_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_3_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(N__13824),
            .in2(_gnd_net_),
            .in3(N__13813),
            .lcout(\HDA_STRAP.countZ0Z_3 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_2 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_3 ),
            .clk(N__32964),
            .ce(N__27394),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_4_LC_1_6_4 .C_ON=1'b1;
    defparam \HDA_STRAP.count_4_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_4_LC_1_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_4_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(N__13810),
            .in2(_gnd_net_),
            .in3(N__13798),
            .lcout(\HDA_STRAP.countZ0Z_4 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_3 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_4 ),
            .clk(N__32964),
            .ce(N__27394),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_5_LC_1_6_5 .C_ON=1'b1;
    defparam \HDA_STRAP.count_5_LC_1_6_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_5_LC_1_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_5_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(N__13795),
            .in2(_gnd_net_),
            .in3(N__13783),
            .lcout(\HDA_STRAP.countZ0Z_5 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_4 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_5 ),
            .clk(N__32964),
            .ce(N__27394),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_1_6_6 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_1_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(N__15050),
            .in2(_gnd_net_),
            .in3(N__13969),
            .lcout(\HDA_STRAP.un1_count_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_5 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_7_LC_1_6_7 .C_ON=1'b1;
    defparam \HDA_STRAP.count_7_LC_1_6_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_7_LC_1_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_7_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(N__15118),
            .in2(_gnd_net_),
            .in3(N__13966),
            .lcout(\HDA_STRAP.countZ0Z_7 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_6 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_7 ),
            .clk(N__32964),
            .ce(N__27394),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_1_7_0 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_1_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__15430),
            .in2(_gnd_net_),
            .in3(N__13963),
            .lcout(\HDA_STRAP.un1_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_9_LC_1_7_1 .C_ON=1'b1;
    defparam \HDA_STRAP.count_9_LC_1_7_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_9_LC_1_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_9_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(N__15145),
            .in2(_gnd_net_),
            .in3(N__13960),
            .lcout(\HDA_STRAP.countZ0Z_9 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_8 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_9 ),
            .clk(N__32902),
            .ce(N__27387),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_1_7_2 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_1_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_1_7_2  (
            .in0(_gnd_net_),
            .in1(N__13957),
            .in2(_gnd_net_),
            .in3(N__13930),
            .lcout(\HDA_STRAP.un1_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_9 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_1_7_3 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_1_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_1_7_3  (
            .in0(_gnd_net_),
            .in1(N__13927),
            .in2(_gnd_net_),
            .in3(N__13900),
            .lcout(\HDA_STRAP.un1_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_10 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_12_LC_1_7_4 .C_ON=1'b1;
    defparam \HDA_STRAP.count_12_LC_1_7_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_12_LC_1_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_12_LC_1_7_4  (
            .in0(_gnd_net_),
            .in1(N__15132),
            .in2(_gnd_net_),
            .in3(N__13897),
            .lcout(\HDA_STRAP.countZ0Z_12 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_11 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_12 ),
            .clk(N__32902),
            .ce(N__27387),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_13_LC_1_7_5 .C_ON=1'b1;
    defparam \HDA_STRAP.count_13_LC_1_7_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_13_LC_1_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_13_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(N__15157),
            .in2(_gnd_net_),
            .in3(N__13894),
            .lcout(\HDA_STRAP.countZ0Z_13 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_12 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_13 ),
            .clk(N__32902),
            .ce(N__27387),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_14_LC_1_7_6 .C_ON=1'b1;
    defparam \HDA_STRAP.count_14_LC_1_7_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_14_LC_1_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_14_LC_1_7_6  (
            .in0(_gnd_net_),
            .in1(N__15094),
            .in2(_gnd_net_),
            .in3(N__14038),
            .lcout(\HDA_STRAP.countZ0Z_14 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_13 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_14 ),
            .clk(N__32902),
            .ce(N__27387),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_15_LC_1_7_7 .C_ON=1'b1;
    defparam \HDA_STRAP.count_15_LC_1_7_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_15_LC_1_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_15_LC_1_7_7  (
            .in0(_gnd_net_),
            .in1(N__15082),
            .in2(_gnd_net_),
            .in3(N__14035),
            .lcout(\HDA_STRAP.countZ0Z_15 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_14 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_15 ),
            .clk(N__32902),
            .ce(N__27387),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_1_8_0 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_1_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(N__14032),
            .in2(_gnd_net_),
            .in3(N__14005),
            .lcout(\HDA_STRAP.un1_count_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_8_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_17_LC_1_8_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_17_LC_1_8_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_17_LC_1_8_1 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \HDA_STRAP.count_17_LC_1_8_1  (
            .in0(N__15408),
            .in1(N__13998),
            .in2(N__15310),
            .in3(N__14002),
            .lcout(\HDA_STRAP.countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32979),
            .ce(N__27390),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI399J_4_LC_1_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI399J_4_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI399J_4_LC_1_9_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNI399J_4_LC_1_9_0  (
            .in0(N__33942),
            .in1(N__14103),
            .in2(N__13984),
            .in3(N__16930),
            .lcout(\POWERLED.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_4_LC_1_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_4_LC_1_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_4_LC_1_9_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_4_LC_1_9_1  (
            .in0(N__14104),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32990),
            .ce(N__16934),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_13_LC_1_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_13_LC_1_9_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_13_LC_1_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_13_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14143),
            .lcout(\POWERLED.count_clk_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32990),
            .ce(N__16934),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI7JKB_15_LC_1_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI7JKB_15_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI7JKB_15_LC_1_9_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.count_clk_RNI7JKB_15_LC_1_9_4  (
            .in0(N__33944),
            .in1(N__13975),
            .in2(N__14170),
            .in3(N__16932),
            .lcout(\POWERLED.count_clkZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_15_LC_1_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_15_LC_1_9_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_15_LC_1_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_15_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14166),
            .lcout(\POWERLED.count_clk_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32990),
            .ce(N__16934),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIM1VB_10_LC_1_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIM1VB_10_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIM1VB_10_LC_1_9_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNIM1VB_10_LC_1_9_6  (
            .in0(N__33943),
            .in1(N__14298),
            .in2(N__14074),
            .in3(N__16931),
            .lcout(\POWERLED.count_clkZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_10_LC_1_9_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_10_LC_1_9_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_10_LC_1_9_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_10_LC_1_9_7  (
            .in0(N__14299),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32990),
            .ce(N__16934),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI5GJB_14_LC_1_10_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI5GJB_14_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI5GJB_14_LC_1_10_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.count_clk_RNI5GJB_14_LC_1_10_0  (
            .in0(N__16924),
            .in1(N__14062),
            .in2(N__14206),
            .in3(N__33941),
            .lcout(\POWERLED.count_clkZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_15_LC_1_10_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_15_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_15_LC_1_10_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNI_15_LC_1_10_1  (
            .in0(N__14313),
            .in1(N__14184),
            .in2(N__14128),
            .in3(N__15826),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_168_0_0_o2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_11_LC_1_10_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_11_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_11_LC_1_10_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNI_11_LC_1_10_2  (
            .in0(N__14283),
            .in1(N__14253),
            .in2(N__14065),
            .in3(N__14220),
            .lcout(\POWERLED.N_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIV6GB_11_LC_1_10_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIV6GB_11_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIV6GB_11_LC_1_10_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNIV6GB_11_LC_1_10_3  (
            .in0(N__33939),
            .in1(N__14268),
            .in2(N__14056),
            .in3(N__16922),
            .lcout(\POWERLED.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_14_LC_1_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_14_LC_1_10_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_14_LC_1_10_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_14_LC_1_10_4  (
            .in0(N__14205),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33018),
            .ce(N__16935),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI1AHB_12_LC_1_10_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI1AHB_12_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI1AHB_12_LC_1_10_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNI1AHB_12_LC_1_10_5  (
            .in0(N__33940),
            .in1(N__14238),
            .in2(N__14047),
            .in3(N__16923),
            .lcout(\POWERLED.count_clkZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_11_LC_1_10_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_11_LC_1_10_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_11_LC_1_10_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_11_LC_1_10_6  (
            .in0(N__14269),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33018),
            .ce(N__16935),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_12_LC_1_10_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_12_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_12_LC_1_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_12_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14239),
            .lcout(\POWERLED.count_clk_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33018),
            .ce(N__16935),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_1_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__15823),
            .in2(N__15790),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_1_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_1_11_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_1_11_1  (
            .in0(N__15869),
            .in1(N__15663),
            .in2(_gnd_net_),
            .in3(N__14110),
            .lcout(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_1 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_1_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_1_11_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_1_11_2  (
            .in0(N__15873),
            .in1(N__15508),
            .in2(_gnd_net_),
            .in3(N__14107),
            .lcout(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_2 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_1_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_1_11_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_1_11_3  (
            .in0(N__15870),
            .in1(_gnd_net_),
            .in2(N__15484),
            .in3(N__14092),
            .lcout(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_3 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_1_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_1_11_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_1_11_4  (
            .in0(N__15874),
            .in1(N__15579),
            .in2(_gnd_net_),
            .in3(N__14089),
            .lcout(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_4 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_1_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_1_11_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_1_11_5  (
            .in0(N__15871),
            .in1(N__15738),
            .in2(_gnd_net_),
            .in3(N__14086),
            .lcout(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_5 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_1_11_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_1_11_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_1_11_6  (
            .in0(N__15875),
            .in1(N__16117),
            .in2(_gnd_net_),
            .in3(N__14083),
            .lcout(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_6 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_1_11_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_1_11_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_1_11_7  (
            .in0(N__15872),
            .in1(N__15699),
            .in2(_gnd_net_),
            .in3(N__14080),
            .lcout(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_7 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_1_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_1_12_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_1_12_0  (
            .in0(N__15901),
            .in1(N__15606),
            .in2(_gnd_net_),
            .in3(N__14077),
            .lcout(\POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_9_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_1_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_1_12_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_1_12_1  (
            .in0(N__15904),
            .in1(_gnd_net_),
            .in2(N__14317),
            .in3(N__14287),
            .lcout(\POWERLED.count_clk_1_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_9_cZ0 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_1_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_1_12_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_1_12_2  (
            .in0(N__15902),
            .in1(N__14284),
            .in2(_gnd_net_),
            .in3(N__14257),
            .lcout(\POWERLED.count_clk_1_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_10 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_1_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_1_12_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_1_12_3  (
            .in0(N__15905),
            .in1(N__14254),
            .in2(_gnd_net_),
            .in3(N__14227),
            .lcout(\POWERLED.count_clk_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_11 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_1_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_1_12_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_1_12_4  (
            .in0(N__15903),
            .in1(N__14121),
            .in2(_gnd_net_),
            .in3(N__14224),
            .lcout(\POWERLED.count_clk_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_12 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_1_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_1_12_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_1_12_5  (
            .in0(N__15906),
            .in1(N__14221),
            .in2(_gnd_net_),
            .in3(N__14191),
            .lcout(\POWERLED.count_clk_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_13 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_1_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_1_12_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_1_12_6  (
            .in0(N__14188),
            .in1(N__15907),
            .in2(_gnd_net_),
            .in3(N__14173),
            .lcout(\POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI3DIB_13_LC_1_12_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI3DIB_13_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI3DIB_13_LC_1_12_7 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \POWERLED.count_clk_RNI3DIB_13_LC_1_12_7  (
            .in0(N__14152),
            .in1(N__14139),
            .in2(N__33923),
            .in3(N__16920),
            .lcout(\POWERLED.count_clkZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_c_LC_1_13_0 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_c_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_c_LC_1_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.counter_1_cry_1_c_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__17380),
            .in2(N__18519),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\COUNTER.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_1_13_1 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_1_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__18592),
            .in2(_gnd_net_),
            .in3(N__14344),
            .lcout(\COUNTER.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_1 ),
            .carryout(\COUNTER.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_1_13_2 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_1_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__17041),
            .in2(_gnd_net_),
            .in3(N__14341),
            .lcout(\COUNTER.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_2 ),
            .carryout(\COUNTER.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_1_13_3 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_1_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__17308),
            .in2(_gnd_net_),
            .in3(N__14338),
            .lcout(\COUNTER.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_3 ),
            .carryout(\COUNTER.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_1_13_4 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_1_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__17359),
            .in2(_gnd_net_),
            .in3(N__14335),
            .lcout(\COUNTER.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_4 ),
            .carryout(\COUNTER.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_1_13_5 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_1_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__17278),
            .in2(_gnd_net_),
            .in3(N__14332),
            .lcout(\COUNTER.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_5 ),
            .carryout(\COUNTER.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_7_LC_1_13_6 .C_ON=1'b1;
    defparam \COUNTER.counter_7_LC_1_13_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_7_LC_1_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_7_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__17340),
            .in2(_gnd_net_),
            .in3(N__14329),
            .lcout(\COUNTER.counterZ0Z_7 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_6 ),
            .carryout(\COUNTER.counter_1_cry_7 ),
            .clk(N__33037),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_8_LC_1_13_7 .C_ON=1'b1;
    defparam \COUNTER.counter_8_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_8_LC_1_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_8_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__16060),
            .in2(_gnd_net_),
            .in3(N__14326),
            .lcout(\COUNTER.counterZ0Z_8 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_7 ),
            .carryout(\COUNTER.counter_1_cry_8 ),
            .clk(N__33037),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_9_LC_1_14_0 .C_ON=1'b1;
    defparam \COUNTER.counter_9_LC_1_14_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_9_LC_1_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_9_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__16021),
            .in2(_gnd_net_),
            .in3(N__14323),
            .lcout(\COUNTER.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\COUNTER.counter_1_cry_9 ),
            .clk(N__33044),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_10_LC_1_14_1 .C_ON=1'b1;
    defparam \COUNTER.counter_10_LC_1_14_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_10_LC_1_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_10_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__16035),
            .in2(_gnd_net_),
            .in3(N__14320),
            .lcout(\COUNTER.counterZ0Z_10 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_9 ),
            .carryout(\COUNTER.counter_1_cry_10 ),
            .clk(N__33044),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_11_LC_1_14_2 .C_ON=1'b1;
    defparam \COUNTER.counter_11_LC_1_14_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_11_LC_1_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_11_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__16048),
            .in2(_gnd_net_),
            .in3(N__14371),
            .lcout(\COUNTER.counterZ0Z_11 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_10 ),
            .carryout(\COUNTER.counter_1_cry_11 ),
            .clk(N__33044),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_12_LC_1_14_3 .C_ON=1'b1;
    defparam \COUNTER.counter_12_LC_1_14_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_12_LC_1_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_12_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__15970),
            .in2(_gnd_net_),
            .in3(N__14368),
            .lcout(\COUNTER.counterZ0Z_12 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_11 ),
            .carryout(\COUNTER.counter_1_cry_12 ),
            .clk(N__33044),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_13_LC_1_14_4 .C_ON=1'b1;
    defparam \COUNTER.counter_13_LC_1_14_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_13_LC_1_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_13_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__15997),
            .in2(_gnd_net_),
            .in3(N__14365),
            .lcout(\COUNTER.counterZ0Z_13 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_12 ),
            .carryout(\COUNTER.counter_1_cry_13 ),
            .clk(N__33044),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_14_LC_1_14_5 .C_ON=1'b1;
    defparam \COUNTER.counter_14_LC_1_14_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_14_LC_1_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_14_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__16009),
            .in2(_gnd_net_),
            .in3(N__14362),
            .lcout(\COUNTER.counterZ0Z_14 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_13 ),
            .carryout(\COUNTER.counter_1_cry_14 ),
            .clk(N__33044),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_15_LC_1_14_6 .C_ON=1'b1;
    defparam \COUNTER.counter_15_LC_1_14_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_15_LC_1_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_15_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__15984),
            .in2(_gnd_net_),
            .in3(N__14359),
            .lcout(\COUNTER.counterZ0Z_15 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_14 ),
            .carryout(\COUNTER.counter_1_cry_15 ),
            .clk(N__33044),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_16_LC_1_14_7 .C_ON=1'b1;
    defparam \COUNTER.counter_16_LC_1_14_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_16_LC_1_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_16_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__15919),
            .in2(_gnd_net_),
            .in3(N__14356),
            .lcout(\COUNTER.counterZ0Z_16 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_15 ),
            .carryout(\COUNTER.counter_1_cry_16 ),
            .clk(N__33044),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_17_LC_1_15_0 .C_ON=1'b1;
    defparam \COUNTER.counter_17_LC_1_15_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_17_LC_1_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_17_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__15946),
            .in2(_gnd_net_),
            .in3(N__14353),
            .lcout(\COUNTER.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\COUNTER.counter_1_cry_17 ),
            .clk(N__33022),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_18_LC_1_15_1 .C_ON=1'b1;
    defparam \COUNTER.counter_18_LC_1_15_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_18_LC_1_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_18_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__15958),
            .in2(_gnd_net_),
            .in3(N__14350),
            .lcout(\COUNTER.counterZ0Z_18 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_17 ),
            .carryout(\COUNTER.counter_1_cry_18 ),
            .clk(N__33022),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_19_LC_1_15_2 .C_ON=1'b1;
    defparam \COUNTER.counter_19_LC_1_15_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_19_LC_1_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_19_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__15933),
            .in2(_gnd_net_),
            .in3(N__14347),
            .lcout(\COUNTER.counterZ0Z_19 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_18 ),
            .carryout(\COUNTER.counter_1_cry_19 ),
            .clk(N__33022),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_20_LC_1_15_3 .C_ON=1'b1;
    defparam \COUNTER.counter_20_LC_1_15_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_20_LC_1_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_20_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__16372),
            .in2(_gnd_net_),
            .in3(N__14401),
            .lcout(\COUNTER.counterZ0Z_20 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_19 ),
            .carryout(\COUNTER.counter_1_cry_20 ),
            .clk(N__33022),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_21_LC_1_15_4 .C_ON=1'b1;
    defparam \COUNTER.counter_21_LC_1_15_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_21_LC_1_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_21_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__16345),
            .in2(_gnd_net_),
            .in3(N__14398),
            .lcout(\COUNTER.counterZ0Z_21 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_20 ),
            .carryout(\COUNTER.counter_1_cry_21 ),
            .clk(N__33022),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_22_LC_1_15_5 .C_ON=1'b1;
    defparam \COUNTER.counter_22_LC_1_15_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_22_LC_1_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_22_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__16384),
            .in2(_gnd_net_),
            .in3(N__14395),
            .lcout(\COUNTER.counterZ0Z_22 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_21 ),
            .carryout(\COUNTER.counter_1_cry_22 ),
            .clk(N__33022),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_23_LC_1_15_6 .C_ON=1'b1;
    defparam \COUNTER.counter_23_LC_1_15_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_23_LC_1_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_23_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(N__16359),
            .in2(_gnd_net_),
            .in3(N__14392),
            .lcout(\COUNTER.counterZ0Z_23 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_22 ),
            .carryout(\COUNTER.counter_1_cry_23 ),
            .clk(N__33022),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_24_LC_1_15_7 .C_ON=1'b1;
    defparam \COUNTER.counter_24_LC_1_15_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_24_LC_1_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_24_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__16270),
            .in2(_gnd_net_),
            .in3(N__14389),
            .lcout(\COUNTER.counterZ0Z_24 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_23 ),
            .carryout(\COUNTER.counter_1_cry_24 ),
            .clk(N__33022),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_25_LC_1_16_0 .C_ON=1'b1;
    defparam \COUNTER.counter_25_LC_1_16_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_25_LC_1_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_25_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__16282),
            .in2(_gnd_net_),
            .in3(N__14386),
            .lcout(\COUNTER.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\COUNTER.counter_1_cry_25 ),
            .clk(N__33064),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_26_LC_1_16_1 .C_ON=1'b1;
    defparam \COUNTER.counter_26_LC_1_16_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_26_LC_1_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_26_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__16257),
            .in2(_gnd_net_),
            .in3(N__14383),
            .lcout(\COUNTER.counterZ0Z_26 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_25 ),
            .carryout(\COUNTER.counter_1_cry_26 ),
            .clk(N__33064),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_27_LC_1_16_2 .C_ON=1'b1;
    defparam \COUNTER.counter_27_LC_1_16_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_27_LC_1_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_27_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(N__16243),
            .in2(_gnd_net_),
            .in3(N__14380),
            .lcout(\COUNTER.counterZ0Z_27 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_26 ),
            .carryout(\COUNTER.counter_1_cry_27 ),
            .clk(N__33064),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_28_LC_1_16_3 .C_ON=1'b1;
    defparam \COUNTER.counter_28_LC_1_16_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_28_LC_1_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_28_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(N__16333),
            .in2(_gnd_net_),
            .in3(N__14377),
            .lcout(\COUNTER.counterZ0Z_28 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_27 ),
            .carryout(\COUNTER.counter_1_cry_28 ),
            .clk(N__33064),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_29_LC_1_16_4 .C_ON=1'b1;
    defparam \COUNTER.counter_29_LC_1_16_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_29_LC_1_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_29_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(N__16308),
            .in2(_gnd_net_),
            .in3(N__14374),
            .lcout(\COUNTER.counterZ0Z_29 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_28 ),
            .carryout(\COUNTER.counter_1_cry_29 ),
            .clk(N__33064),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_30_LC_1_16_5 .C_ON=1'b1;
    defparam \COUNTER.counter_30_LC_1_16_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_30_LC_1_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_30_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(N__16321),
            .in2(_gnd_net_),
            .in3(N__14470),
            .lcout(\COUNTER.counterZ0Z_30 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_29 ),
            .carryout(\COUNTER.counter_1_cry_30 ),
            .clk(N__33064),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_31_LC_1_16_6 .C_ON=1'b0;
    defparam \COUNTER.counter_31_LC_1_16_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_31_LC_1_16_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.counter_31_LC_1_16_6  (
            .in0(_gnd_net_),
            .in1(N__16294),
            .in2(_gnd_net_),
            .in3(N__14467),
            .lcout(\COUNTER.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33064),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_0_LC_2_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_0_LC_2_1_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_0_LC_2_1_0 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \PCH_PWRGD.count_0_LC_2_1_0  (
            .in0(N__14725),
            .in1(N__20930),
            .in2(N__14415),
            .in3(N__14529),
            .lcout(\PCH_PWRGD.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32800),
            .ce(N__21146),
            .sr(N__20976));
    defparam \PCH_PWRGD.count_RNIRP9H1_1_LC_2_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIRP9H1_1_LC_2_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIRP9H1_1_LC_2_1_1 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \PCH_PWRGD.count_RNIRP9H1_1_LC_2_1_1  (
            .in0(N__14461),
            .in1(_gnd_net_),
            .in2(N__20972),
            .in3(N__14432),
            .lcout(\PCH_PWRGD.count_rst_13 ),
            .ltout(\PCH_PWRGD.count_rst_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNILOMR3_1_LC_2_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNILOMR3_1_LC_2_1_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNILOMR3_1_LC_2_1_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.count_RNILOMR3_1_LC_2_1_2  (
            .in0(_gnd_net_),
            .in1(N__14565),
            .in2(N__14464),
            .in3(N__21126),
            .lcout(\PCH_PWRGD.un2_count_1_axb_1 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_1_LC_2_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_1_LC_2_1_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_1_LC_2_1_3 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \PCH_PWRGD.count_1_LC_2_1_3  (
            .in0(N__20929),
            .in1(_gnd_net_),
            .in2(N__14449),
            .in3(N__14433),
            .lcout(\PCH_PWRGD.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32800),
            .ce(N__21146),
            .sr(N__20976));
    defparam \PCH_PWRGD.count_RNI6HKKG_1_LC_2_1_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI6HKKG_1_LC_2_1_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI6HKKG_1_LC_2_1_4 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \PCH_PWRGD.count_RNI6HKKG_1_LC_2_1_4  (
            .in0(N__14724),
            .in1(N__20925),
            .in2(N__14416),
            .in3(N__14528),
            .lcout(),
            .ltout(\PCH_PWRGD.count_RNI6HKKGZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIVE1VI_0_LC_2_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIVE1VI_0_LC_2_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIVE1VI_0_LC_2_1_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNIVE1VI_0_LC_2_1_5  (
            .in0(N__21125),
            .in1(_gnd_net_),
            .in2(N__14446),
            .in3(N__14443),
            .lcout(\PCH_PWRGD.countZ0Z_0 ),
            .ltout(\PCH_PWRGD.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI_0_LC_2_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI_0_LC_2_1_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI_0_LC_2_1_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \PCH_PWRGD.count_RNI_0_LC_2_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14419),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.N_2093_i ),
            .ltout(\PCH_PWRGD.N_2093_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIBNA3F_0_1_LC_2_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIBNA3F_0_1_LC_2_1_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIBNA3F_0_1_LC_2_1_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \PCH_PWRGD.count_RNIBNA3F_0_1_LC_2_1_7  (
            .in0(N__14530),
            .in1(_gnd_net_),
            .in2(N__14584),
            .in3(N__14723),
            .lcout(\PCH_PWRGD.N_540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIELSI2_0_14_LC_2_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIELSI2_0_14_LC_2_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIELSI2_0_14_LC_2_2_0 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \PCH_PWRGD.count_RNIELSI2_0_14_LC_2_2_0  (
            .in0(N__21151),
            .in1(N__14500),
            .in2(N__14518),
            .in3(N__14581),
            .lcout(\PCH_PWRGD.count_1_i_a2_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNILOMR3_0_1_LC_2_2_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNILOMR3_0_1_LC_2_2_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNILOMR3_0_1_LC_2_2_1 .LUT_INIT=16'b0000001100010001;
    LogicCell40 \PCH_PWRGD.count_RNILOMR3_0_1_LC_2_2_1  (
            .in0(N__14566),
            .in1(N__16597),
            .in2(N__14554),
            .in3(N__21152),
            .lcout(),
            .ltout(\PCH_PWRGD.count_1_i_a2_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIBNA3F_1_LC_2_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIBNA3F_1_LC_2_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIBNA3F_1_LC_2_2_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNIBNA3F_1_LC_2_2_2  (
            .in0(N__14545),
            .in1(N__14539),
            .in2(N__14533),
            .in3(N__14488),
            .lcout(\PCH_PWRGD.count_1_i_a2_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_14_LC_2_2_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_14_LC_2_2_4 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_14_LC_2_2_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_14_LC_2_2_4  (
            .in0(N__14514),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32651),
            .ce(N__21150),
            .sr(N__21005));
    defparam \PCH_PWRGD.count_RNIEGTB4_0_11_LC_2_2_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIEGTB4_0_11_LC_2_2_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIEGTB4_0_11_LC_2_2_5 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \PCH_PWRGD.count_RNIEGTB4_0_11_LC_2_2_5  (
            .in0(N__14478),
            .in1(N__21112),
            .in2(N__14665),
            .in3(N__14618),
            .lcout(\PCH_PWRGD.count_1_i_a2_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIEGTB4_11_LC_2_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIEGTB4_11_LC_2_2_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIEGTB4_11_LC_2_2_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \PCH_PWRGD.count_RNIEGTB4_11_LC_2_2_6  (
            .in0(N__21113),
            .in1(N__14479),
            .in2(_gnd_net_),
            .in3(N__14661),
            .lcout(\PCH_PWRGD.un2_count_1_axb_11 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_11_LC_2_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_11_LC_2_2_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_11_LC_2_2_7 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \PCH_PWRGD.count_11_LC_2_2_7  (
            .in0(N__20971),
            .in1(N__15003),
            .in2(N__14482),
            .in3(N__14677),
            .lcout(\PCH_PWRGD.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32651),
            .ce(N__21150),
            .sr(N__21005));
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNI3U0P1_LC_2_3_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNI3U0P1_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNI3U0P1_LC_2_3_0 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_c_RNI3U0P1_LC_2_3_0  (
            .in0(N__15006),
            .in1(N__14689),
            .in2(N__20947),
            .in3(N__14676),
            .lcout(\PCH_PWRGD.count_rst_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIMC9U1_LC_2_3_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIMC9U1_LC_2_3_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIMC9U1_LC_2_3_1 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_c_RNIMC9U1_LC_2_3_1  (
            .in0(N__14801),
            .in1(N__14649),
            .in2(N__20965),
            .in3(N__15005),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIKFM84_5_LC_2_3_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIKFM84_5_LC_2_3_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIKFM84_5_LC_2_3_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNIKFM84_5_LC_2_3_2  (
            .in0(N__21073),
            .in1(_gnd_net_),
            .in2(N__14638),
            .in3(N__14635),
            .lcout(\PCH_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIQKDU1_LC_2_3_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIQKDU1_LC_2_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIQKDU1_LC_2_3_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_c_RNIQKDU1_LC_2_3_3  (
            .in0(N__14602),
            .in1(N__20892),
            .in2(N__14623),
            .in3(N__15004),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNISRQ84_9_LC_2_3_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNISRQ84_9_LC_2_3_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNISRQ84_9_LC_2_3_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNISRQ84_9_LC_2_3_4  (
            .in0(N__21072),
            .in1(_gnd_net_),
            .in2(N__14626),
            .in3(N__14590),
            .lcout(\PCH_PWRGD.countZ0Z_9 ),
            .ltout(\PCH_PWRGD.countZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_9_LC_2_3_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_9_LC_2_3_5 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_9_LC_2_3_5 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.count_9_LC_2_3_5  (
            .in0(N__14601),
            .in1(N__20998),
            .in2(N__14593),
            .in3(N__15007),
            .lcout(\PCH_PWRGD.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32875),
            .ce(N__21076),
            .sr(N__20997));
    defparam \PCH_PWRGD.count_RNIGJUB4_12_LC_2_3_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIGJUB4_12_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIGJUB4_12_LC_2_3_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \PCH_PWRGD.count_RNIGJUB4_12_LC_2_3_6  (
            .in0(N__21075),
            .in1(_gnd_net_),
            .in2(N__14698),
            .in3(N__14709),
            .lcout(\PCH_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIMIN84_6_LC_2_3_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIMIN84_6_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIMIN84_6_LC_2_3_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \PCH_PWRGD.count_RNIMIN84_6_LC_2_3_7  (
            .in0(N__21172),
            .in1(N__21074),
            .in2(_gnd_net_),
            .in3(N__21183),
            .lcout(\PCH_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_2_LC_2_4_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_2_LC_2_4_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_2_LC_2_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_2_LC_2_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14884),
            .lcout(\PCH_PWRGD.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32652),
            .ce(N__21097),
            .sr(N__21010));
    defparam \PCH_PWRGD.count_10_LC_2_4_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_10_LC_2_4_1 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_10_LC_2_4_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_10_LC_2_4_1  (
            .in0(N__14860),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32652),
            .ce(N__21097),
            .sr(N__21010));
    defparam \PCH_PWRGD.count_RNIE6J84_2_LC_2_4_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIE6J84_2_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIE6J84_2_LC_2_4_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \PCH_PWRGD.count_RNIE6J84_2_LC_2_4_2  (
            .in0(N__21096),
            .in1(N__14890),
            .in2(_gnd_net_),
            .in3(N__14883),
            .lcout(\PCH_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNISDK72_0_LC_2_4_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNISDK72_0_LC_2_4_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNISDK72_0_LC_2_4_3 .LUT_INIT=16'b1010101100000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNISDK72_0_LC_2_4_3  (
            .in0(N__20891),
            .in1(N__14908),
            .in2(N__16508),
            .in3(N__28142),
            .lcout(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ),
            .ltout(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI58BH4_10_LC_2_4_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI58BH4_10_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI58BH4_10_LC_2_4_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \PCH_PWRGD.count_RNI58BH4_10_LC_2_4_4  (
            .in0(_gnd_net_),
            .in1(N__14869),
            .in2(N__14863),
            .in3(N__14859),
            .lcout(\PCH_PWRGD.countZ0Z_10 ),
            .ltout(\PCH_PWRGD.countZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI_2_LC_2_4_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI_2_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI_2_LC_2_4_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \PCH_PWRGD.count_RNI_2_LC_2_4_5  (
            .in0(N__14844),
            .in1(N__14830),
            .in2(N__14818),
            .in3(N__14815),
            .lcout(),
            .ltout(\PCH_PWRGD.count_1_i_a2_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI_3_LC_2_4_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI_3_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI_3_LC_2_4_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNI_3_LC_2_4_6  (
            .in0(N__14802),
            .in1(N__14776),
            .in2(N__14752),
            .in3(N__14747),
            .lcout(\PCH_PWRGD.count_1_i_a2_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_12_LC_2_4_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_12_LC_2_4_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_12_LC_2_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_12_LC_2_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14710),
            .lcout(\PCH_PWRGD.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32652),
            .ce(N__21097),
            .sr(N__21010));
    defparam \PCH_PWRGD.curr_state_0_LC_2_5_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_0_LC_2_5_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_0_LC_2_5_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \PCH_PWRGD.curr_state_0_LC_2_5_0  (
            .in0(N__14925),
            .in1(N__16484),
            .in2(N__15024),
            .in3(N__19478),
            .lcout(\PCH_PWRGD.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32978),
            .ce(N__32290),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_1_LC_2_5_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_1_LC_2_5_1 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_1_LC_2_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \PCH_PWRGD.curr_state_1_LC_2_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14941),
            .lcout(\PCH_PWRGD.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32978),
            .ce(N__32290),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_2_5_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_2_5_2 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_2_5_2  (
            .in0(N__14926),
            .in1(N__19477),
            .in2(N__15025),
            .in3(N__16485),
            .lcout(),
            .ltout(\PCH_PWRGD.curr_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIB48V1_0_LC_2_5_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIB48V1_0_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIB48V1_0_LC_2_5_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.curr_state_RNIB48V1_0_LC_2_5_3  (
            .in0(_gnd_net_),
            .in1(N__15037),
            .in2(N__15031),
            .in3(N__33877),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_0 ),
            .ltout(\PCH_PWRGD.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_LC_2_5_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_LC_2_5_4 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m6_i_LC_2_5_4  (
            .in0(N__14924),
            .in1(N__14907),
            .in2(N__15028),
            .in3(N__15017),
            .lcout(\PCH_PWRGD.N_205 ),
            .ltout(\PCH_PWRGD.N_205_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIVGBJ_1_LC_2_5_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIVGBJ_1_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIVGBJ_1_LC_2_5_5 .LUT_INIT=16'b0000111111001100;
    LogicCell40 \PCH_PWRGD.curr_state_RNIVGBJ_1_LC_2_5_5  (
            .in0(_gnd_net_),
            .in1(N__14935),
            .in2(N__14929),
            .in3(N__33878),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_1 ),
            .ltout(\PCH_PWRGD.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_2_5_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_2_5_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_1_LC_2_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14914),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.N_2110_i ),
            .ltout(\PCH_PWRGD.N_2110_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIRP9H1_0_LC_2_5_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIRP9H1_0_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIRP9H1_0_LC_2_5_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNIRP9H1_0_LC_2_5_7  (
            .in0(N__16483),
            .in1(N__16536),
            .in2(N__14911),
            .in3(N__33879),
            .lcout(\PCH_PWRGD.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_LC_2_6_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_LC_2_6_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(N__15184),
            .in2(_gnd_net_),
            .in3(N__25008),
            .lcout(N_355),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIDKSB1_1_LC_2_6_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIDKSB1_1_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIDKSB1_1_LC_2_6_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNIDKSB1_1_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(N__16548),
            .in2(_gnd_net_),
            .in3(N__16535),
            .lcout(\PCH_PWRGD.N_562 ),
            .ltout(\PCH_PWRGD.N_562_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_0_0_LC_2_6_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_0_0_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_0_0_LC_2_6_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_0_0_LC_2_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14893),
            .in3(N__16486),
            .lcout(\PCH_PWRGD.N_38_f0 ),
            .ltout(\PCH_PWRGD.N_38_f0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIT2822_LC_2_6_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIT2822_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIT2822_LC_2_6_3 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNIT2822_LC_2_6_3  (
            .in0(N__19441),
            .in1(N__32316),
            .in2(N__15187),
            .in3(N__19479),
            .lcout(\PCH_PWRGD.delayed_vccin_okZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_2_6_4 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_2_6_4 .LUT_INIT=16'b0000001001010010;
    LogicCell40 \HDA_STRAP.curr_state_RNO_0_0_LC_2_6_4  (
            .in0(N__15221),
            .in1(N__15178),
            .in2(N__15255),
            .in3(N__15293),
            .lcout(),
            .ltout(\HDA_STRAP.m14_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_0_LC_2_6_5 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_0_LC_2_6_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_0_LC_2_6_5 .LUT_INIT=16'b1111000011111001;
    LogicCell40 \HDA_STRAP.curr_state_0_LC_2_6_5  (
            .in0(N__15250),
            .in1(N__15222),
            .in2(N__15160),
            .in3(N__20770),
            .lcout(\HDA_STRAP.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32762),
            .ce(N__27381),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIH91A_0_LC_2_6_6 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIH91A_0_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIH91A_0_LC_2_6_6 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \HDA_STRAP.curr_state_RNIH91A_0_LC_2_6_6  (
            .in0(N__15220),
            .in1(_gnd_net_),
            .in2(N__15254),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.N_336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIH91A_0_0_LC_2_6_7 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIH91A_0_0_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIH91A_0_0_LC_2_6_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \HDA_STRAP.curr_state_RNIH91A_0_0_LC_2_6_7  (
            .in0(_gnd_net_),
            .in1(N__15219),
            .in2(_gnd_net_),
            .in3(N__15243),
            .lcout(\HDA_STRAP.curr_state_RNIH91A_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_2_7_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_2_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \HDA_STRAP.count_RNIBJB61_7_LC_2_7_0  (
            .in0(N__15156),
            .in1(N__15144),
            .in2(N__15133),
            .in3(N__15117),
            .lcout(\HDA_STRAP.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_2_7_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_2_7_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \HDA_STRAP.count_RNIDLB61_6_LC_2_7_1  (
            .in0(N__15093),
            .in1(N__15428),
            .in2(N__15055),
            .in3(N__15081),
            .lcout(\HDA_STRAP.un4_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_6_LC_2_7_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_6_LC_2_7_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_6_LC_2_7_2 .LUT_INIT=16'b0000011001100110;
    LogicCell40 \HDA_STRAP.count_6_LC_2_7_2  (
            .in0(N__15061),
            .in1(N__15054),
            .in2(N__15415),
            .in3(N__15305),
            .lcout(\HDA_STRAP.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32884),
            .ce(N__27380),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_8_LC_2_7_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_8_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_8_LC_2_7_3 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \HDA_STRAP.count_8_LC_2_7_3  (
            .in0(N__15304),
            .in1(N__15429),
            .in2(N__15399),
            .in3(N__15439),
            .lcout(\HDA_STRAP.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32884),
            .ce(N__27380),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_2_7_4 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_2_7_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \HDA_STRAP.curr_state_RNO_0_2_LC_2_7_4  (
            .in0(_gnd_net_),
            .in1(N__15376),
            .in2(_gnd_net_),
            .in3(N__15302),
            .lcout(),
            .ltout(\HDA_STRAP.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_2_LC_2_7_5 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_2_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_2_LC_2_7_5 .LUT_INIT=16'b0000101000001110;
    LogicCell40 \HDA_STRAP.curr_state_2_LC_2_7_5  (
            .in0(N__15331),
            .in1(N__20772),
            .in2(N__15343),
            .in3(N__15340),
            .lcout(\HDA_STRAP.curr_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32884),
            .ce(N__27380),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_2_7_6 .C_ON=1'b0;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_2_7_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_2_7_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \HDA_STRAP.HDA_SDO_ATP_LC_2_7_6  (
            .in0(N__15339),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15330),
            .lcout(hda_sdo_atp),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32884),
            .ce(N__27380),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_1_LC_2_7_7 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_1_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_1_LC_2_7_7 .LUT_INIT=16'b0011111110100000;
    LogicCell40 \HDA_STRAP.curr_state_1_LC_2_7_7  (
            .in0(N__15303),
            .in1(N__20771),
            .in2(N__15259),
            .in3(N__15223),
            .lcout(\HDA_STRAP.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32884),
            .ce(N__27380),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_0_sqmuxa_0_o2_1_LC_2_8_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_0_sqmuxa_0_o2_1_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_0_sqmuxa_0_o2_1_LC_2_8_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \PCH_PWRGD.count_0_sqmuxa_0_o2_1_LC_2_8_3  (
            .in0(N__15202),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24999),
            .lcout(\PCH_PWRGD.N_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_2_LC_2_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_2_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_2_LC_2_9_0 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \POWERLED.count_clk_RNI_2_LC_2_9_0  (
            .in0(N__16120),
            .in1(N__15744),
            .in2(N__15709),
            .in3(N__15669),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_168_0_0_o3_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_3_LC_2_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_3_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_3_LC_2_9_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNI_3_LC_2_9_1  (
            .in0(N__15592),
            .in1(N__15479),
            .in2(N__15190),
            .in3(N__15507),
            .lcout(\POWERLED.N_335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_3_LC_2_9_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_3_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_3_LC_2_9_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_3_LC_2_9_2  (
            .in0(N__15529),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33023),
            .ce(N__16933),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI168J_3_LC_2_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI168J_3_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI168J_3_LC_2_9_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNI168J_3_LC_2_9_3  (
            .in0(N__33880),
            .in1(N__15528),
            .in2(N__15517),
            .in3(N__16896),
            .lcout(\POWERLED.count_clkZ0Z_3 ),
            .ltout(\POWERLED.count_clkZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_2_LC_2_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_2_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_2_LC_2_9_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \POWERLED.count_clk_RNI_0_2_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15487),
            .in3(N__15670),
            .lcout(),
            .ltout(\POWERLED.un1_count_clk_1_sqmuxa_i_i_a2_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_4_LC_2_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_4_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_4_LC_2_9_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.count_clk_RNI_4_LC_2_9_5  (
            .in0(N__15745),
            .in1(N__15480),
            .in2(N__15463),
            .in3(N__15708),
            .lcout(\POWERLED.N_515 ),
            .ltout(\POWERLED.N_515_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_7_LC_2_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_7_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_7_LC_2_9_6 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \POWERLED.count_clk_RNI_7_LC_2_9_6  (
            .in0(N__16119),
            .in1(_gnd_net_),
            .in2(N__15460),
            .in3(N__15591),
            .lcout(\POWERLED.count_clk_RNIZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_9_LC_2_9_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_9_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_9_LC_2_9_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.count_clk_RNI_9_LC_2_9_7  (
            .in0(N__15610),
            .in1(N__15556),
            .in2(N__15457),
            .in3(N__16118),
            .lcout(\POWERLED.count_clk_RNIZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIDPQG4_1_LC_2_10_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIDPQG4_1_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIDPQG4_1_LC_2_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.func_state_RNIDPQG4_1_LC_2_10_0  (
            .in0(N__15616),
            .in1(N__15622),
            .in2(N__18427),
            .in3(N__15628),
            .lcout(\POWERLED.N_47_i ),
            .ltout(\POWERLED.N_47_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_0_LC_2_10_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_0_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_0_LC_2_10_1 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \POWERLED.count_clk_RNI_0_0_LC_2_10_1  (
            .in0(N__15825),
            .in1(_gnd_net_),
            .in2(N__15448),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.count_clk_RNI_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI8LLG_0_LC_2_10_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI8LLG_0_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI8LLG_0_LC_2_10_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \POWERLED.count_clk_RNI8LLG_0_LC_2_10_2  (
            .in0(N__15634),
            .in1(N__33900),
            .in2(N__15445),
            .in3(N__16921),
            .lcout(\POWERLED.count_clkZ0Z_0 ),
            .ltout(\POWERLED.count_clkZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_1_LC_2_10_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_1_LC_2_10_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_1_LC_2_10_3 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \POWERLED.count_clk_1_LC_2_10_3  (
            .in0(N__15789),
            .in1(_gnd_net_),
            .in2(N__15442),
            .in3(N__15883),
            .lcout(\POWERLED.count_clk_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32874),
            .ce(N__16925),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_0_LC_2_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_0_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_0_LC_2_10_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.count_clk_0_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__15882),
            .in2(_gnd_net_),
            .in3(N__15824),
            .lcout(\POWERLED.count_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32874),
            .ce(N__16925),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_1_LC_2_10_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_1_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_1_LC_2_10_5 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \POWERLED.func_state_RNI5DLR_1_LC_2_10_5  (
            .in0(N__28863),
            .in1(N__18235),
            .in2(N__26731),
            .in3(N__18449),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_0_1_LC_2_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_0_1_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_0_1_LC_2_10_6 .LUT_INIT=16'b0100010001001110;
    LogicCell40 \POWERLED.func_state_RNI5DLR_0_1_LC_2_10_6  (
            .in0(N__26726),
            .in1(N__18251),
            .in2(N__30698),
            .in3(N__28862),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_i_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_3_1_LC_2_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_3_1_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_3_1_LC_2_10_7 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \POWERLED.func_state_RNI5DLR_3_1_LC_2_10_7  (
            .in0(N__30571),
            .in1(N__16786),
            .in2(N__30391),
            .in3(N__19906),
            .lcout(\POWERLED.N_415 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIDOEJ_9_LC_2_11_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIDOEJ_9_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIDOEJ_9_LC_2_11_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNIDOEJ_9_LC_2_11_0  (
            .in0(N__33910),
            .in1(N__15762),
            .in2(N__15754),
            .in3(N__16928),
            .lcout(\POWERLED.count_clkZ0Z_9 ),
            .ltout(\POWERLED.count_clkZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_1_LC_2_11_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_1_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_1_LC_2_11_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \POWERLED.count_clk_RNI_1_LC_2_11_1  (
            .in0(N__15580),
            .in1(N__15568),
            .in2(N__15595),
            .in3(N__15783),
            .lcout(\POWERLED.N_320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI5CAJ_5_LC_2_11_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI5CAJ_5_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI5CAJ_5_LC_2_11_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNI5CAJ_5_LC_2_11_2  (
            .in0(N__33909),
            .in1(N__15546),
            .in2(N__15538),
            .in3(N__16927),
            .lcout(\POWERLED.count_clkZ0Z_5 ),
            .ltout(\POWERLED.count_clkZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_1_LC_2_11_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_1_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_1_LC_2_11_3 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_1_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__15567),
            .in2(N__15559),
            .in3(N__15784),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_i_i_a2_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_5_LC_2_11_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_5_LC_2_11_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_5_LC_2_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_5_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15547),
            .lcout(\POWERLED.count_clk_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32973),
            .ce(N__16929),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_LC_2_11_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_LC_2_11_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.count_clk_RNI_0_LC_2_11_5  (
            .in0(N__15884),
            .in1(N__15822),
            .in2(_gnd_net_),
            .in3(N__15785),
            .lcout(),
            .ltout(\POWERLED.count_clk_RNIZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI9MLG_1_LC_2_11_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI9MLG_1_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI9MLG_1_LC_2_11_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \POWERLED.count_clk_RNI9MLG_1_LC_2_11_6  (
            .in0(N__15799),
            .in1(N__33901),
            .in2(N__15793),
            .in3(N__16926),
            .lcout(\POWERLED.count_clkZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_9_LC_2_11_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_9_LC_2_11_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_9_LC_2_11_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_9_LC_2_11_7  (
            .in0(N__15763),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32973),
            .ce(N__16929),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI7FBJ_6_LC_2_12_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI7FBJ_6_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI7FBJ_6_LC_2_12_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNI7FBJ_6_LC_2_12_0  (
            .in0(N__33850),
            .in1(N__15726),
            .in2(N__15718),
            .in3(N__16918),
            .lcout(\POWERLED.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_6_LC_2_12_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_6_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_6_LC_2_12_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_6_LC_2_12_1  (
            .in0(N__15727),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33043),
            .ce(N__16936),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIBLDJ_8_LC_2_12_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIBLDJ_8_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIBLDJ_8_LC_2_12_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNIBLDJ_8_LC_2_12_2  (
            .in0(N__33851),
            .in1(N__15687),
            .in2(N__15679),
            .in3(N__16919),
            .lcout(\POWERLED.count_clkZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_8_LC_2_12_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_8_LC_2_12_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_8_LC_2_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_8_LC_2_12_3  (
            .in0(N__15688),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33043),
            .ce(N__16936),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIV27J_2_LC_2_12_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIV27J_2_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIV27J_2_LC_2_12_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNIV27J_2_LC_2_12_4  (
            .in0(N__33849),
            .in1(N__15651),
            .in2(N__15643),
            .in3(N__16917),
            .lcout(\POWERLED.count_clkZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_2_LC_2_12_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_2_LC_2_12_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_2_LC_2_12_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_2_LC_2_12_5  (
            .in0(N__15652),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33043),
            .ce(N__16936),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI9ICJ_7_LC_2_12_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI9ICJ_7_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI9ICJ_7_LC_2_12_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \POWERLED.count_clk_RNI9ICJ_7_LC_2_12_6  (
            .in0(N__16087),
            .in1(N__33826),
            .in2(N__16099),
            .in3(N__16916),
            .lcout(\POWERLED.count_clkZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_7_LC_2_12_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_7_LC_2_12_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_7_LC_2_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_7_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16095),
            .lcout(\POWERLED.count_clk_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33043),
            .ce(N__16936),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_LC_2_13_2 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_LC_2_13_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_LC_2_13_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.tmp_0_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__33861),
            .in2(_gnd_net_),
            .in3(N__21748),
            .lcout(suswarn_n),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33060),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_vddq_en_LC_2_13_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_vddq_en_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_vddq_en_LC_2_13_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \VPP_VDDQ.un1_vddq_en_LC_2_13_6  (
            .in0(N__16081),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23384),
            .lcout(vddq_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_RNO_LC_2_14_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_2_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_2_c_RNO_LC_2_14_0  (
            .in0(N__16059),
            .in1(N__16047),
            .in2(N__16036),
            .in3(N__16020),
            .lcout(\COUNTER.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_RNO_LC_2_14_1 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_2_14_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_3_c_RNO_LC_2_14_1  (
            .in0(N__16008),
            .in1(N__15996),
            .in2(N__15985),
            .in3(N__15969),
            .lcout(\COUNTER.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_RNO_LC_2_14_2 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_2_14_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_4_c_RNO_LC_2_14_2  (
            .in0(N__15957),
            .in1(N__15945),
            .in2(N__15934),
            .in3(N__15918),
            .lcout(\COUNTER.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIH71P_2_LC_2_14_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIH71P_2_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIH71P_2_LC_2_14_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DSW_PWRGD.count_RNIH71P_2_LC_2_14_3  (
            .in0(N__17497),
            .in1(N__17191),
            .in2(N__17173),
            .in3(N__17533),
            .lcout(\DSW_PWRGD.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIKA1P_1_LC_2_14_4 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIKA1P_1_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIKA1P_1_LC_2_14_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DSW_PWRGD.count_RNIKA1P_1_LC_2_14_4  (
            .in0(N__17212),
            .in1(N__17515),
            .in2(N__17149),
            .in3(N__17458),
            .lcout(\DSW_PWRGD.un4_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIBCB91_0_LC_2_15_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIBCB91_0_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIBCB91_0_LC_2_15_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \DSW_PWRGD.count_RNIBCB91_0_LC_2_15_0  (
            .in0(N__17437),
            .in1(N__17476),
            .in2(N__17233),
            .in3(N__17419),
            .lcout(\DSW_PWRGD.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.DSW_PWROK_LC_2_15_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.DSW_PWROK_LC_2_15_1 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.DSW_PWROK_LC_2_15_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \DSW_PWRGD.DSW_PWROK_LC_2_15_1  (
            .in0(N__16144),
            .in1(N__16188),
            .in2(_gnd_net_),
            .in3(N__16165),
            .lcout(dsw_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32963),
            .ce(N__27398),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_RNIADII_0_LC_2_15_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_RNIADII_0_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_RNIADII_0_LC_2_15_2 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \DSW_PWRGD.curr_state_RNIADII_0_LC_2_15_2  (
            .in0(N__16161),
            .in1(N__16191),
            .in2(_gnd_net_),
            .in3(N__16140),
            .lcout(\DSW_PWRGD.un1_curr_state10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_0_LC_2_15_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_0_LC_2_15_3 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.curr_state_0_LC_2_15_3 .LUT_INIT=16'b0100010010100000;
    LogicCell40 \DSW_PWRGD.curr_state_0_LC_2_15_3  (
            .in0(N__16145),
            .in1(N__16189),
            .in2(N__16405),
            .in3(N__16164),
            .lcout(\DSW_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32963),
            .ce(N__27398),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_1_LC_2_15_4 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_1_LC_2_15_4 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.curr_state_1_LC_2_15_4 .LUT_INIT=16'b0000010101000100;
    LogicCell40 \DSW_PWRGD.curr_state_1_LC_2_15_4  (
            .in0(N__16163),
            .in1(N__16190),
            .in2(N__16404),
            .in3(N__16146),
            .lcout(\DSW_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32963),
            .ce(N__27398),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_RNILLF15_0_LC_2_15_5 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_RNILLF15_0_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_RNILLF15_0_LC_2_15_5 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \DSW_PWRGD.curr_state_RNILLF15_0_LC_2_15_5  (
            .in0(N__16192),
            .in1(N__16162),
            .in2(N__16147),
            .in3(N__16397),
            .lcout(),
            .ltout(DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_28_LC_2_15_6 .C_ON=1'b0;
    defparam \POWERLED.G_28_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_28_LC_2_15_6 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \POWERLED.G_28_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16126),
            .in3(N__27526),
            .lcout(G_28),
            .ltout(G_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_esr_RNO_0_15_LC_2_15_7 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_esr_RNO_0_15_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_esr_RNO_0_15_LC_2_15_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \DSW_PWRGD.count_esr_RNO_0_15_LC_2_15_7  (
            .in0(N__27527),
            .in1(_gnd_net_),
            .in2(N__16123),
            .in3(_gnd_net_),
            .lcout(\DSW_PWRGD.N_42_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_16_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_16_0  (
            .in0(N__17401),
            .in1(N__17605),
            .in2(N__17653),
            .in3(N__17629),
            .lcout(),
            .ltout(\DSW_PWRGD.un4_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIB8TE4_0_LC_2_16_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIB8TE4_0_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIB8TE4_0_LC_2_16_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DSW_PWRGD.count_RNIB8TE4_0_LC_2_16_1  (
            .in0(N__16432),
            .in1(N__16426),
            .in2(N__16417),
            .in3(N__16414),
            .lcout(\DSW_PWRGD.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_RNO_LC_2_16_2 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_2_16_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_5_c_RNO_LC_2_16_2  (
            .in0(N__16383),
            .in1(N__16371),
            .in2(N__16360),
            .in3(N__16344),
            .lcout(\COUNTER.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_RNO_LC_2_16_3 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_2_16_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_7_c_RNO_LC_2_16_3  (
            .in0(N__16332),
            .in1(N__16320),
            .in2(N__16309),
            .in3(N__16293),
            .lcout(\COUNTER.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_RNO_LC_2_16_4 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_2_16_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_6_c_RNO_LC_2_16_4  (
            .in0(N__16281),
            .in1(N__16269),
            .in2(N__16258),
            .in3(N__16242),
            .lcout(\COUNTER.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNI1KAM_0_LC_4_1_0 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI1KAM_0_LC_4_1_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI1KAM_0_LC_4_1_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \POWERLED.curr_state_RNI1KAM_0_LC_4_1_0  (
            .in0(_gnd_net_),
            .in1(N__32319),
            .in2(_gnd_net_),
            .in3(N__22382),
            .lcout(\POWERLED.g0_i_o3_0 ),
            .ltout(\POWERLED.g0_i_o3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_LC_4_1_1 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_LC_4_1_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.pwm_out_LC_4_1_1 .LUT_INIT=16'b0010001100100010;
    LogicCell40 \POWERLED.pwm_out_LC_4_1_1  (
            .in0(N__16227),
            .in1(N__17721),
            .in2(N__16231),
            .in3(N__22421),
            .lcout(\POWERLED.pwm_outZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32549),
            .ce(),
            .sr(N__17728));
    defparam \POWERLED.pwm_out_RNIB7P12_LC_4_1_2 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNIB7P12_LC_4_1_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNIB7P12_LC_4_1_2 .LUT_INIT=16'b0100010001010100;
    LogicCell40 \POWERLED.pwm_out_RNIB7P12_LC_4_1_2  (
            .in0(N__17722),
            .in1(N__16228),
            .in2(N__22426),
            .in3(N__16219),
            .lcout(pwrbtn_led),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_4_1_3 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_4_1_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_4_1_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_4_1_3  (
            .in0(N__22383),
            .in1(N__22352),
            .in2(_gnd_net_),
            .in3(N__22420),
            .lcout(),
            .ltout(\POWERLED.curr_state_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNI2P6L_0_LC_4_1_4 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI2P6L_0_LC_4_1_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI2P6L_0_LC_4_1_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.curr_state_RNI2P6L_0_LC_4_1_4  (
            .in0(_gnd_net_),
            .in1(N__22333),
            .in2(N__16462),
            .in3(N__33983),
            .lcout(\POWERLED.curr_stateZ0Z_0 ),
            .ltout(\POWERLED.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNIE5D5_0_LC_4_1_5 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNIE5D5_0_LC_4_1_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNIE5D5_0_LC_4_1_5 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \POWERLED.curr_state_RNIE5D5_0_LC_4_1_5  (
            .in0(N__33984),
            .in1(_gnd_net_),
            .in2(N__16459),
            .in3(N__22351),
            .lcout(\POWERLED.count_0_sqmuxa_i ),
            .ltout(\POWERLED.count_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_0_LC_4_1_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_0_LC_4_1_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_0_LC_4_1_6 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \POWERLED.count_RNI_0_LC_4_1_6  (
            .in0(N__18746),
            .in1(_gnd_net_),
            .in2(N__16456),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.count_RNIZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIFAFE_0_LC_4_1_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNIFAFE_0_LC_4_1_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIFAFE_0_LC_4_1_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.count_RNIFAFE_0_LC_4_1_7  (
            .in0(N__33985),
            .in1(_gnd_net_),
            .in2(N__16453),
            .in3(N__16438),
            .lcout(\POWERLED.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_1_LC_4_2_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_1_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_1_LC_4_2_0 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \POWERLED.count_RNI_1_LC_4_2_0  (
            .in0(N__18701),
            .in1(N__18743),
            .in2(_gnd_net_),
            .in3(N__17812),
            .lcout(),
            .ltout(\POWERLED.count_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIGBFE_1_LC_4_2_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNIGBFE_1_LC_4_2_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIGBFE_1_LC_4_2_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.count_RNIGBFE_1_LC_4_2_1  (
            .in0(N__34022),
            .in1(_gnd_net_),
            .in2(N__16450),
            .in3(N__16444),
            .lcout(\POWERLED.countZ0Z_1 ),
            .ltout(\POWERLED.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_1_LC_4_2_2 .C_ON=1'b0;
    defparam \POWERLED.count_1_LC_4_2_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_1_LC_4_2_2 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \POWERLED.count_1_LC_4_2_2  (
            .in0(_gnd_net_),
            .in1(N__18745),
            .in2(N__16447),
            .in3(N__17816),
            .lcout(\POWERLED.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32536),
            .ce(N__32285),
            .sr(_gnd_net_));
    defparam \POWERLED.count_0_LC_4_2_3 .C_ON=1'b0;
    defparam \POWERLED.count_0_LC_4_2_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_0_LC_4_2_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \POWERLED.count_0_LC_4_2_3  (
            .in0(N__18744),
            .in1(_gnd_net_),
            .in2(N__17824),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32536),
            .ce(N__32285),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIUHGN_3_LC_4_2_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNIUHGN_3_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIUHGN_3_LC_4_2_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIUHGN_3_LC_4_2_4  (
            .in0(N__16609),
            .in1(N__34021),
            .in2(_gnd_net_),
            .in3(N__17706),
            .lcout(\POWERLED.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_3_LC_4_2_5 .C_ON=1'b0;
    defparam \POWERLED.count_3_LC_4_2_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_3_LC_4_2_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_3_LC_4_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17710),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32536),
            .ce(N__32285),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIUI5O_12_LC_4_2_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNIUI5O_12_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIUI5O_12_LC_4_2_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNIUI5O_12_LC_4_2_6  (
            .in0(N__17854),
            .in1(N__16603),
            .in2(_gnd_net_),
            .in3(N__34023),
            .lcout(\POWERLED.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_12_LC_4_2_7 .C_ON=1'b0;
    defparam \POWERLED.count_12_LC_4_2_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_12_LC_4_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_12_LC_4_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17853),
            .lcout(\POWERLED.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32536),
            .ce(N__32285),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIMS1C4_15_LC_4_3_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIMS1C4_15_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIMS1C4_15_LC_4_3_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNIMS1C4_15_LC_4_3_0  (
            .in0(N__21154),
            .in1(_gnd_net_),
            .in2(N__16576),
            .in3(N__16561),
            .lcout(\PCH_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_15_LC_4_3_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_15_LC_4_3_1 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_15_LC_4_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_15_LC_4_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16572),
            .lcout(\PCH_PWRGD.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32660),
            .ce(N__21153),
            .sr(N__20978));
    defparam \PCH_PWRGD.curr_state_RNIDKSB1_0_LC_4_3_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIDKSB1_0_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIDKSB1_0_LC_4_3_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \PCH_PWRGD.curr_state_RNIDKSB1_0_LC_4_3_2  (
            .in0(N__16510),
            .in1(N__16555),
            .in2(_gnd_net_),
            .in3(N__16537),
            .lcout(\PCH_PWRGD.curr_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_4_3_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_4_3_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_0_LC_4_3_3  (
            .in0(_gnd_net_),
            .in1(N__16509),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.N_2091_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI0LHN_4_LC_4_3_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI0LHN_4_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI0LHN_4_LC_4_3_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI0LHN_4_LC_4_3_4  (
            .in0(N__16636),
            .in1(N__34024),
            .in2(_gnd_net_),
            .in3(N__17691),
            .lcout(\POWERLED.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI0M6O_13_LC_4_3_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNI0M6O_13_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI0M6O_13_LC_4_3_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \POWERLED.count_RNI0M6O_13_LC_4_3_5  (
            .in0(N__34026),
            .in1(N__17842),
            .in2(_gnd_net_),
            .in3(N__16645),
            .lcout(\POWERLED.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI2OIN_5_LC_4_3_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNI2OIN_5_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI2OIN_5_LC_4_3_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI2OIN_5_LC_4_3_6  (
            .in0(N__16627),
            .in1(N__34025),
            .in2(_gnd_net_),
            .in3(N__17673),
            .lcout(\POWERLED.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI2P7O_14_LC_4_3_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNI2P7O_14_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI2P7O_14_LC_4_3_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNI2P7O_14_LC_4_3_7  (
            .in0(N__34027),
            .in1(N__17737),
            .in2(_gnd_net_),
            .in3(N__17749),
            .lcout(\POWERLED.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_13_LC_4_4_0 .C_ON=1'b0;
    defparam \POWERLED.count_13_LC_4_4_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_13_LC_4_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_13_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17841),
            .lcout(\POWERLED.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32766),
            .ce(N__32288),
            .sr(_gnd_net_));
    defparam \POWERLED.count_4_LC_4_4_1 .C_ON=1'b0;
    defparam \POWERLED.count_4_LC_4_4_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_4_LC_4_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_4_LC_4_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17695),
            .lcout(\POWERLED.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32766),
            .ce(N__32288),
            .sr(_gnd_net_));
    defparam \POWERLED.count_5_LC_4_4_2 .C_ON=1'b0;
    defparam \POWERLED.count_5_LC_4_4_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_5_LC_4_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_5_LC_4_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17677),
            .lcout(\POWERLED.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32766),
            .ce(N__32288),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_5_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_5_0  (
            .in0(_gnd_net_),
            .in1(N__21268),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_5_0_),
            .carryout(\POWERLED.mult1_un138_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_5_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_5_1  (
            .in0(_gnd_net_),
            .in1(N__19372),
            .in2(N__16755),
            .in3(N__16621),
            .lcout(\POWERLED.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_5_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_5_2  (
            .in0(_gnd_net_),
            .in1(N__16751),
            .in2(N__16705),
            .in3(N__16618),
            .lcout(\POWERLED.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_5_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(N__16693),
            .in2(N__17919),
            .in3(N__16615),
            .lcout(\POWERLED.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_5_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(N__17915),
            .in2(N__16684),
            .in3(N__16612),
            .lcout(\POWERLED.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_5_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_5_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_5_5  (
            .in0(N__17996),
            .in1(N__16672),
            .in2(N__16756),
            .in3(N__16711),
            .lcout(\POWERLED.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_5_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_5_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16774),
            .in3(N__16708),
            .lcout(\POWERLED.mult1_un138_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_5_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18081),
            .lcout(\POWERLED.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(N__21250),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_6_0_),
            .carryout(\POWERLED.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(N__19351),
            .in2(N__16662),
            .in3(N__16696),
            .lcout(\POWERLED.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(N__16658),
            .in2(N__17953),
            .in3(N__16687),
            .lcout(\POWERLED.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_6_3  (
            .in0(_gnd_net_),
            .in1(N__17941),
            .in2(N__18090),
            .in3(N__16675),
            .lcout(\POWERLED.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_6_4  (
            .in0(_gnd_net_),
            .in1(N__18086),
            .in2(N__17932),
            .in3(N__16666),
            .lcout(\POWERLED.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_6_5  (
            .in0(N__17911),
            .in1(N__18115),
            .in2(N__16663),
            .in3(N__16765),
            .lcout(\POWERLED.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_6_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18106),
            .in3(N__16762),
            .lcout(\POWERLED.mult1_un131_sum_s_8 ),
            .ltout(\POWERLED.mult1_un131_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_6_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_6_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16759),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIF2ST9_4_LC_4_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIF2ST9_4_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIF2ST9_4_LC_4_9_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \POWERLED.count_off_RNIF2ST9_4_LC_4_9_0  (
            .in0(N__20326),
            .in1(N__20196),
            .in2(N__16732),
            .in3(N__20606),
            .lcout(\POWERLED.count_offZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2O4A1_1_LC_4_9_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2O4A1_1_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2O4A1_1_LC_4_9_1 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \POWERLED.func_state_RNI2O4A1_1_LC_4_9_1  (
            .in0(N__24813),
            .in1(_gnd_net_),
            .in2(N__21828),
            .in3(N__28818),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_0_sqmuxa_4_i_0_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBITL2_0_LC_4_9_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBITL2_0_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBITL2_0_LC_4_9_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \POWERLED.func_state_RNIBITL2_0_LC_4_9_2  (
            .in0(N__16720),
            .in1(N__18258),
            .in2(N__16738),
            .in3(N__18456),
            .lcout(\POWERLED.N_96 ),
            .ltout(\POWERLED.N_96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_4_LC_4_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_4_LC_4_9_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_4_LC_4_9_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \POWERLED.count_off_4_LC_4_9_3  (
            .in0(N__20197),
            .in1(_gnd_net_),
            .in2(N__16735),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32885),
            .ce(N__20625),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI9QOB1_0_LC_4_9_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI9QOB1_0_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI9QOB1_0_LC_4_9_4 .LUT_INIT=16'b0000010000001000;
    LogicCell40 \POWERLED.func_state_RNI9QOB1_0_LC_4_9_4  (
            .in0(N__28817),
            .in1(N__16993),
            .in2(N__19905),
            .in3(N__22893),
            .lcout(\POWERLED.un1_count_off_0_sqmuxa_4_i_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2O4A1_0_0_LC_4_9_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2O4A1_0_0_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2O4A1_0_0_LC_4_9_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.func_state_RNI2O4A1_0_0_LC_4_9_5  (
            .in0(N__24812),
            .in1(N__19897),
            .in2(N__22897),
            .in3(N__28816),
            .lcout(),
            .ltout(\POWERLED.N_455_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIEB7T2_0_LC_4_9_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIEB7T2_0_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIEB7T2_0_LC_4_9_6 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \POWERLED.func_state_RNIEB7T2_0_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(N__32314),
            .in2(N__16714),
            .in3(N__22989),
            .lcout(),
            .ltout(\POWERLED.count_clk_en_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI81TV4_1_LC_4_9_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI81TV4_1_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI81TV4_1_LC_4_9_7 .LUT_INIT=16'b0010000000110000;
    LogicCell40 \POWERLED.func_state_RNI81TV4_1_LC_4_9_7  (
            .in0(N__31061),
            .in1(N__19759),
            .in2(N__16939),
            .in3(N__23038),
            .lcout(\POWERLED.func_state_RNI81TV4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_1_sqmuxa_i_i_o2_LC_4_10_0 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_i_i_o2_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_i_i_o2_LC_4_10_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \POWERLED.un1_count_clk_1_sqmuxa_i_i_o2_LC_4_10_0  (
            .in0(N__30475),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30376),
            .lcout(\POWERLED.N_239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_0_LC_4_10_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_0_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_0_LC_4_10_1 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \POWERLED.func_state_RNI5DLR_0_LC_4_10_1  (
            .in0(N__19889),
            .in1(N__22885),
            .in2(_gnd_net_),
            .in3(N__19749),
            .lcout(\POWERLED.N_480 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIAG3J3_1_LC_4_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIAG3J3_1_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIAG3J3_1_LC_4_10_2 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \POWERLED.func_state_RNIAG3J3_1_LC_4_10_2  (
            .in0(N__28844),
            .in1(N__17008),
            .in2(_gnd_net_),
            .in3(N__18420),
            .lcout(),
            .ltout(\POWERLED.func_state_1_ss0_i_0_o3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNILFRF4_0_LC_4_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNILFRF4_0_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNILFRF4_0_LC_4_10_3 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \POWERLED.func_state_RNILFRF4_0_LC_4_10_3  (
            .in0(N__25144),
            .in1(N__16795),
            .in2(N__16789),
            .in3(N__19828),
            .lcout(\POWERLED.func_state_RNILFRF4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNICP854_0_LC_4_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNICP854_0_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNICP854_0_LC_4_10_4 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \POWERLED.func_state_RNICP854_0_LC_4_10_4  (
            .in0(N__19750),
            .in1(N__16975),
            .in2(N__22896),
            .in3(N__19890),
            .lcout(\POWERLED.func_state_1_m0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI34G9_0_1_LC_4_10_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI34G9_0_1_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI34G9_0_1_LC_4_10_5 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \POWERLED.func_state_RNI34G9_0_1_LC_4_10_5  (
            .in0(N__31790),
            .in1(N__31860),
            .in2(_gnd_net_),
            .in3(N__28843),
            .lcout(\POWERLED.N_217 ),
            .ltout(\POWERLED.N_217_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIV0AS_1_LC_4_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIV0AS_1_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIV0AS_1_LC_4_10_6 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \POWERLED.func_state_RNIV0AS_1_LC_4_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16777),
            .in3(N__24995),
            .lcout(\POWERLED.N_487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_4_0_LC_4_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_4_0_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_4_0_LC_4_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_4_0_LC_4_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18234),
            .lcout(\POWERLED.N_2168_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI34G9_1_LC_4_11_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI34G9_1_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI34G9_1_LC_4_11_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \POWERLED.func_state_RNI34G9_1_LC_4_11_0  (
            .in0(N__31791),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28860),
            .lcout(\POWERLED.N_321 ),
            .ltout(\POWERLED.N_321_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNICU8L1_1_LC_4_11_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNICU8L1_1_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNICU8L1_1_LC_4_11_1 .LUT_INIT=16'b1010101110001011;
    LogicCell40 \POWERLED.func_state_RNICU8L1_1_LC_4_11_1  (
            .in0(N__16992),
            .in1(N__19888),
            .in2(N__17011),
            .in3(N__31894),
            .lcout(\POWERLED.func_state_1_ss0_i_0_o3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_EN_i_0_i_LC_4_11_4 .C_ON=1'b0;
    defparam \POWERLED.VCCST_EN_i_0_i_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_EN_i_0_i_LC_4_11_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.VCCST_EN_i_0_i_LC_4_11_4  (
            .in0(N__25146),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30451),
            .lcout(vccst_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_LC_4_11_5 .C_ON=1'b0;
    defparam \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_LC_4_11_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_LC_4_11_5  (
            .in0(N__30358),
            .in1(N__33945),
            .in2(N__31795),
            .in3(N__23374),
            .lcout(\POWERLED.N_516 ),
            .ltout(\POWERLED.N_516_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI7CJ93_1_LC_4_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI7CJ93_1_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI7CJ93_1_LC_4_11_6 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \POWERLED.func_state_RNI7CJ93_1_LC_4_11_6  (
            .in0(_gnd_net_),
            .in1(N__28861),
            .in2(N__16978),
            .in3(N__18419),
            .lcout(\POWERLED.N_403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_LC_4_12_0 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_0_c_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_LC_4_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17020),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(\COUNTER.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_LC_4_12_1 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_1_c_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_LC_4_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_1_c_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17326),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_0 ),
            .carryout(\COUNTER.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_LC_4_12_2 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_2_c_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_LC_4_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_2_c_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16969),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_1 ),
            .carryout(\COUNTER.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_LC_4_12_3 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_3_c_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_LC_4_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_3_c_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16954),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_2 ),
            .carryout(\COUNTER.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_LC_4_12_4 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_4_c_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_LC_4_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_4_c_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17125),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_3 ),
            .carryout(\COUNTER.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_LC_4_12_5 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_5_c_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_LC_4_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_5_c_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17110),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_4 ),
            .carryout(\COUNTER.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_LC_4_12_6 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_6_c_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_LC_4_12_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_6_c_LC_4_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17095),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_5 ),
            .carryout(\COUNTER.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_LC_4_12_7 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_7_c_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_LC_4_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_7_c_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17080),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_6 ),
            .carryout(COUNTER_un4_counter_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_13_0.C_ON=1'b0;
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_13_0.SEQ_MODE=4'b0000;
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_13_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_13_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17065),
            .lcout(COUNTER_un4_counter_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_LC_4_13_1 .C_ON=1'b0;
    defparam \COUNTER.counter_1_LC_4_13_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_1_LC_4_13_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_1_LC_4_13_1  (
            .in0(N__18501),
            .in1(N__17379),
            .in2(_gnd_net_),
            .in3(N__21724),
            .lcout(\COUNTER.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32972),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_5_LC_4_13_2 .C_ON=1'b0;
    defparam \COUNTER.counter_5_LC_4_13_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_5_LC_4_13_2 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \COUNTER.counter_5_LC_4_13_2  (
            .in0(N__17355),
            .in1(_gnd_net_),
            .in2(N__21747),
            .in3(N__17062),
            .lcout(\COUNTER.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32972),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_3_LC_4_13_3 .C_ON=1'b0;
    defparam \COUNTER.counter_3_LC_4_13_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_3_LC_4_13_3 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \COUNTER.counter_3_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__17053),
            .in2(N__17040),
            .in3(N__21722),
            .lcout(\COUNTER.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32972),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_RNO_LC_4_13_4 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_4_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_RNO_LC_4_13_4  (
            .in0(N__17300),
            .in1(N__17033),
            .in2(N__18591),
            .in3(N__18500),
            .lcout(\COUNTER.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_RNO_LC_4_13_5 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_4_13_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \COUNTER.un4_counter_1_c_RNO_LC_4_13_5  (
            .in0(N__17375),
            .in1(N__17354),
            .in2(N__17277),
            .in3(N__17341),
            .lcout(\COUNTER.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_4_LC_4_13_6 .C_ON=1'b0;
    defparam \COUNTER.counter_4_LC_4_13_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_4_LC_4_13_6 .LUT_INIT=16'b0001010000010100;
    LogicCell40 \COUNTER.counter_4_LC_4_13_6  (
            .in0(N__21718),
            .in1(N__17317),
            .in2(N__17307),
            .in3(_gnd_net_),
            .lcout(\COUNTER.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32972),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_6_LC_4_13_7 .C_ON=1'b0;
    defparam \COUNTER.counter_6_LC_4_13_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_6_LC_4_13_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_6_LC_4_13_7  (
            .in0(N__17287),
            .in1(N__17276),
            .in2(_gnd_net_),
            .in3(N__21723),
            .lcout(\COUNTER.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32972),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_0_LC_4_14_0 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_0_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_0_LC_4_14_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_0_LC_4_14_0  (
            .in0(N__27571),
            .in1(N__17226),
            .in2(N__17254),
            .in3(N__17253),
            .lcout(\DSW_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\DSW_PWRGD.un1_count_1_cry_0 ),
            .clk(N__33058),
            .ce(),
            .sr(N__17574));
    defparam \DSW_PWRGD.count_1_LC_4_14_1 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_1_LC_4_14_1 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_1_LC_4_14_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_1_LC_4_14_1  (
            .in0(N__27567),
            .in1(N__17208),
            .in2(_gnd_net_),
            .in3(N__17194),
            .lcout(\DSW_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_0 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_1 ),
            .clk(N__33058),
            .ce(),
            .sr(N__17574));
    defparam \DSW_PWRGD.count_2_LC_4_14_2 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_2_LC_4_14_2 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_2_LC_4_14_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_2_LC_4_14_2  (
            .in0(N__27572),
            .in1(N__17190),
            .in2(_gnd_net_),
            .in3(N__17176),
            .lcout(\DSW_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_1 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_2 ),
            .clk(N__33058),
            .ce(),
            .sr(N__17574));
    defparam \DSW_PWRGD.count_3_LC_4_14_3 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_3_LC_4_14_3 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_3_LC_4_14_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_3_LC_4_14_3  (
            .in0(N__27568),
            .in1(N__17166),
            .in2(_gnd_net_),
            .in3(N__17152),
            .lcout(\DSW_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_2 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_3 ),
            .clk(N__33058),
            .ce(),
            .sr(N__17574));
    defparam \DSW_PWRGD.count_4_LC_4_14_4 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_4_LC_4_14_4 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_4_LC_4_14_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_4_LC_4_14_4  (
            .in0(N__27573),
            .in1(N__17142),
            .in2(_gnd_net_),
            .in3(N__17128),
            .lcout(\DSW_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_3 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_4 ),
            .clk(N__33058),
            .ce(),
            .sr(N__17574));
    defparam \DSW_PWRGD.count_5_LC_4_14_5 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_5_LC_4_14_5 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_5_LC_4_14_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_5_LC_4_14_5  (
            .in0(N__27569),
            .in1(N__17532),
            .in2(_gnd_net_),
            .in3(N__17518),
            .lcout(\DSW_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_4 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_5 ),
            .clk(N__33058),
            .ce(),
            .sr(N__17574));
    defparam \DSW_PWRGD.count_6_LC_4_14_6 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_6_LC_4_14_6 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_6_LC_4_14_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_6_LC_4_14_6  (
            .in0(N__27574),
            .in1(N__17514),
            .in2(_gnd_net_),
            .in3(N__17500),
            .lcout(\DSW_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_5 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_6 ),
            .clk(N__33058),
            .ce(),
            .sr(N__17574));
    defparam \DSW_PWRGD.count_7_LC_4_14_7 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_7_LC_4_14_7 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_7_LC_4_14_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_7_LC_4_14_7  (
            .in0(N__27570),
            .in1(N__17496),
            .in2(_gnd_net_),
            .in3(N__17479),
            .lcout(\DSW_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_6 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_7 ),
            .clk(N__33058),
            .ce(),
            .sr(N__17574));
    defparam \DSW_PWRGD.count_8_LC_4_15_0 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_8_LC_4_15_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_8_LC_4_15_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_8_LC_4_15_0  (
            .in0(N__27566),
            .in1(N__17475),
            .in2(_gnd_net_),
            .in3(N__17461),
            .lcout(\DSW_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_4_15_0_),
            .carryout(\DSW_PWRGD.un1_count_1_cry_8 ),
            .clk(N__32974),
            .ce(),
            .sr(N__17567));
    defparam \DSW_PWRGD.count_9_LC_4_15_1 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_9_LC_4_15_1 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_9_LC_4_15_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_9_LC_4_15_1  (
            .in0(N__27558),
            .in1(N__17457),
            .in2(_gnd_net_),
            .in3(N__17440),
            .lcout(\DSW_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_8 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_9 ),
            .clk(N__32974),
            .ce(),
            .sr(N__17567));
    defparam \DSW_PWRGD.count_10_LC_4_15_2 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_10_LC_4_15_2 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_10_LC_4_15_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_10_LC_4_15_2  (
            .in0(N__27563),
            .in1(N__17436),
            .in2(_gnd_net_),
            .in3(N__17422),
            .lcout(\DSW_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_9 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_10 ),
            .clk(N__32974),
            .ce(),
            .sr(N__17567));
    defparam \DSW_PWRGD.count_11_LC_4_15_3 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_11_LC_4_15_3 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_11_LC_4_15_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_11_LC_4_15_3  (
            .in0(N__27556),
            .in1(N__17418),
            .in2(_gnd_net_),
            .in3(N__17404),
            .lcout(\DSW_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_10 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_11 ),
            .clk(N__32974),
            .ce(),
            .sr(N__17567));
    defparam \DSW_PWRGD.count_12_LC_4_15_4 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_12_LC_4_15_4 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_12_LC_4_15_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_12_LC_4_15_4  (
            .in0(N__27564),
            .in1(N__17397),
            .in2(_gnd_net_),
            .in3(N__17383),
            .lcout(\DSW_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_11 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_12 ),
            .clk(N__32974),
            .ce(),
            .sr(N__17567));
    defparam \DSW_PWRGD.count_13_LC_4_15_5 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_13_LC_4_15_5 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_13_LC_4_15_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_13_LC_4_15_5  (
            .in0(N__27557),
            .in1(N__17646),
            .in2(_gnd_net_),
            .in3(N__17632),
            .lcout(\DSW_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_12 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_13 ),
            .clk(N__32974),
            .ce(),
            .sr(N__17567));
    defparam \DSW_PWRGD.count_14_LC_4_15_6 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_14_LC_4_15_6 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_14_LC_4_15_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_14_LC_4_15_6  (
            .in0(N__27565),
            .in1(N__17628),
            .in2(_gnd_net_),
            .in3(N__17611),
            .lcout(\DSW_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_13 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_14 ),
            .clk(N__32974),
            .ce(),
            .sr(N__17567));
    defparam \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_4_15_7 .C_ON=1'b1;
    defparam \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_4_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(N__27254),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_14 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_esr_15_LC_4_16_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_esr_15_LC_4_16_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_esr_15_LC_4_16_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DSW_PWRGD.count_esr_15_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__17601),
            .in2(_gnd_net_),
            .in3(N__17608),
            .lcout(\DSW_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33059),
            .ce(N__17587),
            .sr(N__17575));
    defparam \POWERLED.count_RNI_2_LC_5_1_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_2_LC_5_1_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_2_LC_5_1_0 .LUT_INIT=16'b0000000100000001;
    LogicCell40 \POWERLED.count_RNI_2_LC_5_1_0  (
            .in0(N__19076),
            .in1(N__19043),
            .in2(N__19012),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlt6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_5_LC_5_1_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_5_LC_5_1_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_5_LC_5_1_1 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \POWERLED.count_RNI_5_LC_5_1_1  (
            .in0(N__18914),
            .in1(N__18888),
            .in2(N__17548),
            .in3(N__18960),
            .lcout(\POWERLED.un79_clk_100khzlto15_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_10_LC_5_1_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_10_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_10_LC_5_1_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_RNI_10_LC_5_1_2  (
            .in0(N__19188),
            .in1(N__19261),
            .in2(N__19224),
            .in3(N__19286),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlto15_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_15_LC_5_1_3 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_15_LC_5_1_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_15_LC_5_1_3 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \POWERLED.count_RNI_15_LC_5_1_3  (
            .in0(N__19155),
            .in1(_gnd_net_),
            .in2(N__17545),
            .in3(N__19118),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlto15_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_8_LC_5_1_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_8_LC_5_1_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_8_LC_5_1_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.count_RNI_8_LC_5_1_4  (
            .in0(N__19313),
            .in1(N__18851),
            .in2(N__17542),
            .in3(N__17539),
            .lcout(\POWERLED.count_RNIZ0Z_8 ),
            .ltout(\POWERLED.count_RNIZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_0_LC_5_1_5 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_0_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_0_LC_5_1_5 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \POWERLED.pwm_out_RNO_0_LC_5_1_5  (
            .in0(_gnd_net_),
            .in1(N__33998),
            .in2(N__17731),
            .in3(N__22381),
            .lcout(\POWERLED.pwm_out_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNIFPNR_0_LC_5_1_6 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNIFPNR_0_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNIFPNR_0_LC_5_1_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.curr_state_RNIFPNR_0_LC_5_1_6  (
            .in0(N__22380),
            .in1(N__32317),
            .in2(N__34020),
            .in3(N__22353),
            .lcout(\POWERLED.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_LC_5_2_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_LC_5_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_LC_5_2_0  (
            .in0(_gnd_net_),
            .in1(N__18702),
            .in2(N__18750),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_2_0_),
            .carryout(\POWERLED.un1_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_5_2_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_5_2_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_RNIB209_LC_5_2_1  (
            .in0(N__17790),
            .in1(N__19077),
            .in2(_gnd_net_),
            .in3(N__17713),
            .lcout(\POWERLED.un1_count_cry_1_c_RNIBZ0Z209 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_1 ),
            .carryout(\POWERLED.un1_count_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_2_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_2_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_2_2  (
            .in0(N__17793),
            .in1(N__19050),
            .in2(_gnd_net_),
            .in3(N__17698),
            .lcout(\POWERLED.un1_count_cry_2_c_RNICZ0Z419 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_2 ),
            .carryout(\POWERLED.un1_count_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_5_2_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_5_2_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_3_c_RNID629_LC_5_2_3  (
            .in0(N__17789),
            .in1(N__19010),
            .in2(_gnd_net_),
            .in3(N__17680),
            .lcout(\POWERLED.un1_count_cry_3_c_RNIDZ0Z629 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_3 ),
            .carryout(\POWERLED.un1_count_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_2_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_2_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_2_4  (
            .in0(N__17795),
            .in1(N__18959),
            .in2(_gnd_net_),
            .in3(N__17662),
            .lcout(\POWERLED.un1_count_cry_4_c_RNIEZ0Z839 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_4 ),
            .carryout(\POWERLED.un1_count_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_5_2_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_5_2_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_5_c_RNIFA49_LC_5_2_5  (
            .in0(N__17791),
            .in1(N__18918),
            .in2(_gnd_net_),
            .in3(N__17659),
            .lcout(\POWERLED.un1_count_cry_5_c_RNIFAZ0Z49 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_5 ),
            .carryout(\POWERLED.un1_count_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_5_2_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_5_2_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_6_c_RNIGC59_LC_5_2_6  (
            .in0(N__17794),
            .in1(N__18887),
            .in2(_gnd_net_),
            .in3(N__17656),
            .lcout(\POWERLED.un1_count_cry_6_c_RNIGCZ0Z59 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_6 ),
            .carryout(\POWERLED.un1_count_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_5_2_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_5_2_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_5_2_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_7_c_RNIHE69_LC_5_2_7  (
            .in0(N__17792),
            .in1(N__18852),
            .in2(_gnd_net_),
            .in3(N__17866),
            .lcout(\POWERLED.un1_count_cry_7_c_RNIHEZ0Z69 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_7 ),
            .carryout(\POWERLED.un1_count_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_5_3_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_5_3_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_8_c_RNIIG79_LC_5_3_0  (
            .in0(N__17817),
            .in1(N__19317),
            .in2(_gnd_net_),
            .in3(N__17863),
            .lcout(\POWERLED.un1_count_cry_8_c_RNIIGZ0Z79 ),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(\POWERLED.un1_count_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_5_3_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_5_3_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_9_c_RNIJI89_LC_5_3_1  (
            .in0(N__17821),
            .in1(N__19287),
            .in2(_gnd_net_),
            .in3(N__17860),
            .lcout(\POWERLED.un1_count_cry_9_c_RNIJIZ0Z89 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_9 ),
            .carryout(\POWERLED.un1_count_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_5_3_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_5_3_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_5_3_2  (
            .in0(N__17818),
            .in1(N__19259),
            .in2(_gnd_net_),
            .in3(N__17857),
            .lcout(\POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_10 ),
            .carryout(\POWERLED.un1_count_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_5_3_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_5_3_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_11_c_RNISEH7_LC_5_3_3  (
            .in0(N__17820),
            .in1(N__19220),
            .in2(_gnd_net_),
            .in3(N__17845),
            .lcout(\POWERLED.un1_count_cry_11_c_RNISEHZ0Z7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_11 ),
            .carryout(\POWERLED.un1_count_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_5_3_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_5_3_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_12_c_RNITGI7_LC_5_3_4  (
            .in0(N__17819),
            .in1(N__19181),
            .in2(_gnd_net_),
            .in3(N__17830),
            .lcout(\POWERLED.un1_count_cry_12_c_RNITGIZ0Z7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_12 ),
            .carryout(\POWERLED.un1_count_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_5_3_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_5_3_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_5_3_5  (
            .in0(N__17822),
            .in1(N__19148),
            .in2(_gnd_net_),
            .in3(N__17827),
            .lcout(\POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_13 ),
            .carryout(\POWERLED.un1_count_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_5_3_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_5_3_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_5_3_6  (
            .in0(N__19126),
            .in1(N__17823),
            .in2(_gnd_net_),
            .in3(N__17752),
            .lcout(\POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_14_LC_5_3_7 .C_ON=1'b0;
    defparam \POWERLED.count_14_LC_5_3_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_14_LC_5_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_14_LC_5_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17748),
            .lcout(\POWERLED.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32659),
            .ce(N__32286),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_4_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18091),
            .lcout(\POWERLED.un85_clk_100khz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_4_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_4_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17920),
            .lcout(\POWERLED.un85_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_4_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_4_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17997),
            .lcout(\POWERLED.un85_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_4_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_4_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18343),
            .lcout(\POWERLED.un85_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_4_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_4_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18307),
            .lcout(\POWERLED.un85_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_PWRGD_LC_5_4_7 .C_ON=1'b0;
    defparam \POWERLED.VCCST_PWRGD_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_PWRGD_LC_5_4_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.VCCST_PWRGD_LC_5_4_7  (
            .in0(_gnd_net_),
            .in1(N__27787),
            .in2(_gnd_net_),
            .in3(N__20784),
            .lcout(vccst_pwrgd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_5_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_5_0  (
            .in0(_gnd_net_),
            .in1(N__21282),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_5_0_),
            .carryout(\POWERLED.mult1_un145_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_5_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(N__19363),
            .in2(N__17970),
            .in3(N__17881),
            .lcout(\POWERLED.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_5_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(N__17966),
            .in2(N__17878),
            .in3(N__17869),
            .lcout(\POWERLED.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_5_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(N__17992),
            .in2(N__18040),
            .in3(N__18031),
            .lcout(\POWERLED.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_5_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(N__18028),
            .in2(N__17998),
            .in3(N__18022),
            .lcout(\POWERLED.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_5_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_5_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_5_5  (
            .in0(N__18306),
            .in1(N__18019),
            .in2(N__17971),
            .in3(N__18013),
            .lcout(\POWERLED.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_5_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_5_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18010),
            .in3(N__18001),
            .lcout(\POWERLED.mult1_un145_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_5_5_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_5_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_5_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17991),
            .lcout(\POWERLED.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_5_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_5_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(N__21469),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_6_0_),
            .carryout(\POWERLED.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_5_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_5_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_5_6_1  (
            .in0(_gnd_net_),
            .in1(N__19357),
            .in2(N__19390),
            .in3(N__17944),
            .lcout(\POWERLED.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_5_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_5_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__19515),
            .in2(N__19501),
            .in3(N__17935),
            .lcout(\POWERLED.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_5_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_5_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(N__19417),
            .in2(N__19330),
            .in3(N__17923),
            .lcout(\POWERLED.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_5_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_5_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_5_6_4  (
            .in0(_gnd_net_),
            .in1(N__19570),
            .in2(N__19423),
            .in3(N__18109),
            .lcout(\POWERLED.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_5_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_5_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_5_6_5  (
            .in0(N__18082),
            .in1(N__19560),
            .in2(N__18058),
            .in3(N__18097),
            .lcout(\POWERLED.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_5_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_5_6_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_5_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19531),
            .in3(N__18094),
            .lcout(\POWERLED.mult1_un124_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_5_6_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_5_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(N__19561),
            .in2(_gnd_net_),
            .in3(N__19416),
            .lcout(\POWERLED.mult1_un124_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_5_7_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_5_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21286),
            .lcout(\POWERLED.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_5_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_5_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(N__31547),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(\POWERLED.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_5_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_5_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__21517),
            .in2(N__18201),
            .in3(N__18049),
            .lcout(\POWERLED.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_5_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_5_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_5_8_2  (
            .in0(_gnd_net_),
            .in1(N__18197),
            .in2(N__18175),
            .in3(N__18046),
            .lcout(\POWERLED.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_5_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_5_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_5_8_3  (
            .in0(_gnd_net_),
            .in1(N__18334),
            .in2(N__18151),
            .in3(N__18043),
            .lcout(\POWERLED.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_5_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_5_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_5_8_4  (
            .in0(_gnd_net_),
            .in1(N__18124),
            .in2(N__18342),
            .in3(N__18211),
            .lcout(\POWERLED.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_5_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_5_8_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_5_8_5  (
            .in0(N__19610),
            .in1(N__18385),
            .in2(N__18202),
            .in3(N__18208),
            .lcout(\POWERLED.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_5_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_5_8_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_5_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18367),
            .in3(N__18205),
            .lcout(\POWERLED.mult1_un159_sum_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_5_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_5_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_5_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18333),
            .lcout(\POWERLED.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_2_LC_5_9_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_5_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_2_LC_5_9_0  (
            .in0(_gnd_net_),
            .in1(N__26414),
            .in2(_gnd_net_),
            .in3(N__29338),
            .lcout(\POWERLED.N_505 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\POWERLED.mult1_un152_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_5_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_5_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(N__18184),
            .in2(N__18282),
            .in3(N__18166),
            .lcout(\POWERLED.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_5_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_5_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__18278),
            .in2(N__18163),
            .in3(N__18142),
            .lcout(\POWERLED.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_5_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_5_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(N__18309),
            .in2(N__18139),
            .in3(N__18118),
            .lcout(\POWERLED.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_5_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_5_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(N__18394),
            .in2(N__18313),
            .in3(N__18379),
            .lcout(\POWERLED.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_5_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_5_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_5_9_5  (
            .in0(N__18338),
            .in1(N__18376),
            .in2(N__18283),
            .in3(N__18358),
            .lcout(\POWERLED.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_5_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_5_9_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(N__18355),
            .in2(_gnd_net_),
            .in3(N__18346),
            .lcout(\POWERLED.mult1_un152_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18308),
            .lcout(\POWERLED.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_0_LC_5_10_0 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_0_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_0_LC_5_10_0 .LUT_INIT=16'b0010000010000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_0_LC_5_10_0  (
            .in0(N__19720),
            .in1(N__22862),
            .in2(N__18265),
            .in3(N__28851),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_o_N_423_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_2_LC_5_10_1 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_2_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_2_LC_5_10_1 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_2_LC_5_10_1  (
            .in0(N__31080),
            .in1(N__24724),
            .in2(N__18238),
            .in3(N__23059),
            .lcout(\POWERLED.un1_func_state25_6_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_LC_5_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_LC_5_10_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.func_state_RNI_0_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__19886),
            .in2(_gnd_net_),
            .in3(N__22861),
            .lcout(\POWERLED.N_348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_0_0_LC_5_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_0_0_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_0_0_LC_5_10_3 .LUT_INIT=16'b0100100000000000;
    LogicCell40 \POWERLED.func_state_RNI5DLR_0_0_LC_5_10_3  (
            .in0(N__30532),
            .in1(N__24723),
            .in2(N__30384),
            .in3(N__23058),
            .lcout(\POWERLED.func_state_RNI5DLR_0Z0Z_0 ),
            .ltout(\POWERLED.func_state_RNI5DLR_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIIBB64_0_LC_5_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIIBB64_0_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIIBB64_0_LC_5_10_4 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \POWERLED.func_state_RNIIBB64_0_LC_5_10_4  (
            .in0(N__18220),
            .in1(N__19887),
            .in2(N__18214),
            .in3(N__25125),
            .lcout(),
            .ltout(\POWERLED.func_state_1_m0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIU8CJB_0_LC_5_10_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIU8CJB_0_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIU8CJB_0_LC_5_10_5 .LUT_INIT=16'b0000000001110010;
    LogicCell40 \POWERLED.func_state_RNIU8CJB_0_LC_5_10_5  (
            .in0(N__21778),
            .in1(N__19806),
            .in2(N__18463),
            .in3(N__23338),
            .lcout(\POWERLED.func_state_RNIU8CJBZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_S4n_RNI5DLR_0_LC_5_10_6.C_ON=1'b0;
    defparam SLP_S4n_RNI5DLR_0_LC_5_10_6.SEQ_MODE=4'b0000;
    defparam SLP_S4n_RNI5DLR_0_LC_5_10_6.LUT_INIT=16'b0000000001000000;
    LogicCell40 SLP_S4n_RNI5DLR_0_LC_5_10_6 (
            .in0(N__30354),
            .in1(N__30533),
            .in2(N__31893),
            .in3(N__28850),
            .lcout(m3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_2_LC_5_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_2_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_2_LC_5_10_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_2_LC_5_10_7  (
            .in0(N__24814),
            .in1(N__31875),
            .in2(N__28864),
            .in3(N__18460),
            .lcout(\POWERLED.un1_func_state25_6_0_o_N_425_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_10_LC_5_11_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_10_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_10_LC_5_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_10_LC_5_11_0  (
            .in0(N__20281),
            .in1(N__20097),
            .in2(N__20067),
            .in3(N__20457),
            .lcout(),
            .ltout(\POWERLED.un34_clk_100khz_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_0_10_LC_5_11_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_0_10_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_0_10_LC_5_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.count_off_RNI_0_10_LC_5_11_1  (
            .in0(N__18433),
            .in1(N__18400),
            .in2(N__18436),
            .in3(N__18472),
            .lcout(\POWERLED.count_off_RNI_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIBITL2_0_LC_5_11_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIBITL2_0_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIBITL2_0_LC_5_11_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.count_off_RNIBITL2_0_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__20332),
            .in2(_gnd_net_),
            .in3(N__20013),
            .lcout(\POWERLED.count_off_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_3_LC_5_11_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_3_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_3_LC_5_11_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_3_LC_5_11_4  (
            .in0(N__20677),
            .in1(N__20217),
            .in2(N__19942),
            .in3(N__20236),
            .lcout(\POWERLED.un34_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_1_sqmuxa_i_i_o3_LC_5_11_5 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_i_i_o3_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_i_i_o3_LC_5_11_5 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \POWERLED.un1_count_clk_1_sqmuxa_i_i_o3_LC_5_11_5  (
            .in0(N__30527),
            .in1(N__24405),
            .in2(N__30380),
            .in3(N__33933),
            .lcout(\POWERLED.N_322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_0_1_LC_5_11_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_0_1_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_0_1_LC_5_11_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.count_off_RNI_0_1_LC_5_11_7  (
            .in0(N__19966),
            .in1(N__19990),
            .in2(N__20146),
            .in3(N__20179),
            .lcout(\POWERLED.un34_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIDVQT9_3_LC_5_12_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIDVQT9_3_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIDVQT9_3_LC_5_12_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \POWERLED.count_off_RNIDVQT9_3_LC_5_12_0  (
            .in0(N__20348),
            .in1(N__19926),
            .in2(N__18544),
            .in3(N__20587),
            .lcout(\POWERLED.count_offZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_3_LC_5_12_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_3_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_3_LC_5_12_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \POWERLED.count_off_3_LC_5_12_1  (
            .in0(N__19927),
            .in1(N__20351),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33045),
            .ce(N__20610),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_1_LC_5_12_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_1_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_1_LC_5_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_off_1_LC_5_12_2  (
            .in0(N__20349),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18487),
            .lcout(\POWERLED.count_off_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33045),
            .ce(N__20610),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIIIPE9_0_LC_5_12_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIIIPE9_0_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIIIPE9_0_LC_5_12_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIIIPE9_0_LC_5_12_6  (
            .in0(N__18526),
            .in1(N__18535),
            .in2(_gnd_net_),
            .in3(N__20586),
            .lcout(\POWERLED.count_offZ0Z_0 ),
            .ltout(\POWERLED.count_offZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_0_LC_5_12_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_0_LC_5_12_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_0_LC_5_12_7 .LUT_INIT=16'b0000110000001100;
    LogicCell40 \POWERLED.count_off_0_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__20350),
            .in2(N__18529),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33045),
            .ce(N__20610),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_0_LC_5_13_0 .C_ON=1'b0;
    defparam \COUNTER.counter_0_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_0_LC_5_13_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \COUNTER.counter_0_LC_5_13_0  (
            .in0(N__21725),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18520),
            .lcout(\COUNTER.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32971),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_1_LC_5_13_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_1_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_1_LC_5_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.count_off_RNI_1_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(N__19985),
            .in2(_gnd_net_),
            .in3(N__20012),
            .lcout(\POWERLED.count_off_RNIZ0Z_1 ),
            .ltout(\POWERLED.count_off_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIJJPE9_1_LC_5_13_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIJJPE9_1_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIJJPE9_1_LC_5_13_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \POWERLED.count_off_RNIJJPE9_1_LC_5_13_3  (
            .in0(N__18481),
            .in1(N__20364),
            .in2(N__18475),
            .in3(N__20588),
            .lcout(\POWERLED.count_offZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_15_LC_5_13_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_15_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_15_LC_5_13_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_15_LC_5_13_4  (
            .in0(N__20406),
            .in1(N__20430),
            .in2(N__20017),
            .in3(N__20262),
            .lcout(\POWERLED.un34_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_2_LC_5_13_5 .C_ON=1'b0;
    defparam \COUNTER.counter_2_LC_5_13_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_2_LC_5_13_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \COUNTER.counter_2_LC_5_13_5  (
            .in0(N__18604),
            .in1(N__21726),
            .in2(_gnd_net_),
            .in3(N__18590),
            .lcout(\COUNTER.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32971),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_5_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_5_13_6 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_5_13_6  (
            .in0(N__30469),
            .in1(N__30295),
            .in2(_gnd_net_),
            .in3(N__25143),
            .lcout(\POWERLED.N_292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIF9MQ9_13_LC_5_14_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIF9MQ9_13_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIF9MQ9_13_LC_5_14_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_off_RNIF9MQ9_13_LC_5_14_0  (
            .in0(N__20419),
            .in1(N__18568),
            .in2(_gnd_net_),
            .in3(N__20595),
            .lcout(\POWERLED.count_offZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_13_LC_5_14_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_13_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_13_LC_5_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_13_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20418),
            .lcout(\POWERLED.count_off_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33042),
            .ce(N__20626),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIH5TT9_5_LC_5_14_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIH5TT9_5_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIH5TT9_5_LC_5_14_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIH5TT9_5_LC_5_14_2  (
            .in0(N__18562),
            .in1(N__20160),
            .in2(_gnd_net_),
            .in3(N__20593),
            .lcout(\POWERLED.count_offZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_5_LC_5_14_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_5_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_5_LC_5_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_5_LC_5_14_3  (
            .in0(N__20161),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33042),
            .ce(N__20626),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIHCNQ9_14_LC_5_14_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIHCNQ9_14_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIHCNQ9_14_LC_5_14_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \POWERLED.count_off_RNIHCNQ9_14_LC_5_14_4  (
            .in0(N__20395),
            .in1(N__20596),
            .in2(_gnd_net_),
            .in3(N__18556),
            .lcout(\POWERLED.count_offZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_14_LC_5_14_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_14_LC_5_14_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_14_LC_5_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_14_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20394),
            .lcout(\POWERLED.count_off_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33042),
            .ce(N__20626),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIJ8UT9_6_LC_5_14_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIJ8UT9_6_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIJ8UT9_6_LC_5_14_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIJ8UT9_6_LC_5_14_6  (
            .in0(N__18550),
            .in1(N__20124),
            .in2(_gnd_net_),
            .in3(N__20594),
            .lcout(\POWERLED.count_offZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_6_LC_5_14_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_6_LC_5_14_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_6_LC_5_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_6_LC_5_14_7  (
            .in0(N__20125),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33042),
            .ce(N__20626),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI4RJN_6_LC_6_1_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI4RJN_6_LC_6_1_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI4RJN_6_LC_6_1_0 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \POWERLED.count_RNI4RJN_6_LC_6_1_0  (
            .in0(N__18667),
            .in1(N__33987),
            .in2(N__18679),
            .in3(_gnd_net_),
            .lcout(\POWERLED.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_6_LC_6_1_1 .C_ON=1'b0;
    defparam \POWERLED.count_6_LC_6_1_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_6_LC_6_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_6_LC_6_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18678),
            .lcout(\POWERLED.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32368),
            .ce(N__32284),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI4S8O_15_LC_6_1_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNI4S8O_15_LC_6_1_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI4S8O_15_LC_6_1_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI4S8O_15_LC_6_1_2  (
            .in0(N__18646),
            .in1(N__33986),
            .in2(_gnd_net_),
            .in3(N__18657),
            .lcout(\POWERLED.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_15_LC_6_1_3 .C_ON=1'b0;
    defparam \POWERLED.count_15_LC_6_1_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_15_LC_6_1_3 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_15_LC_6_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18661),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32368),
            .ce(N__32284),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI6UKN_7_LC_6_1_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI6UKN_7_LC_6_1_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI6UKN_7_LC_6_1_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI6UKN_7_LC_6_1_4  (
            .in0(N__18628),
            .in1(N__33988),
            .in2(_gnd_net_),
            .in3(N__18636),
            .lcout(\POWERLED.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_7_LC_6_1_5 .C_ON=1'b0;
    defparam \POWERLED.count_7_LC_6_1_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_7_LC_6_1_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_7_LC_6_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18640),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32368),
            .ce(N__32284),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI81MN_8_LC_6_1_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNI81MN_8_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI81MN_8_LC_6_1_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI81MN_8_LC_6_1_6  (
            .in0(N__18610),
            .in1(N__33989),
            .in2(_gnd_net_),
            .in3(N__18618),
            .lcout(\POWERLED.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_8_LC_6_1_7 .C_ON=1'b0;
    defparam \POWERLED.count_8_LC_6_1_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_8_LC_6_1_7 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_8_LC_6_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18622),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32368),
            .ce(N__32284),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIA4NN_9_LC_6_2_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNIA4NN_9_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIA4NN_9_LC_6_2_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNIA4NN_9_LC_6_2_0  (
            .in0(N__34001),
            .in1(N__18814),
            .in2(_gnd_net_),
            .in3(N__18822),
            .lcout(\POWERLED.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_9_LC_6_2_1 .C_ON=1'b0;
    defparam \POWERLED.count_9_LC_6_2_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_9_LC_6_2_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_9_LC_6_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18826),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32535),
            .ce(N__32287),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIJKSP_10_LC_6_2_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNIJKSP_10_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIJKSP_10_LC_6_2_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \POWERLED.count_RNIJKSP_10_LC_6_2_2  (
            .in0(N__34002),
            .in1(N__18808),
            .in2(_gnd_net_),
            .in3(N__18796),
            .lcout(\POWERLED.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_10_LC_6_2_3 .C_ON=1'b0;
    defparam \POWERLED.count_10_LC_6_2_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_10_LC_6_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_10_LC_6_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18807),
            .lcout(\POWERLED.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32535),
            .ce(N__32287),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNISEFN_2_LC_6_2_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNISEFN_2_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNISEFN_2_LC_6_2_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \POWERLED.count_RNISEFN_2_LC_6_2_4  (
            .in0(_gnd_net_),
            .in1(N__34000),
            .in2(N__18790),
            .in3(N__18778),
            .lcout(\POWERLED.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_2_LC_6_2_5 .C_ON=1'b0;
    defparam \POWERLED.count_2_LC_6_2_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_2_LC_6_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_2_LC_6_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18789),
            .lcout(\POWERLED.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32535),
            .ce(N__32287),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNISF4O_11_LC_6_2_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNISF4O_11_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNISF4O_11_LC_6_2_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \POWERLED.count_RNISF4O_11_LC_6_2_6  (
            .in0(N__34003),
            .in1(N__18772),
            .in2(_gnd_net_),
            .in3(N__18760),
            .lcout(\POWERLED.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_11_LC_6_2_7 .C_ON=1'b0;
    defparam \POWERLED.count_11_LC_6_2_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_11_LC_6_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_11_LC_6_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18771),
            .lcout(\POWERLED.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32535),
            .ce(N__32287),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_6_3_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_6_3_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_6_3_0  (
            .in0(N__18754),
            .in1(N__18715),
            .in2(N__19627),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_cry_0_i ),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_6_3_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_6_3_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_6_3_1  (
            .in0(N__18709),
            .in1(N__18685),
            .in2(N__19585),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4698_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_0 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_6_3_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_6_3_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_6_3_2  (
            .in0(_gnd_net_),
            .in1(N__19060),
            .in2(N__19087),
            .in3(N__19078),
            .lcout(\POWERLED.N_4699_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_1 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_6_3_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_6_3_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_6_3_3  (
            .in0(N__19054),
            .in1(N__19027),
            .in2(N__19021),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4700_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_2 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_6_3_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_6_3_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_6_3_4  (
            .in0(N__19011),
            .in1(N__18985),
            .in2(N__18979),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4701_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_3 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_6_3_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_6_3_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_6_3_5  (
            .in0(_gnd_net_),
            .in1(N__18970),
            .in2(N__18937),
            .in3(N__18964),
            .lcout(\POWERLED.N_4702_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_4 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_6_3_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_6_3_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_6_3_6  (
            .in0(_gnd_net_),
            .in1(N__18898),
            .in2(N__18928),
            .in3(N__18919),
            .lcout(\POWERLED.N_4703_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_5 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_6_3_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_6_3_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_6_3_7  (
            .in0(_gnd_net_),
            .in1(N__19381),
            .in2(N__18868),
            .in3(N__18892),
            .lcout(\POWERLED.N_4704_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_6 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_6_4_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_6_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_6_4_0  (
            .in0(_gnd_net_),
            .in1(N__21223),
            .in2(N__18835),
            .in3(N__18859),
            .lcout(\POWERLED.N_4705_i ),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_6_4_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_6_4_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_6_4_1  (
            .in0(N__19318),
            .in1(N__21229),
            .in2(N__19297),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4706_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_8 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_6_4_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_6_4_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_6_4_2  (
            .in0(N__19288),
            .in1(N__19267),
            .in2(N__20473),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4707_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_9 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_6_4_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_6_4_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_6_4_3  (
            .in0(N__19260),
            .in1(N__20482),
            .in2(N__19237),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_4708_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_10 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_6_4_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_6_4_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_6_4_4  (
            .in0(_gnd_net_),
            .in1(N__21292),
            .in2(N__19201),
            .in3(N__19228),
            .lcout(\POWERLED.N_4709_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_11 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_6_4_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_6_4_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_6_4_5  (
            .in0(_gnd_net_),
            .in1(N__19165),
            .in2(N__20707),
            .in3(N__19192),
            .lcout(\POWERLED.N_4710_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_12 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_6_4_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_6_4_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_6_4_6  (
            .in0(_gnd_net_),
            .in1(N__20716),
            .in2(N__19135),
            .in3(N__19159),
            .lcout(\POWERLED.N_4711_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_13 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_6_4_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_6_4_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_6_4_7  (
            .in0(_gnd_net_),
            .in1(N__23962),
            .in2(N__19102),
            .in3(N__19125),
            .lcout(\POWERLED.N_4712_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_14 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_6_5_0 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_6_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19090),
            .lcout(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_5_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_5_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_5_1  (
            .in0(N__19422),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_5_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_5_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21246),
            .lcout(\POWERLED.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_5_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21267),
            .lcout(\POWERLED.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_5_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_5_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21448),
            .lcout(\POWERLED.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_6_5_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_6_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_6_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21432),
            .lcout(\POWERLED.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_5_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_5_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21468),
            .lcout(\POWERLED.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_6_5_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_6_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_6_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21313),
            .lcout(\POWERLED.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__21447),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(\POWERLED.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__19339),
            .in2(N__19548),
            .in3(N__19333),
            .lcout(\POWERLED.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__19544),
            .in2(N__21208),
            .in3(N__19321),
            .lcout(\POWERLED.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__21400),
            .in2(N__21325),
            .in3(N__19564),
            .lcout(\POWERLED.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(N__21324),
            .in2(N__21388),
            .in3(N__19552),
            .lcout(\POWERLED.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_6_5  (
            .in0(N__19421),
            .in1(N__21373),
            .in2(N__19549),
            .in3(N__19522),
            .lcout(\POWERLED.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_6_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(N__21340),
            .in2(_gnd_net_),
            .in3(N__19519),
            .lcout(\POWERLED.mult1_un117_sum_s_8 ),
            .ltout(\POWERLED.mult1_un117_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_6_6_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_6_6_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_6_6_7  (
            .in0(N__19516),
            .in1(_gnd_net_),
            .in2(N__19504),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un124_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_6_7_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_6_7_0 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_LC_6_7_0  (
            .in0(N__19492),
            .in1(N__19480),
            .in2(N__32323),
            .in3(N__19437),
            .lcout(\PCH_PWRGD.delayed_vccin_ok_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32508),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_7_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19415),
            .lcout(\POWERLED.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_1_LC_6_7_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_1_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_1_LC_6_7_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.func_state_RNI_0_1_LC_6_7_6  (
            .in0(_gnd_net_),
            .in1(N__31879),
            .in2(_gnd_net_),
            .in3(N__28815),
            .lcout(\POWERLED.N_341 ),
            .ltout(\POWERLED.N_341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_3_1_LC_6_7_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_3_1_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_3_1_LC_6_7_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.func_state_RNI_3_1_LC_6_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19687),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_341_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_1_LC_6_8_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_5_1_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_1_LC_6_8_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \POWERLED.dutycycle_RNI_5_1_LC_6_8_0  (
            .in0(_gnd_net_),
            .in1(N__31470),
            .in2(_gnd_net_),
            .in3(N__31548),
            .lcout(\POWERLED.dutycycle_RNI_5Z0Z_1 ),
            .ltout(),
            .carryin(bfn_6_8_0_),
            .carryout(\POWERLED.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_6_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_6_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_6_8_1  (
            .in0(_gnd_net_),
            .in1(N__21523),
            .in2(N__19656),
            .in3(N__19606),
            .lcout(G_2129),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_0 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_6_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_6_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_6_8_2  (
            .in0(_gnd_net_),
            .in1(N__19652),
            .in2(N__19684),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_6_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_6_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_6_8_3  (
            .in0(_gnd_net_),
            .in1(N__19675),
            .in2(N__19615),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_6_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_6_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_6_8_4  (
            .in0(_gnd_net_),
            .in1(N__19669),
            .in2(N__19614),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_6_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_6_8_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_6_8_5  (
            .in0(_gnd_net_),
            .in1(N__19663),
            .in2(N__19657),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_6_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_6_8_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_6_8_6  (
            .in0(N__19636),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19630),
            .lcout(\POWERLED.un85_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_6_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_6_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_6_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19605),
            .lcout(\POWERLED.un85_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_LC_6_9_0 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_LC_6_9_0 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_LC_6_9_0  (
            .in0(N__19719),
            .in1(N__19726),
            .in2(N__19904),
            .in3(N__30748),
            .lcout(\POWERLED.un1_func_state25_6_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_1_1_LC_6_9_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_1_1_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_1_1_LC_6_9_1 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \POWERLED.func_state_RNI5DLR_1_1_LC_6_9_1  (
            .in0(N__28760),
            .in1(N__30381),
            .in2(_gnd_net_),
            .in3(N__30522),
            .lcout(\POWERLED.func_state_RNI5DLR_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_0_LC_6_9_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_0_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_0_LC_6_9_2 .LUT_INIT=16'b0000101011101110;
    LogicCell40 \POWERLED.func_state_RNI_1_0_LC_6_9_2  (
            .in0(N__19891),
            .in1(N__31851),
            .in2(N__22874),
            .in3(N__28759),
            .lcout(),
            .ltout(\POWERLED.N_394_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI25Q51_0_LC_6_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI25Q51_0_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI25Q51_0_LC_6_9_3 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \POWERLED.func_state_RNI25Q51_0_LC_6_9_3  (
            .in0(N__31787),
            .in1(_gnd_net_),
            .in2(N__19762),
            .in3(N__25000),
            .lcout(\POWERLED.N_453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI0N7A2_1_LC_6_9_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI0N7A2_1_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI0N7A2_1_LC_6_9_4 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \POWERLED.func_state_RNI0N7A2_1_LC_6_9_4  (
            .in0(N__19740),
            .in1(N__33924),
            .in2(N__28830),
            .in3(N__21508),
            .lcout(\POWERLED.func_state_1_m0_i_o2_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_0_0_LC_6_9_5 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_0_0_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_0_0_LC_6_9_5 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_0_0_LC_6_9_5  (
            .in0(N__31789),
            .in1(N__30383),
            .in2(_gnd_net_),
            .in3(N__23369),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_0_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_LC_6_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_LC_6_9_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_LC_6_9_6  (
            .in0(N__22857),
            .in1(N__19896),
            .in2(N__19729),
            .in3(N__28761),
            .lcout(\POWERLED.un1_func_state25_6_0_o_N_422_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_count_off_0_sqmuxa_4_i_0_a2_LC_6_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_count_off_0_sqmuxa_4_i_0_a2_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_count_off_0_sqmuxa_4_i_0_a2_LC_6_9_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_count_off_0_sqmuxa_4_i_0_a2_LC_6_9_7  (
            .in0(N__31788),
            .in1(N__30382),
            .in2(_gnd_net_),
            .in3(N__23368),
            .lcout(\POWERLED.un1_func_state25_6_0_o_N_516_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_en_LC_6_10_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_en_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_en_LC_6_10_0 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \POWERLED.count_off_en_LC_6_10_0  (
            .in0(N__19708),
            .in1(N__19702),
            .in2(N__19696),
            .in3(N__28026),
            .lcout(\POWERLED.count_off_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_EN_i_0_o3_LC_6_10_1 .C_ON=1'b0;
    defparam \POWERLED.VCCST_EN_i_0_o3_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_EN_i_0_o3_LC_6_10_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \POWERLED.VCCST_EN_i_0_o3_LC_6_10_1  (
            .in0(N__30534),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31180),
            .lcout(VCCST_EN_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_LC_6_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_0_LC_6_10_2 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \POWERLED.func_state_0_LC_6_10_2  (
            .in0(N__19789),
            .in1(N__19780),
            .in2(N__22988),
            .in3(N__28027),
            .lcout(\POWERLED.func_stateZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32630),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIOGRS_0_LC_6_10_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIOGRS_0_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIOGRS_0_LC_6_10_3 .LUT_INIT=16'b1000010101010101;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_fast_RNIOGRS_0_LC_6_10_3  (
            .in0(N__21502),
            .in1(N__26421),
            .in2(N__19915),
            .in3(N__31181),
            .lcout(\RSMRST_PWRGD.N_8_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI0N7A2_0_1_LC_6_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI0N7A2_0_1_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI0N7A2_0_1_LC_6_10_4 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \POWERLED.func_state_RNI0N7A2_0_1_LC_6_10_4  (
            .in0(N__19895),
            .in1(N__19827),
            .in2(_gnd_net_),
            .in3(N__19816),
            .lcout(),
            .ltout(\POWERLED.N_143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNICK8N9_1_LC_6_10_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNICK8N9_1_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNICK8N9_1_LC_6_10_5 .LUT_INIT=16'b0000000010001101;
    LogicCell40 \POWERLED.func_state_RNICK8N9_1_LC_6_10_5  (
            .in0(N__21774),
            .in1(N__19810),
            .in2(N__19792),
            .in3(N__23339),
            .lcout(\POWERLED.func_state_RNICK8N9Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIE4QDD_0_LC_6_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIE4QDD_0_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIE4QDD_0_LC_6_10_6 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \POWERLED.func_state_RNIE4QDD_0_LC_6_10_6  (
            .in0(N__19788),
            .in1(N__28025),
            .in2(N__22987),
            .in3(N__19779),
            .lcout(\POWERLED.func_stateZ0Z_0 ),
            .ltout(\POWERLED.func_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_2_0_LC_6_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_2_0_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_2_0_LC_6_10_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.func_state_RNI_2_0_LC_6_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19771),
            .in3(_gnd_net_),
            .lcout(func_state_RNI_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI2S6S9_10_LC_6_11_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI2S6S9_10_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI2S6S9_10_LC_6_11_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \POWERLED.count_off_RNI2S6S9_10_LC_6_11_0  (
            .in0(N__19768),
            .in1(_gnd_net_),
            .in2(N__20086),
            .in3(N__20590),
            .lcout(\POWERLED.count_offZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_10_LC_6_11_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_10_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_10_LC_6_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_10_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20082),
            .lcout(\POWERLED.count_off_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32650),
            .ce(N__20621),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIB3KQ9_11_LC_6_11_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIB3KQ9_11_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIB3KQ9_11_LC_6_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_off_RNIB3KQ9_11_LC_6_11_2  (
            .in0(N__20050),
            .in1(N__20035),
            .in2(_gnd_net_),
            .in3(N__20591),
            .lcout(\POWERLED.count_offZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_11_LC_6_11_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_11_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_11_LC_6_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_11_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20049),
            .lcout(\POWERLED.count_off_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32650),
            .ce(N__20621),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIBSPT9_2_LC_6_11_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIBSPT9_2_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIBSPT9_2_LC_6_11_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIBSPT9_2_LC_6_11_4  (
            .in0(N__20029),
            .in1(N__19953),
            .in2(_gnd_net_),
            .in3(N__20589),
            .lcout(\POWERLED.count_offZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_2_LC_6_11_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_2_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_2_LC_6_11_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_2_LC_6_11_5  (
            .in0(N__19954),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32650),
            .ce(N__20621),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNID6LQ9_12_LC_6_11_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNID6LQ9_12_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNID6LQ9_12_LC_6_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_off_RNID6LQ9_12_LC_6_11_6  (
            .in0(N__20446),
            .in1(N__20023),
            .in2(_gnd_net_),
            .in3(N__20592),
            .lcout(\POWERLED.count_offZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_12_LC_6_11_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_12_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_12_LC_6_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_12_LC_6_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20445),
            .lcout(\POWERLED.count_off_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32650),
            .ce(N__20621),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_6_12_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_6_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_LC_6_12_0  (
            .in0(_gnd_net_),
            .in1(N__20011),
            .in2(N__19989),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_12_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI2QT43_LC_6_12_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI2QT43_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI2QT43_LC_6_12_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_RNI2QT43_LC_6_12_1  (
            .in0(N__20365),
            .in1(N__19965),
            .in2(_gnd_net_),
            .in3(N__19945),
            .lcout(\POWERLED.count_off_1_2 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_1 ),
            .carryout(\POWERLED.un3_count_off_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_6_12_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_6_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(N__19938),
            .in2(_gnd_net_),
            .in3(N__19918),
            .lcout(\POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_2 ),
            .carryout(\POWERLED.un3_count_off_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_6_12_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_6_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_6_12_3  (
            .in0(_gnd_net_),
            .in1(N__20218),
            .in2(_gnd_net_),
            .in3(N__20182),
            .lcout(\POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_3 ),
            .carryout(\POWERLED.un3_count_off_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI50153_LC_6_12_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI50153_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI50153_LC_6_12_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_4_c_RNI50153_LC_6_12_4  (
            .in0(N__20368),
            .in1(N__20178),
            .in2(_gnd_net_),
            .in3(N__20149),
            .lcout(\POWERLED.count_off_1_5 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_4 ),
            .carryout(\POWERLED.un3_count_off_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI62253_LC_6_12_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI62253_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI62253_LC_6_12_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_5_c_RNI62253_LC_6_12_5  (
            .in0(N__20366),
            .in1(N__20142),
            .in2(_gnd_net_),
            .in3(N__20113),
            .lcout(\POWERLED.count_off_1_6 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_5 ),
            .carryout(\POWERLED.un3_count_off_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNI74353_LC_6_12_6 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNI74353_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNI74353_LC_6_12_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_6_c_RNI74353_LC_6_12_6  (
            .in0(N__20369),
            .in1(N__20232),
            .in2(_gnd_net_),
            .in3(N__20110),
            .lcout(\POWERLED.count_off_1_7 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_6 ),
            .carryout(\POWERLED.un3_count_off_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNI86453_LC_6_12_7 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNI86453_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNI86453_LC_6_12_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_7_c_RNI86453_LC_6_12_7  (
            .in0(N__20367),
            .in1(N__20676),
            .in2(_gnd_net_),
            .in3(N__20107),
            .lcout(\POWERLED.count_off_1_8 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_7 ),
            .carryout(\POWERLED.un3_count_off_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNI98553_LC_6_13_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNI98553_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNI98553_LC_6_13_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_8_c_RNI98553_LC_6_13_0  (
            .in0(N__20382),
            .in1(N__20277),
            .in2(_gnd_net_),
            .in3(N__20104),
            .lcout(\POWERLED.count_off_1_9 ),
            .ltout(),
            .carryin(bfn_6_13_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIAA653_LC_6_13_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIAA653_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIAA653_LC_6_13_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_9_c_RNIAA653_LC_6_13_1  (
            .in0(N__20371),
            .in1(N__20101),
            .in2(_gnd_net_),
            .in3(N__20071),
            .lcout(\POWERLED.count_off_1_10 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_9 ),
            .carryout(\POWERLED.un3_count_off_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIIGJ33_LC_6_13_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIIGJ33_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIIGJ33_LC_6_13_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_10_c_RNIIGJ33_LC_6_13_2  (
            .in0(N__20381),
            .in1(N__20068),
            .in2(_gnd_net_),
            .in3(N__20038),
            .lcout(\POWERLED.count_off_1_11 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_10 ),
            .carryout(\POWERLED.un3_count_off_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIJIK33_LC_6_13_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIJIK33_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIJIK33_LC_6_13_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_11_c_RNIJIK33_LC_6_13_3  (
            .in0(N__20370),
            .in1(N__20461),
            .in2(_gnd_net_),
            .in3(N__20434),
            .lcout(\POWERLED.count_off_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_11 ),
            .carryout(\POWERLED.un3_count_off_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNIKKL33_LC_6_13_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNIKKL33_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNIKKL33_LC_6_13_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_12_c_RNIKKL33_LC_6_13_4  (
            .in0(N__20383),
            .in1(N__20431),
            .in2(_gnd_net_),
            .in3(N__20410),
            .lcout(\POWERLED.count_off_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_12 ),
            .carryout(\POWERLED.un3_count_off_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNILMM33_LC_6_13_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNILMM33_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNILMM33_LC_6_13_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_13_c_RNILMM33_LC_6_13_5  (
            .in0(N__20372),
            .in1(N__20407),
            .in2(_gnd_net_),
            .in3(N__20386),
            .lcout(\POWERLED.count_off_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_13 ),
            .carryout(\POWERLED.un3_count_off_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIMON33_LC_6_13_6 .C_ON=1'b0;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIMON33_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIMON33_LC_6_13_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_14_c_RNIMON33_LC_6_13_6  (
            .in0(N__20266),
            .in1(N__20373),
            .in2(_gnd_net_),
            .in3(N__20284),
            .lcout(\POWERLED.un3_count_off_1_cry_14_c_RNIMONZ0Z33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIPH1U9_9_LC_6_13_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIPH1U9_9_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIPH1U9_9_LC_6_13_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_off_RNIPH1U9_9_LC_6_13_7  (
            .in0(N__20644),
            .in1(N__20632),
            .in2(_gnd_net_),
            .in3(N__20605),
            .lcout(\POWERLED.count_offZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIJFOQ9_15_LC_6_14_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIJFOQ9_15_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIJFOQ9_15_LC_6_14_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIJFOQ9_15_LC_6_14_0  (
            .in0(N__20242),
            .in1(N__20250),
            .in2(_gnd_net_),
            .in3(N__20540),
            .lcout(\POWERLED.count_offZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_15_LC_6_14_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_15_LC_6_14_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_15_LC_6_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_15_LC_6_14_1  (
            .in0(N__20251),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33041),
            .ce(N__20617),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNILBVT9_7_LC_6_14_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNILBVT9_7_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNILBVT9_7_LC_6_14_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_off_RNILBVT9_7_LC_6_14_2  (
            .in0(N__20694),
            .in1(N__20683),
            .in2(_gnd_net_),
            .in3(N__20541),
            .lcout(\POWERLED.count_offZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_7_LC_6_14_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_7_LC_6_14_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_7_LC_6_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_7_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20695),
            .lcout(\POWERLED.count_off_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33041),
            .ce(N__20617),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNINE0U9_8_LC_6_14_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNINE0U9_8_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNINE0U9_8_LC_6_14_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_off_RNINE0U9_8_LC_6_14_4  (
            .in0(N__20662),
            .in1(N__20650),
            .in2(_gnd_net_),
            .in3(N__20539),
            .lcout(\POWERLED.count_offZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_8_LC_6_14_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_8_LC_6_14_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_8_LC_6_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_8_LC_6_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20661),
            .lcout(\POWERLED.count_off_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33041),
            .ce(N__20617),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_9_LC_6_14_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_9_LC_6_14_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_9_LC_6_14_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \POWERLED.count_off_9_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(N__20643),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33041),
            .ce(N__20617),
            .sr(_gnd_net_));
    defparam \POWERLED.G_10_LC_6_15_7 .C_ON=1'b0;
    defparam \POWERLED.G_10_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_10_LC_6_15_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.G_10_LC_6_15_7  (
            .in0(_gnd_net_),
            .in1(N__33930),
            .in2(_gnd_net_),
            .in3(N__21753),
            .lcout(G_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_1_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_1_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21964),
            .lcout(\POWERLED.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_7_1_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_7_1_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_7_1_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_7_1_2  (
            .in0(N__22053),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_1_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_1_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_1_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_1_3  (
            .in0(N__22102),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_7_1_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_7_1_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_7_1_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_7_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22470),
            .lcout(\POWERLED.un85_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_6_LC_7_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_6_LC_7_1_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_6_LC_7_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_6_LC_7_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21193),
            .lcout(\PCH_PWRGD.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32367),
            .ce(N__21157),
            .sr(N__20996));
    defparam CONSTANT_ONE_LUT4_LC_7_1_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_1_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_1_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_0_LC_7_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_0_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_0_LC_7_2_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_0_LC_7_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20788),
            .lcout(pch_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_7_2_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_7_2_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_7_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23904),
            .lcout(\POWERLED.mult1_un54_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_7_2_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_7_2_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_7_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26007),
            .lcout(\POWERLED.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_7_2_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_7_2_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_7_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25725),
            .lcout(\POWERLED.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_7_2_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_7_2_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_7_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25623),
            .lcout(\POWERLED.mult1_un68_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_7_2_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_7_2_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_7_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23809),
            .lcout(\POWERLED.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_7_2_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_7_2_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_7_2_6  (
            .in0(N__23704),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un75_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_2_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_2_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_2_7  (
            .in0(N__23601),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_6_LC_7_3_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_6_LC_7_3_0 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_6_LC_7_3_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \POWERLED.dutycycle_6_LC_7_3_0  (
            .in0(N__22746),
            .in1(N__24343),
            .in2(N__28147),
            .in3(N__22762),
            .lcout(\POWERLED.dutycycle_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32418),
            .ce(),
            .sr(N__26632));
    defparam \POWERLED.dutycycle_7_LC_7_3_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_7_LC_7_3_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_7_LC_7_3_1 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \POWERLED.dutycycle_7_LC_7_3_1  (
            .in0(N__24268),
            .in1(N__21544),
            .in2(N__21667),
            .in3(N__31081),
            .lcout(\POWERLED.dutycycleZ1Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32418),
            .ce(),
            .sr(N__26632));
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_3_2 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_3_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24084),
            .lcout(\POWERLED.un1_dutycycle_53_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_3_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_3_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_3_3  (
            .in0(N__22201),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_7_3_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_7_3_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_7_3_4  (
            .in0(N__22492),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_7_3_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_7_3_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_7_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22491),
            .lcout(\POWERLED.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_7_3_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_7_3_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_7_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21320),
            .lcout(\POWERLED.un85_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_4_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_4_0  (
            .in0(_gnd_net_),
            .in1(N__21433),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_4_0_),
            .carryout(\POWERLED.mult1_un110_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_4_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_4_1  (
            .in0(_gnd_net_),
            .in1(N__21217),
            .in2(N__21357),
            .in3(N__21196),
            .lcout(\POWERLED.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_4_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_4_2  (
            .in0(_gnd_net_),
            .in1(N__21353),
            .in2(N__22177),
            .in3(N__21391),
            .lcout(\POWERLED.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_4_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_4_3  (
            .in0(_gnd_net_),
            .in1(N__22156),
            .in2(N__22498),
            .in3(N__21376),
            .lcout(\POWERLED.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_4_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_4_4  (
            .in0(_gnd_net_),
            .in1(N__22497),
            .in2(N__22138),
            .in3(N__21361),
            .lcout(\POWERLED.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_4_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_4_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_4_5  (
            .in0(N__21314),
            .in1(N__22120),
            .in2(N__21358),
            .in3(N__21331),
            .lcout(\POWERLED.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_4_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_4_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22522),
            .in3(N__21328),
            .lcout(\POWERLED.mult1_un110_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_7_4_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_7_4_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_7_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23845),
            .lcout(\POWERLED.un85_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_LC_7_5_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_0_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_LC_7_5_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_LC_7_5_0  (
            .in0(_gnd_net_),
            .in1(N__28966),
            .in2(N__31480),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un145_sum ),
            .ltout(),
            .carryin(bfn_7_5_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_0_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_5_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_5_1  (
            .in0(_gnd_net_),
            .in1(N__31478),
            .in2(N__21535),
            .in3(N__21253),
            .lcout(\POWERLED.mult1_un138_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_0_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_5_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_5_2  (
            .in0(_gnd_net_),
            .in1(N__22594),
            .in2(N__26428),
            .in3(N__21232),
            .lcout(\POWERLED.mult1_un131_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_1_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_5_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_5_3  (
            .in0(_gnd_net_),
            .in1(N__26425),
            .in2(N__21595),
            .in3(N__21451),
            .lcout(\POWERLED.mult1_un124_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_2_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_3_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_5_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_5_4  (
            .in0(_gnd_net_),
            .in1(N__21562),
            .in2(N__21616),
            .in3(N__21436),
            .lcout(\POWERLED.mult1_un117_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_3_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_4_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_5_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_5_5  (
            .in0(_gnd_net_),
            .in1(N__30871),
            .in2(N__22582),
            .in3(N__21418),
            .lcout(\POWERLED.mult1_un110_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_4_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_5_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_5_6  (
            .in0(_gnd_net_),
            .in1(N__27733),
            .in2(N__30879),
            .in3(N__21415),
            .lcout(\POWERLED.mult1_un103_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_5_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_6_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_5_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_5_7  (
            .in0(_gnd_net_),
            .in1(N__26026),
            .in2(N__30019),
            .in3(N__21412),
            .lcout(\POWERLED.mult1_un96_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_6_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__30159),
            .in2(N__22552),
            .in3(N__21409),
            .lcout(\POWERLED.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_7_6_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__29483),
            .in2(N__22537),
            .in3(N__21406),
            .lcout(\POWERLED.mult1_un82_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_8 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__22543),
            .in2(N__26116),
            .in3(N__21403),
            .lcout(\POWERLED.mult1_un75_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__28351),
            .in2(N__28288),
            .in3(N__21496),
            .lcout(\POWERLED.mult1_un68_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(N__28640),
            .in2(N__22603),
            .in3(N__21493),
            .lcout(\POWERLED.mult1_un61_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_6_5  (
            .in0(_gnd_net_),
            .in1(N__26114),
            .in2(N__26056),
            .in3(N__21490),
            .lcout(\POWERLED.mult1_un54_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_6_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(N__24157),
            .in2(N__28357),
            .in3(N__21487),
            .lcout(\POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_6_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_6_7  (
            .in0(_gnd_net_),
            .in1(N__28641),
            .in2(N__24181),
            .in3(N__21484),
            .lcout(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_14 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__28642),
            .in2(N__24208),
            .in3(N__21481),
            .lcout(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\POWERLED.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_7_1 .C_ON=1'b0;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.CO2_THRU_LUT4_0_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21478),
            .lcout(\POWERLED.CO2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_7_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_7_2 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__22276),
            .in2(N__22320),
            .in3(N__22298),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOGRS_4_LC_7_7_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOGRS_4_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOGRS_4_LC_7_7_4 .LUT_INIT=16'b1111111100001100;
    LogicCell40 \POWERLED.dutycycle_RNIOGRS_4_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__31017),
            .in2(N__29261),
            .in3(N__28468),
            .lcout(\POWERLED.N_76_f0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIFOI43_4_LC_7_7_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIFOI43_4_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIFOI43_4_LC_7_7_6 .LUT_INIT=16'b1000000010101010;
    LogicCell40 \POWERLED.dutycycle_RNIFOI43_4_LC_7_7_6  (
            .in0(N__28091),
            .in1(N__28215),
            .in2(N__31775),
            .in3(N__21475),
            .lcout(\POWERLED.dutycycle_en_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_1_LC_7_7_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_1_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_1_LC_7_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_4_1_LC_7_7_7  (
            .in0(N__31460),
            .in1(N__29224),
            .in2(_gnd_net_),
            .in3(N__31524),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_7_8_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_7_8_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_7_8_0  (
            .in0(N__31523),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_8_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26396),
            .lcout(\POWERLED.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_eena_5_0_s_tz_iso_LC_7_8_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_eena_5_0_s_tz_iso_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_eena_5_0_s_tz_iso_LC_7_8_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.dutycycle_eena_5_0_s_tz_iso_LC_7_8_3  (
            .in0(N__23370),
            .in1(N__30374),
            .in2(N__33999),
            .in3(N__31753),
            .lcout(\POWERLED.dutycycle_eena_5_0_s_tz_isoZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_1_LC_7_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_1_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_1_LC_7_8_5 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_1_LC_7_8_5  (
            .in0(_gnd_net_),
            .in1(N__31522),
            .in2(N__29304),
            .in3(N__30852),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNID4591_1_LC_7_8_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNID4591_1_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNID4591_1_LC_7_8_6 .LUT_INIT=16'b0010000011111111;
    LogicCell40 \POWERLED.func_state_RNID4591_1_LC_7_8_6  (
            .in0(N__30375),
            .in1(N__31764),
            .in2(N__26754),
            .in3(N__21808),
            .lcout(\POWERLED.func_state_1_m0_i_o2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_13_LC_7_8_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_13_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_13_LC_7_8_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.dutycycle_RNI_2_13_LC_7_8_7  (
            .in0(N__26110),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_2187_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_LC_7_9_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_LC_7_9_0 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \POWERLED.dutycycle_RNI_9_LC_7_9_0  (
            .in0(N__31287),
            .in1(N__26953),
            .in2(N__29887),
            .in3(N__22693),
            .lcout(N_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNITGMHB_1_LC_7_9_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNITGMHB_1_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNITGMHB_1_LC_7_9_2 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \POWERLED.func_state_RNITGMHB_1_LC_7_9_2  (
            .in0(N__22983),
            .in1(N__28028),
            .in2(N__21574),
            .in3(N__21582),
            .lcout(func_state_RNITGMHB_0_1),
            .ltout(func_state_RNITGMHB_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOGRS_1_LC_7_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOGRS_1_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOGRS_1_LC_7_9_3 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \POWERLED.func_state_RNIOGRS_1_LC_7_9_3  (
            .in0(N__30244),
            .in1(N__30523),
            .in2(N__21619),
            .in3(N__31183),
            .lcout(func_state_RNIOGRS_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_LC_7_9_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_LC_7_9_4 .LUT_INIT=16'b1110100011101000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_LC_7_9_4  (
            .in0(N__21604),
            .in1(N__28923),
            .in2(N__31345),
            .in3(N__21561),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_LC_7_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_LC_7_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_2_LC_7_9_5  (
            .in0(N__26415),
            .in1(N__21603),
            .in2(N__28944),
            .in3(N__31283),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_LC_7_9_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_1_LC_7_9_6 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \POWERLED.func_state_1_LC_7_9_6  (
            .in0(N__21573),
            .in1(N__28029),
            .in2(N__22990),
            .in3(N__21583),
            .lcout(\POWERLED.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32507),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_3_LC_7_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_7_9_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNI_4_3_LC_7_9_7  (
            .in0(N__28922),
            .in1(_gnd_net_),
            .in2(N__29305),
            .in3(N__29027),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_rep1_LC_7_10_0 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_rep1_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_rep1_LC_7_10_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \COUNTER.tmp_0_rep1_LC_7_10_0  (
            .in0(N__23019),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21751),
            .lcout(SUSWARN_N_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32629),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_156_LC_7_10_1 .C_ON=1'b0;
    defparam \POWERLED.G_156_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_156_LC_7_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.G_156_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__23017),
            .in2(_gnd_net_),
            .in3(N__21749),
            .lcout(G_156),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_7_LC_7_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_7_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_7_LC_7_10_2 .LUT_INIT=16'b1011101110111010;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_7_LC_7_10_2  (
            .in0(N__28435),
            .in1(N__29031),
            .in2(N__24807),
            .in3(N__28780),
            .lcout(),
            .ltout(\POWERLED.N_80_f0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI375F3_7_LC_7_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI375F3_7_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI375F3_7_LC_7_10_3 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI375F3_7_LC_7_10_3  (
            .in0(N__28553),
            .in1(N__23018),
            .in2(N__21547),
            .in3(N__21750),
            .lcout(\POWERLED.dutycycle_RNI375F3Z0Z_7 ),
            .ltout(\POWERLED.dutycycle_RNI375F3Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIPENJ4_7_LC_7_10_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIPENJ4_7_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIPENJ4_7_LC_7_10_4 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \POWERLED.dutycycle_RNIPENJ4_7_LC_7_10_4  (
            .in0(N__21666),
            .in1(N__24264),
            .in2(N__21649),
            .in3(N__30983),
            .lcout(\POWERLED.dutycycleZ0Z_4 ),
            .ltout(\POWERLED.dutycycleZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_4_LC_7_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_4_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_4_LC_7_10_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \POWERLED.dutycycle_RNI_2_4_LC_7_10_5  (
            .in0(N__29306),
            .in1(_gnd_net_),
            .in2(N__21646),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(m57_i_o2_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIQ8072_LC_7_10_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIQ8072_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIQ8072_LC_7_10_6 .LUT_INIT=16'b0011001100110101;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_fast_RNIQ8072_LC_7_10_6  (
            .in0(N__21643),
            .in1(N__26899),
            .in2(N__21637),
            .in3(N__24367),
            .lcout(),
            .ltout(\RSMRST_PWRGD.N_4713_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIO5AE5_LC_7_10_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIO5AE5_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIO5AE5_LC_7_10_7 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_fast_RNIO5AE5_LC_7_10_7  (
            .in0(N__24953),
            .in1(N__26665),
            .in2(N__21634),
            .in3(N__28555),
            .lcout(\RSMRST_PWRGD.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_6_0_LC_7_11_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_6_0_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_6_0_LC_7_11_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \POWERLED.func_state_RNI_6_0_LC_7_11_0  (
            .in0(N__30699),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23031),
            .lcout(),
            .ltout(\POWERLED.N_569_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_2_1_LC_7_11_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_2_1_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_2_1_LC_7_11_1 .LUT_INIT=16'b0011001101000000;
    LogicCell40 \POWERLED.func_state_RNI5DLR_2_1_LC_7_11_1  (
            .in0(N__28858),
            .in1(N__30528),
            .in2(N__21631),
            .in3(N__30371),
            .lcout(),
            .ltout(\POWERLED.N_220_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI1PE62_1_LC_7_11_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI1PE62_1_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI1PE62_1_LC_7_11_2 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \POWERLED.func_state_RNI1PE62_1_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__26926),
            .in2(N__21628),
            .in3(N__24684),
            .lcout(\POWERLED.N_282_N ),
            .ltout(\POWERLED.N_282_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIB0O42_3_LC_7_11_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIB0O42_3_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIB0O42_3_LC_7_11_3 .LUT_INIT=16'b1111111100001011;
    LogicCell40 \POWERLED.dutycycle_RNIB0O42_3_LC_7_11_3  (
            .in0(N__28909),
            .in1(N__31052),
            .in2(N__21625),
            .in3(N__28198),
            .lcout(),
            .ltout(\POWERLED.dutycycle_eena_8_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI79E14_3_LC_7_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI79E14_3_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI79E14_3_LC_7_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI79E14_3_LC_7_11_4  (
            .in0(N__21859),
            .in1(N__23020),
            .in2(N__21622),
            .in3(N__21752),
            .lcout(\POWERLED.dutycycle_RNI79E14Z0Z_3 ),
            .ltout(\POWERLED.dutycycle_RNI79E14Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIL4S55_3_LC_7_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIL4S55_3_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIL4S55_3_LC_7_11_5 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \POWERLED.dutycycle_RNIL4S55_3_LC_7_11_5  (
            .in0(N__24306),
            .in1(N__21843),
            .in2(N__21865),
            .in3(N__31049),
            .lcout(\POWERLED.dutycycleZ0Z_6 ),
            .ltout(\POWERLED.dutycycleZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIRKB61_3_LC_7_11_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIRKB61_3_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIRKB61_3_LC_7_11_6 .LUT_INIT=16'b1100110011111101;
    LogicCell40 \POWERLED.dutycycle_RNIRKB61_3_LC_7_11_6  (
            .in0(N__31050),
            .in1(N__31776),
            .in2(N__21862),
            .in3(N__28436),
            .lcout(\POWERLED.dutycycle_eena_8_c ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_3_LC_7_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_3_LC_7_11_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_3_LC_7_11_7 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \POWERLED.dutycycle_3_LC_7_11_7  (
            .in0(N__24307),
            .in1(N__21853),
            .in2(N__21847),
            .in3(N__31051),
            .lcout(\POWERLED.dutycycleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32637),
            .ce(),
            .sr(N__26653));
    defparam \POWERLED.func_state_RNI_1_1_LC_7_12_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_1_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_1_LC_7_12_0 .LUT_INIT=16'b0101110101010101;
    LogicCell40 \POWERLED.func_state_RNI_1_1_LC_7_12_0  (
            .in0(N__30764),
            .in1(N__24757),
            .in2(N__28859),
            .in3(N__24742),
            .lcout(\POWERLED.N_52_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.N_52_i_i_x2_LC_7_12_1 .C_ON=1'b0;
    defparam \POWERLED.N_52_i_i_x2_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.N_52_i_i_x2_LC_7_12_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \POWERLED.N_52_i_i_x2_LC_7_12_1  (
            .in0(N__30547),
            .in1(_gnd_net_),
            .in2(N__30386),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.N_231_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBVNS_1_LC_7_12_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_1_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_1_LC_7_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.func_state_RNIBVNS_1_LC_7_12_2  (
            .in0(N__21832),
            .in1(N__28834),
            .in2(N__21811),
            .in3(N__25124),
            .lcout(),
            .ltout(\POWERLED.N_410_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI1J4E2_1_LC_7_12_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI1J4E2_1_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI1J4E2_1_LC_7_12_3 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \POWERLED.func_state_RNI1J4E2_1_LC_7_12_3  (
            .in0(N__21807),
            .in1(N__21787),
            .in2(N__21781),
            .in3(N__28205),
            .lcout(\POWERLED.func_state_RNI1J4E2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_fast_LC_7_12_4 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_fast_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_fast_LC_7_12_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \COUNTER.tmp_0_fast_LC_7_12_4  (
            .in0(N__24627),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21757),
            .lcout(SUSWARN_N_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32754),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.N_52_i_i_a2_LC_7_12_7 .C_ON=1'b0;
    defparam \POWERLED.N_52_i_i_a2_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.N_52_i_i_a2_LC_7_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.N_52_i_i_a2_LC_7_12_7  (
            .in0(N__30546),
            .in1(N__24626),
            .in2(N__30385),
            .in3(N__31179),
            .lcout(\POWERLED.N_507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_44_LC_7_13_0 .C_ON=1'b0;
    defparam \POWERLED.G_44_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_44_LC_7_13_0 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \POWERLED.G_44_LC_7_13_0  (
            .in0(N__23419),
            .in1(N__23437),
            .in2(N__21898),
            .in3(N__27523),
            .lcout(G_44),
            .ltout(G_44_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_7_13_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_7_13_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \VPP_VDDQ.count_esr_RNO_0_15_LC_7_13_1  (
            .in0(N__27524),
            .in1(_gnd_net_),
            .in2(N__21901),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.N_42_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNI8I855_0_LC_7_13_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNI8I855_0_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNI8I855_0_LC_7_13_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.curr_state_RNI8I855_0_LC_7_13_2  (
            .in0(N__23417),
            .in1(N__23458),
            .in2(_gnd_net_),
            .in3(N__23217),
            .lcout(N_365),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_1_LC_7_13_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_1_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_1_LC_7_13_3 .LUT_INIT=16'b0001101100001010;
    LogicCell40 \VPP_VDDQ.curr_state_1_LC_7_13_3  (
            .in0(N__23461),
            .in1(N__23308),
            .in2(N__23221),
            .in3(N__23420),
            .lcout(\VPP_VDDQ.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32752),
            .ce(N__27386),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_0_LC_7_13_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_0_LC_7_13_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_0_LC_7_13_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \VPP_VDDQ.curr_state_0_LC_7_13_4  (
            .in0(N__23307),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23460),
            .lcout(VPP_VDDQ_curr_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32752),
            .ce(N__27386),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_7_13_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_7_13_5 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_7_13_5  (
            .in0(N__23459),
            .in1(N__23306),
            .in2(_gnd_net_),
            .in3(N__23418),
            .lcout(\VPP_VDDQ.N_464_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_0_LC_7_14_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_0_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_0_LC_7_14_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_0_LC_7_14_0  (
            .in0(N__27541),
            .in1(N__23194),
            .in2(N__21889),
            .in3(N__21888),
            .lcout(\VPP_VDDQ.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_0 ),
            .clk(N__32755),
            .ce(),
            .sr(N__21997));
    defparam \VPP_VDDQ.count_1_LC_7_14_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_1_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_1_LC_7_14_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_1_LC_7_14_1  (
            .in0(N__27533),
            .in1(N__23638),
            .in2(_gnd_net_),
            .in3(N__21874),
            .lcout(\VPP_VDDQ.countZ0Z_1 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_0 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_1 ),
            .clk(N__32755),
            .ce(),
            .sr(N__21997));
    defparam \VPP_VDDQ.count_2_LC_7_14_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_2_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_LC_7_14_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_2_LC_7_14_2  (
            .in0(N__27542),
            .in1(N__23665),
            .in2(_gnd_net_),
            .in3(N__21871),
            .lcout(\VPP_VDDQ.countZ0Z_2 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_2 ),
            .clk(N__32755),
            .ce(),
            .sr(N__21997));
    defparam \VPP_VDDQ.count_3_LC_7_14_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_3_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_3_LC_7_14_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_3_LC_7_14_3  (
            .in0(N__27534),
            .in1(N__23487),
            .in2(_gnd_net_),
            .in3(N__21868),
            .lcout(\VPP_VDDQ.countZ0Z_3 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_3 ),
            .clk(N__32755),
            .ce(),
            .sr(N__21997));
    defparam \VPP_VDDQ.count_4_LC_7_14_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_4_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_4_LC_7_14_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_4_LC_7_14_4  (
            .in0(N__27543),
            .in1(N__23500),
            .in2(_gnd_net_),
            .in3(N__21928),
            .lcout(\VPP_VDDQ.countZ0Z_4 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_4 ),
            .clk(N__32755),
            .ce(),
            .sr(N__21997));
    defparam \VPP_VDDQ.count_5_LC_7_14_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_5_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_5_LC_7_14_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_5_LC_7_14_5  (
            .in0(N__27535),
            .in1(N__23512),
            .in2(_gnd_net_),
            .in3(N__21925),
            .lcout(\VPP_VDDQ.countZ0Z_5 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_5 ),
            .clk(N__32755),
            .ce(),
            .sr(N__21997));
    defparam \VPP_VDDQ.count_6_LC_7_14_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_6_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_6_LC_7_14_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_6_LC_7_14_6  (
            .in0(N__27544),
            .in1(N__23677),
            .in2(_gnd_net_),
            .in3(N__21922),
            .lcout(\VPP_VDDQ.countZ0Z_6 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_6 ),
            .clk(N__32755),
            .ce(),
            .sr(N__21997));
    defparam \VPP_VDDQ.count_7_LC_7_14_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_7_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_7_LC_7_14_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_7_LC_7_14_7  (
            .in0(N__27536),
            .in1(N__23473),
            .in2(_gnd_net_),
            .in3(N__21919),
            .lcout(\VPP_VDDQ.countZ0Z_7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_7 ),
            .clk(N__32755),
            .ce(),
            .sr(N__21997));
    defparam \VPP_VDDQ.count_8_LC_7_15_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_8_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_8_LC_7_15_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_8_LC_7_15_0  (
            .in0(N__27540),
            .in1(N__23181),
            .in2(_gnd_net_),
            .in3(N__21916),
            .lcout(\VPP_VDDQ.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_8 ),
            .clk(N__32753),
            .ce(),
            .sr(N__21986));
    defparam \VPP_VDDQ.count_9_LC_7_15_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_9_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_9_LC_7_15_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_9_LC_7_15_1  (
            .in0(N__27532),
            .in1(N__23206),
            .in2(_gnd_net_),
            .in3(N__21913),
            .lcout(\VPP_VDDQ.countZ0Z_9 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_8 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_9 ),
            .clk(N__32753),
            .ce(),
            .sr(N__21986));
    defparam \VPP_VDDQ.count_10_LC_7_15_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_10_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_10_LC_7_15_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_10_LC_7_15_2  (
            .in0(N__27537),
            .in1(N__23652),
            .in2(_gnd_net_),
            .in3(N__21910),
            .lcout(\VPP_VDDQ.countZ0Z_10 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_10 ),
            .clk(N__32753),
            .ce(),
            .sr(N__21986));
    defparam \VPP_VDDQ.count_11_LC_7_15_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_11_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_11_LC_7_15_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_11_LC_7_15_3  (
            .in0(N__27530),
            .in1(N__23164),
            .in2(_gnd_net_),
            .in3(N__21907),
            .lcout(\VPP_VDDQ.countZ0Z_11 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_11 ),
            .clk(N__32753),
            .ce(),
            .sr(N__21986));
    defparam \VPP_VDDQ.count_12_LC_7_15_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_12_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_12_LC_7_15_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_12_LC_7_15_4  (
            .in0(N__27538),
            .in1(N__23245),
            .in2(_gnd_net_),
            .in3(N__21904),
            .lcout(\VPP_VDDQ.countZ0Z_12 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_12 ),
            .clk(N__32753),
            .ce(),
            .sr(N__21986));
    defparam \VPP_VDDQ.count_13_LC_7_15_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_13_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_13_LC_7_15_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_13_LC_7_15_5  (
            .in0(N__27531),
            .in1(N__23272),
            .in2(_gnd_net_),
            .in3(N__22018),
            .lcout(\VPP_VDDQ.countZ0Z_13 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_13 ),
            .clk(N__32753),
            .ce(),
            .sr(N__21986));
    defparam \VPP_VDDQ.count_14_LC_7_15_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_14_LC_7_15_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_14_LC_7_15_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_14_LC_7_15_6  (
            .in0(N__27539),
            .in1(N__23284),
            .in2(_gnd_net_),
            .in3(N__22015),
            .lcout(\VPP_VDDQ.countZ0Z_14 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14 ),
            .clk(N__32753),
            .ce(),
            .sr(N__21986));
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_7_15_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_7_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(N__27244),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_14 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_15_LC_7_16_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_15_LC_7_16_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_esr_15_LC_7_16_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \VPP_VDDQ.count_esr_15_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__23259),
            .in2(_gnd_net_),
            .in3(N__22012),
            .lcout(\VPP_VDDQ.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32870),
            .ce(N__22009),
            .sr(N__21993));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_8_1_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_8_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_8_1_0  (
            .in0(_gnd_net_),
            .in1(N__21963),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_1_0_),
            .carryout(\POWERLED.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_8_1_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_8_1_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_8_1_1  (
            .in0(_gnd_net_),
            .in1(N__21946),
            .in2(N__22218),
            .in3(N__21940),
            .lcout(\POWERLED.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_8_1_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_8_1_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_8_1_2  (
            .in0(_gnd_net_),
            .in1(N__22214),
            .in2(N__23569),
            .in3(N__21937),
            .lcout(\POWERLED.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_8_1_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_8_1_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_8_1_3  (
            .in0(_gnd_net_),
            .in1(N__23557),
            .in2(N__23841),
            .in3(N__21934),
            .lcout(\POWERLED.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_8_1_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_8_1_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_8_1_4  (
            .in0(_gnd_net_),
            .in1(N__23837),
            .in2(N__23548),
            .in3(N__21931),
            .lcout(\POWERLED.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_8_1_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_8_1_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_8_1_5  (
            .in0(N__22048),
            .in1(N__23536),
            .in2(N__22219),
            .in3(N__22111),
            .lcout(\POWERLED.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_8_1_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_8_1_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_8_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23527),
            .in3(N__22108),
            .lcout(\POWERLED.mult1_un89_sum_s_8 ),
            .ltout(\POWERLED.mult1_un89_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_8_1_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_8_1_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_8_1_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_8_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22105),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_8_2_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_8_2_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_8_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_8_2_0  (
            .in0(_gnd_net_),
            .in1(N__22101),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(\POWERLED.mult1_un96_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_8_2_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_8_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(N__22084),
            .in2(N__22251),
            .in3(N__22078),
            .lcout(\POWERLED.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_8_2_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_8_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_8_2_2  (
            .in0(_gnd_net_),
            .in1(N__22247),
            .in2(N__22075),
            .in3(N__22066),
            .lcout(\POWERLED.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_8_2_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_8_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_8_2_3  (
            .in0(_gnd_net_),
            .in1(N__22063),
            .in2(N__22054),
            .in3(N__22057),
            .lcout(\POWERLED.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_8_2_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_8_2_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_8_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_8_2_4  (
            .in0(_gnd_net_),
            .in1(N__22052),
            .in2(N__22030),
            .in3(N__22021),
            .lcout(\POWERLED.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_8_2_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_8_2_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_8_2_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_8_2_5  (
            .in0(N__22469),
            .in1(N__22258),
            .in2(N__22252),
            .in3(N__22234),
            .lcout(\POWERLED.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_8_2_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_8_2_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_8_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22231),
            .in3(N__22222),
            .lcout(\POWERLED.mult1_un96_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_8_2_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_8_2_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_8_2_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_8_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23832),
            .lcout(\POWERLED.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_8_3_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_8_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__22200),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\POWERLED.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_8_3_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_8_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(N__22186),
            .in2(N__22443),
            .in3(N__22168),
            .lcout(\POWERLED.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_8_3_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_8_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_8_3_2  (
            .in0(_gnd_net_),
            .in1(N__22439),
            .in2(N__22165),
            .in3(N__22150),
            .lcout(\POWERLED.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_8_3_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_8_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(N__22465),
            .in2(N__22147),
            .in3(N__22129),
            .lcout(\POWERLED.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_8_3_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_8_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_8_3_4  (
            .in0(_gnd_net_),
            .in1(N__22126),
            .in2(N__22471),
            .in3(N__22114),
            .lcout(\POWERLED.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_8_3_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_8_3_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_8_3_5  (
            .in0(N__22493),
            .in1(N__22528),
            .in2(N__22444),
            .in3(N__22513),
            .lcout(\POWERLED.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_8_3_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_8_3_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_8_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22510),
            .in3(N__22501),
            .lcout(\POWERLED.mult1_un103_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_3_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_3_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22464),
            .lcout(\POWERLED.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_0_LC_8_4_0 .C_ON=1'b0;
    defparam \POWERLED.curr_state_0_LC_8_4_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.curr_state_0_LC_8_4_0 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \POWERLED.curr_state_0_LC_8_4_0  (
            .in0(_gnd_net_),
            .in1(N__22425),
            .in2(N__22393),
            .in3(N__22360),
            .lcout(\POWERLED.curr_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32714),
            .ce(N__32289),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_8_4_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_8_4_1 .LUT_INIT=16'b1111000010100101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_8_4_1  (
            .in0(N__22281),
            .in1(_gnd_net_),
            .in2(N__22321),
            .in3(N__22300),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_4_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_4_3 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22282),
            .in3(N__22299),
            .lcout(\POWERLED.mult1_un47_sum_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_8_4_4 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_8_4_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_8_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22277),
            .lcout(\POWERLED.un1_dutycycle_53_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIPM861_8_LC_8_4_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIPM861_8_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIPM861_8_LC_8_4_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \VPP_VDDQ.count_2_RNIPM861_8_LC_8_4_5  (
            .in0(_gnd_net_),
            .in1(N__31985),
            .in2(N__23095),
            .in3(N__23080),
            .lcout(\VPP_VDDQ.count_2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_7_LC_8_4_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_7_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_7_LC_8_4_6 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_7_LC_8_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24100),
            .in3(N__29128),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_1_LC_8_5_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_1_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_1_LC_8_5_0 .LUT_INIT=16'b1111010100001010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_1_LC_8_5_0  (
            .in0(N__31537),
            .in1(N__26426),
            .in2(N__29285),
            .in3(N__30870),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_3_LC_8_5_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_8_5_1 .LUT_INIT=16'b0001001100110111;
    LogicCell40 \POWERLED.dutycycle_RNI_5_3_LC_8_5_1  (
            .in0(N__28964),
            .in1(N__29245),
            .in2(N__29153),
            .in3(N__29675),
            .lcout(\POWERLED.g0_1_1 ),
            .ltout(\POWERLED.g0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_7_LC_8_5_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_7_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_7_LC_8_5_2 .LUT_INIT=16'b1100111000001000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_7_LC_8_5_2  (
            .in0(N__29829),
            .in1(N__29122),
            .in2(N__22585),
            .in3(N__31343),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_3_LC_8_5_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_8_5_3 .LUT_INIT=16'b1101101100100100;
    LogicCell40 \POWERLED.dutycycle_RNI_3_3_LC_8_5_3  (
            .in0(N__28965),
            .in1(N__29249),
            .in2(N__29154),
            .in3(N__29676),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_LC_8_5_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_LC_8_5_4 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_LC_8_5_4  (
            .in0(N__29830),
            .in1(N__29123),
            .in2(N__22573),
            .in3(N__31344),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNIZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_7_LC_8_5_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_7_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_7_LC_8_5_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.dutycycle_RNI_9_7_LC_8_5_5  (
            .in0(N__27871),
            .in1(_gnd_net_),
            .in2(N__22564),
            .in3(N__22561),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_9Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_LC_8_5_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_LC_8_5_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNI_11_LC_8_5_6  (
            .in0(N__29677),
            .in1(N__30158),
            .in2(N__22555),
            .in3(N__29127),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_13_LC_8_5_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_8_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_13_LC_8_5_7  (
            .in0(N__26097),
            .in1(N__29831),
            .in2(N__30018),
            .in3(N__27775),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_12_LC_8_6_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_8_6_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_12_LC_8_6_0  (
            .in0(N__29752),
            .in1(N__29484),
            .in2(N__29674),
            .in3(N__22645),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_4_LC_8_6_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_4_LC_8_6_3 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_4_LC_8_6_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \POWERLED.dutycycle_4_LC_8_6_3  (
            .in0(N__24286),
            .in1(N__31079),
            .in2(N__22639),
            .in3(N__22624),
            .lcout(\POWERLED.dutycycleZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32715),
            .ce(),
            .sr(N__26641));
    defparam \POWERLED.dutycycle_RNI_5_4_LC_8_6_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_4_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_4_LC_8_6_4 .LUT_INIT=16'b0000001100111111;
    LogicCell40 \POWERLED.dutycycle_RNI_5_4_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__29256),
            .in2(N__29815),
            .in3(N__31322),
            .lcout(),
            .ltout(\POWERLED.N_9_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_7_LC_8_6_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_7_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_7_LC_8_6_5 .LUT_INIT=16'b1100111010001100;
    LogicCell40 \POWERLED.dutycycle_RNI_1_7_LC_8_6_5  (
            .in0(N__31323),
            .in1(N__29103),
            .in2(N__22648),
            .in3(N__29648),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIVM194_4_LC_8_6_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIVM194_4_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIVM194_4_LC_8_6_6 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \POWERLED.dutycycle_RNIVM194_4_LC_8_6_6  (
            .in0(N__22635),
            .in1(N__22623),
            .in2(N__31109),
            .in3(N__24285),
            .lcout(\POWERLED.dutycycleZ0Z_8 ),
            .ltout(\POWERLED.dutycycleZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_4_LC_8_6_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_4_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_4_LC_8_6_7 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \POWERLED.dutycycle_RNI_1_4_LC_8_6_7  (
            .in0(N__29079),
            .in1(N__29748),
            .in2(N__22612),
            .in3(N__29647),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_4_LC_8_7_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_4_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_4_LC_8_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.dutycycle_RNI_7_4_LC_8_7_0  (
            .in0(N__29075),
            .in1(N__30149),
            .in2(N__29885),
            .in3(N__29257),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_7Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_4_LC_8_7_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_4_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_4_LC_8_7_1 .LUT_INIT=16'b0011011000110011;
    LogicCell40 \POWERLED.dutycycle_RNI_8_4_LC_8_7_1  (
            .in0(N__22717),
            .in1(N__22699),
            .in2(N__22609),
            .in3(N__26188),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_15_LC_8_7_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_8_7_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_15_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22606),
            .in3(N__28639),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_15_LC_8_7_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_15_LC_8_7_3 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_15_LC_8_7_3 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \POWERLED.dutycycle_15_LC_8_7_3  (
            .in0(N__22711),
            .in1(N__24421),
            .in2(N__28107),
            .in3(N__28384),
            .lcout(\POWERLED.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32716),
            .ce(),
            .sr(N__26602));
    defparam \POWERLED.dutycycle_RNI_8_10_LC_8_7_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_10_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_10_LC_8_7_4 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \POWERLED.dutycycle_RNI_8_10_LC_8_7_4  (
            .in0(N__29074),
            .in1(_gnd_net_),
            .in2(N__29683),
            .in3(N__30006),
            .lcout(\POWERLED.dutycycle_RNI_8Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIDB0M4_15_LC_8_7_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIDB0M4_15_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIDB0M4_15_LC_8_7_5 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.dutycycle_RNIDB0M4_15_LC_8_7_5  (
            .in0(N__22710),
            .in1(N__28383),
            .in2(N__28106),
            .in3(N__24420),
            .lcout(\POWERLED.dutycycleZ0Z_12 ),
            .ltout(\POWERLED.dutycycleZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_15_LC_8_7_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_15_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_15_LC_8_7_6 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \POWERLED.dutycycle_RNI_15_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(N__29478),
            .in2(N__22702),
            .in3(N__30148),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_12_LC_8_7_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_12_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_12_LC_8_7_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.dutycycle_RNI_12_LC_8_7_7  (
            .in0(N__29479),
            .in1(N__30153),
            .in2(N__30017),
            .in3(N__29681),
            .lcout(\POWERLED.m69_0_o2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_LC_8_8_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_LC_8_8_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_1_LC_8_8_0 .LUT_INIT=16'b0111111101000000;
    LogicCell40 \POWERLED.dutycycle_1_LC_8_8_0  (
            .in0(N__22681),
            .in1(N__22657),
            .in2(N__28169),
            .in3(N__22675),
            .lcout(\POWERLED.dutycycleZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32942),
            .ce(),
            .sr(N__26648));
    defparam \POWERLED.func_state_RNI2O4A1_0_LC_8_8_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2O4A1_0_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2O4A1_0_LC_8_8_1 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \POWERLED.func_state_RNI2O4A1_0_LC_8_8_1  (
            .in0(N__22895),
            .in1(N__24798),
            .in2(N__31471),
            .in3(N__28784),
            .lcout(\POWERLED.N_81 ),
            .ltout(\POWERLED.N_81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIG11I4_0_LC_8_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIG11I4_0_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIG11I4_0_LC_8_8_2 .LUT_INIT=16'b0010111010101010;
    LogicCell40 \POWERLED.dutycycle_RNIG11I4_0_LC_8_8_2  (
            .in0(N__22776),
            .in1(N__28067),
            .in2(N__22684),
            .in3(N__22792),
            .lcout(\POWERLED.dutycycleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_8_8_3 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_8_8_3 .LUT_INIT=16'b1110110011101111;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_8_8_3  (
            .in0(N__22894),
            .in1(N__24797),
            .in2(N__28829),
            .in3(N__24148),
            .lcout(\POWERLED.N_85 ),
            .ltout(\POWERLED.N_85_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKCVI4_1_LC_8_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKCVI4_1_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKCVI4_1_LC_8_8_4 .LUT_INIT=16'b0010111010101010;
    LogicCell40 \POWERLED.dutycycle_RNIKCVI4_1_LC_8_8_4  (
            .in0(N__22674),
            .in1(N__28068),
            .in2(N__22663),
            .in3(N__22656),
            .lcout(\POWERLED.dutycycle ),
            .ltout(\POWERLED.dutycycle_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIVRVA2_1_LC_8_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIVRVA2_1_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIVRVA2_1_LC_8_8_5 .LUT_INIT=16'b1111111101010100;
    LogicCell40 \POWERLED.dutycycle_RNIVRVA2_1_LC_8_8_5  (
            .in0(N__24655),
            .in1(N__24966),
            .in2(N__22660),
            .in3(N__28563),
            .lcout(\POWERLED.dutycycle_eena_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIVRVA2_0_LC_8_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIVRVA2_0_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIVRVA2_0_LC_8_8_6 .LUT_INIT=16'b1111000011111110;
    LogicCell40 \POWERLED.dutycycle_RNIVRVA2_0_LC_8_8_6  (
            .in0(N__31459),
            .in1(N__24976),
            .in2(N__28587),
            .in3(N__24654),
            .lcout(\POWERLED.dutycycle_eena ),
            .ltout(\POWERLED.dutycycle_eena_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_0_LC_8_8_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_0_LC_8_8_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_0_LC_8_8_7 .LUT_INIT=16'b0010101011101010;
    LogicCell40 \POWERLED.dutycycle_0_LC_8_8_7  (
            .in0(N__22777),
            .in1(N__28143),
            .in2(N__22786),
            .in3(N__22783),
            .lcout(\POWERLED.dutycycleZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32942),
            .ce(),
            .sr(N__26648));
    defparam \POWERLED.func_state_RNI99TE_1_LC_8_9_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI99TE_1_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI99TE_1_LC_8_9_0 .LUT_INIT=16'b0000000010111111;
    LogicCell40 \POWERLED.func_state_RNI99TE_1_LC_8_9_0  (
            .in0(N__28757),
            .in1(N__30555),
            .in2(N__25145),
            .in3(N__31288),
            .lcout(),
            .ltout(\POWERLED.N_441_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIHCGC2_1_LC_8_9_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIHCGC2_1_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIHCGC2_1_LC_8_9_1 .LUT_INIT=16'b1100110011001101;
    LogicCell40 \POWERLED.func_state_RNIHCGC2_1_LC_8_9_1  (
            .in0(N__22726),
            .in1(N__28565),
            .in2(N__22765),
            .in3(N__28457),
            .lcout(\POWERLED.dutycycle_eena_13 ),
            .ltout(\POWERLED.dutycycle_eena_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKVA67_6_LC_8_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKVA67_6_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKVA67_6_LC_8_9_2 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.dutycycle_RNIKVA67_6_LC_8_9_2  (
            .in0(N__28039),
            .in1(N__22750),
            .in2(N__22732),
            .in3(N__24336),
            .lcout(\POWERLED.dutycycleZ1Z_6 ),
            .ltout(\POWERLED.dutycycleZ1Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI88TE_1_LC_8_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI88TE_1_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI88TE_1_LC_8_9_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.func_state_RNI88TE_1_LC_8_9_3  (
            .in0(N__30373),
            .in1(N__25132),
            .in2(N__22729),
            .in3(N__28756),
            .lcout(\POWERLED.N_442 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_2_LC_8_9_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_2_LC_8_9_4 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_2_LC_8_9_4 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \POWERLED.dutycycle_2_LC_8_9_4  (
            .in0(N__22912),
            .in1(N__22921),
            .in2(_gnd_net_),
            .in3(N__24375),
            .lcout(\POWERLED.dutycycleZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32931),
            .ce(),
            .sr(N__26651));
    defparam \POWERLED.dutycycle_RNI88TE_2_LC_8_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI88TE_2_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI88TE_2_LC_8_9_5 .LUT_INIT=16'b0000100010000000;
    LogicCell40 \POWERLED.dutycycle_RNI88TE_2_LC_8_9_5  (
            .in0(N__30372),
            .in1(N__25136),
            .in2(N__26419),
            .in3(N__28758),
            .lcout(),
            .ltout(\POWERLED.N_429_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI9NTJ2_2_LC_8_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI9NTJ2_2_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI9NTJ2_2_LC_8_9_6 .LUT_INIT=16'b1010101100000000;
    LogicCell40 \POWERLED.dutycycle_RNI9NTJ2_2_LC_8_9_6  (
            .in0(N__28564),
            .in1(N__24653),
            .in2(N__22720),
            .in3(N__28030),
            .lcout(\POWERLED.dutycycle_RNI9NTJ2Z0Z_2 ),
            .ltout(\POWERLED.dutycycle_RNI9NTJ2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNINBHJ5_2_LC_8_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNINBHJ5_2_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNINBHJ5_2_LC_8_9_7 .LUT_INIT=16'b0101111101010000;
    LogicCell40 \POWERLED.dutycycle_RNINBHJ5_2_LC_8_9_7  (
            .in0(N__24376),
            .in1(_gnd_net_),
            .in2(N__22915),
            .in3(N__22911),
            .lcout(dutycycle_RNINBHJ5_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_5_LC_8_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_5_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_5_LC_8_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_2_5_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30829),
            .lcout(N_2145_i),
            .ltout(N_2145_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_6_LC_8_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_6_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_6_LC_8_10_1 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_6_LC_8_10_1  (
            .in0(N__31290),
            .in1(_gnd_net_),
            .in2(N__22903),
            .in3(N__26802),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_6 ),
            .ltout(\POWERLED.dutycycle_RNI_3Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_0_LC_8_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_0_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_0_LC_8_10_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.func_state_RNI_0_0_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22900),
            .in3(N__22889),
            .lcout(\POWERLED.func_state_RNI_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_5_LC_8_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_5_LC_8_10_3 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_5_LC_8_10_3 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.dutycycle_5_LC_8_10_3  (
            .in0(N__22816),
            .in1(N__22810),
            .in2(N__28105),
            .in3(N__24316),
            .lcout(\POWERLED.dutycycle_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32839),
            .ce(),
            .sr(N__26633));
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIB7P1F_LC_8_10_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIB7P1F_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIB7P1F_LC_8_10_4 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_fast_RNIB7P1F_LC_8_10_4  (
            .in0(N__24637),
            .in1(N__22822),
            .in2(N__22936),
            .in3(N__30781),
            .lcout(POWERLED_dutycycle_eena_14_0),
            .ltout(POWERLED_dutycycle_eena_14_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKBMSJ_5_LC_8_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKBMSJ_5_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKBMSJ_5_LC_8_10_5 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \POWERLED.dutycycle_RNIKBMSJ_5_LC_8_10_5  (
            .in0(N__22809),
            .in1(N__24315),
            .in2(N__22798),
            .in3(N__28011),
            .lcout(dutycycle_RNIKBMSJ_0_5),
            .ltout(dutycycle_RNIKBMSJ_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_5_LC_8_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_5_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_5_LC_8_10_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_5_LC_8_10_6  (
            .in0(N__26343),
            .in1(_gnd_net_),
            .in2(N__22795),
            .in3(N__31289),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_5 ),
            .ltout(\POWERLED.dutycycle_RNI_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_5_0_LC_8_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_5_0_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_5_0_LC_8_10_7 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \POWERLED.func_state_RNI_5_0_LC_8_10_7  (
            .in0(N__31891),
            .in1(N__23057),
            .in2(N__23041),
            .in3(N__24741),
            .lcout(\POWERLED.func_state_RNI_5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.slp_s3n_signal_i_0_o3_2_LC_8_11_0 .C_ON=1'b0;
    defparam \POWERLED.slp_s3n_signal_i_0_o3_2_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.slp_s3n_signal_i_0_o3_2_LC_8_11_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \POWERLED.slp_s3n_signal_i_0_o3_2_LC_8_11_0  (
            .in0(N__30367),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26924),
            .lcout(v5s_enn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_i_i_o3_0_LC_8_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_i_i_o3_0_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_i_i_o3_0_LC_8_11_1 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_i_i_o3_0_LC_8_11_1  (
            .in0(N__26925),
            .in1(N__30548),
            .in2(_gnd_net_),
            .in3(N__30365),
            .lcout(\POWERLED.N_258 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_clk_100khz_52_and_i_0_a3_0_LC_8_11_2 .C_ON=1'b0;
    defparam \POWERLED.un1_clk_100khz_52_and_i_0_a3_0_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_clk_100khz_52_and_i_0_a3_0_LC_8_11_2 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \POWERLED.un1_clk_100khz_52_and_i_0_a3_0_LC_8_11_2  (
            .in0(N__30550),
            .in1(_gnd_net_),
            .in2(N__30387),
            .in3(N__25099),
            .lcout(\POWERLED.N_443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI56A8_0_LC_8_11_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI56A8_0_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI56A8_0_LC_8_11_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.func_state_RNI56A8_0_LC_8_11_3  (
            .in0(N__23016),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31884),
            .lcout(\POWERLED.func_state_RNI56A8Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_eena_5_0_s_tz_1_LC_8_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_eena_5_0_s_tz_1_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_eena_5_0_s_tz_1_LC_8_11_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \POWERLED.dutycycle_eena_5_0_s_tz_1_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__30549),
            .in2(_gnd_net_),
            .in3(N__31786),
            .lcout(),
            .ltout(\POWERLED.dutycycle_eena_5_0_s_tzZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_eena_5_0_s_tz_LC_8_11_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_eena_5_0_s_tz_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_eena_5_0_s_tz_LC_8_11_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.dutycycle_eena_5_0_s_tz_LC_8_11_6  (
            .in0(N__30366),
            .in1(N__23015),
            .in2(N__22993),
            .in3(N__31148),
            .lcout(POWERLED_func_state_0_sqmuxa),
            .ltout(POWERLED_func_state_0_sqmuxa_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIARN73_1_LC_8_11_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIARN73_1_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIARN73_1_LC_8_11_7 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \POWERLED.func_state_RNIARN73_1_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__22960),
            .in2(N__22939),
            .in3(N__24688),
            .lcout(N_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_8_12_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_8_12_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_8_12_0  (
            .in0(N__33287),
            .in1(N__33613),
            .in2(N__33521),
            .in3(N__25020),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIHA461_4_LC_8_12_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIHA461_4_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIHA461_4_LC_8_12_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIHA461_4_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__23110),
            .in2(N__22924),
            .in3(N__32009),
            .lcout(\VPP_VDDQ.count_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_4_LC_8_12_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_4_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_4_LC_8_12_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.count_2_4_LC_8_12_2  (
            .in0(N__33290),
            .in1(N__25021),
            .in2(N__33522),
            .in3(N__33622),
            .lcout(\VPP_VDDQ.count_2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32994),
            .ce(N__32059),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_5_LC_8_12_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_5_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_5_LC_8_12_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.count_2_5_LC_8_12_3  (
            .in0(N__33511),
            .in1(N__33294),
            .in2(N__33677),
            .in3(N__25380),
            .lcout(\VPP_VDDQ.count_2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32994),
            .ce(N__32059),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_8_12_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_8_12_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_8_12_4  (
            .in0(N__33288),
            .in1(N__33614),
            .in2(N__25381),
            .in3(N__33509),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIJD561_5_LC_8_12_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIJD561_5_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIJD561_5_LC_8_12_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNIJD561_5_LC_8_12_5  (
            .in0(N__23104),
            .in1(_gnd_net_),
            .in2(N__23098),
            .in3(N__32010),
            .lcout(\VPP_VDDQ.count_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_8_LC_8_12_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_8_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_8_LC_8_12_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.count_2_8_LC_8_12_6  (
            .in0(N__25330),
            .in1(N__33618),
            .in2(N__33301),
            .in3(N__33512),
            .lcout(\VPP_VDDQ.count_2_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32994),
            .ce(N__32059),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_8_12_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_8_12_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_8_12_7  (
            .in0(N__33510),
            .in1(N__25329),
            .in2(N__33676),
            .in3(N__33289),
            .lcout(\VPP_VDDQ.count_2_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_2_LC_8_13_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_2_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_2_LC_8_13_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.count_2_2_LC_8_13_0  (
            .in0(N__33284),
            .in1(N__25050),
            .in2(N__33518),
            .in3(N__33609),
            .lcout(\VPP_VDDQ.count_2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32999),
            .ce(N__32074),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_8_13_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_8_13_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_8_13_1  (
            .in0(N__33606),
            .in1(N__33481),
            .in2(N__25051),
            .in3(N__33282),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNID4261_2_LC_8_13_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNID4261_2_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNID4261_2_LC_8_13_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNID4261_2_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__23068),
            .in2(N__23062),
            .in3(N__32008),
            .lcout(\VPP_VDDQ.count_2Z0Z_2 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_2_LC_8_13_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_2_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_2_LC_8_13_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNI_2_LC_8_13_3  (
            .in0(N__27679),
            .in1(N__25393),
            .in2(N__23146),
            .in3(N__25354),
            .lcout(\VPP_VDDQ.un9_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_15_LC_8_13_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_15_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_15_LC_8_13_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.count_2_15_LC_8_13_4  (
            .in0(N__33283),
            .in1(N__33608),
            .in2(N__33517),
            .in3(N__25488),
            .lcout(\VPP_VDDQ.count_2_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32999),
            .ce(N__32074),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_8_13_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_8_13_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_8_13_5  (
            .in0(N__25489),
            .in1(N__33488),
            .in2(N__33675),
            .in3(N__33286),
            .lcout(),
            .ltout(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIL79C1_15_LC_8_13_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIL79C1_15_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIL79C1_15_LC_8_13_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \VPP_VDDQ.count_2_RNIL79C1_15_LC_8_13_6  (
            .in0(N__32075),
            .in1(_gnd_net_),
            .in2(N__23143),
            .in3(N__23140),
            .lcout(\VPP_VDDQ.count_2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_3_LC_8_13_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_3_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_3_LC_8_13_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.count_2_3_LC_8_13_7  (
            .in0(N__33607),
            .in1(N__33285),
            .in2(N__33523),
            .in3(N__27711),
            .lcout(\VPP_VDDQ.count_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32999),
            .ce(N__32074),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_8_14_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_8_14_0 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_LC_8_14_0  (
            .in0(N__27529),
            .in1(N__23134),
            .in2(N__23395),
            .in3(N__23305),
            .lcout(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32941),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_8_14_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_8_14_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_8_14_1  (
            .in0(N__23457),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23421),
            .lcout(\VPP_VDDQ.N_551 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_8_14_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_8_14_2 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_8_14_2  (
            .in0(N__23386),
            .in1(N__23431),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vpp_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_8_14_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_8_14_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_8_14_3  (
            .in0(N__33513),
            .in1(N__25749),
            .in2(N__33722),
            .in3(N__33295),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIJ48C1_14_LC_8_14_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIJ48C1_14_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIJ48C1_14_LC_8_14_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIJ48C1_14_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__25738),
            .in2(N__23113),
            .in3(N__32016),
            .lcout(\VPP_VDDQ.count_2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_8_14_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_8_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_RNIVJP51_3_LC_8_14_5  (
            .in0(N__23511),
            .in1(N__23499),
            .in2(N__23488),
            .in3(N__23472),
            .lcout(\VPP_VDDQ.un6_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNILLP51_1_LC_8_14_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNILLP51_1_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNILLP51_1_LC_8_14_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \VPP_VDDQ.curr_state_RNILLP51_1_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__23456),
            .in2(_gnd_net_),
            .in3(N__23304),
            .lcout(N_325),
            .ltout(N_325_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_8_14_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_8_14_7 .LUT_INIT=16'b0011100010101010;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_8_14_7  (
            .in0(N__23430),
            .in1(N__23422),
            .in2(N__23398),
            .in3(N__27528),
            .lcout(\VPP_VDDQ.delayed_vddq_pwrgd_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_0_sqmuxa_0_a2_LC_8_15_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_0_sqmuxa_0_a2_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_0_sqmuxa_0_a2_LC_8_15_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_0_sqmuxa_0_a2_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__33122),
            .in2(_gnd_net_),
            .in3(N__23385),
            .lcout(\VPP_VDDQ.N_541 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_8_15_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_8_15_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_esr_RNI7CQO_15_LC_8_15_2  (
            .in0(N__23283),
            .in1(N__23271),
            .in2(N__23260),
            .in3(N__23244),
            .lcout(),
            .ltout(\VPP_VDDQ.un6_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_8_15_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_8_15_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_esr_RNIRFM64_15_LC_8_15_3  (
            .in0(N__23233),
            .in1(N__23152),
            .in2(N__23224),
            .in3(N__23626),
            .lcout(\VPP_VDDQ.un6_count ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_8_15_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_8_15_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \VPP_VDDQ.count_RNIFC141_11_LC_8_15_4  (
            .in0(N__23205),
            .in1(N__23193),
            .in2(N__23182),
            .in3(N__23163),
            .lcout(\VPP_VDDQ.un6_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI63141_10_LC_8_15_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_8_15_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_RNI63141_10_LC_8_15_5  (
            .in0(N__23676),
            .in1(N__23664),
            .in2(N__23653),
            .in3(N__23637),
            .lcout(\VPP_VDDQ.un6_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PRIMARY_VOLTAGES_EN.N_171_i_LC_8_15_7 .C_ON=1'b0;
    defparam \PRIMARY_VOLTAGES_EN.N_171_i_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \PRIMARY_VOLTAGES_EN.N_171_i_LC_8_15_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \PRIMARY_VOLTAGES_EN.N_171_i_LC_8_15_7  (
            .in0(N__24860),
            .in1(N__24837),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(v1p8a_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_9_1_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_9_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_9_1_0  (
            .in0(_gnd_net_),
            .in1(N__23605),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_1_0_),
            .carryout(\POWERLED.mult1_un82_sum_cry_2_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_9_1_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_9_1_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_9_1_1  (
            .in0(_gnd_net_),
            .in1(N__23581),
            .in2(N__23922),
            .in3(N__23560),
            .lcout(\POWERLED.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_2_c ),
            .carryout(\POWERLED.mult1_un82_sum_cry_3_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_9_1_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_9_1_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_9_1_2  (
            .in0(_gnd_net_),
            .in1(N__23918),
            .in2(N__23779),
            .in3(N__23551),
            .lcout(\POWERLED.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_3_c ),
            .carryout(\POWERLED.mult1_un82_sum_cry_4_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_9_1_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_9_1_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_9_1_3  (
            .in0(_gnd_net_),
            .in1(N__23767),
            .in2(N__23703),
            .in3(N__23539),
            .lcout(\POWERLED.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_4_c ),
            .carryout(\POWERLED.mult1_un82_sum_cry_5_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_9_1_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_9_1_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_9_1_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_9_1_4  (
            .in0(_gnd_net_),
            .in1(N__23699),
            .in2(N__23758),
            .in3(N__23530),
            .lcout(\POWERLED.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_5_c ),
            .carryout(\POWERLED.mult1_un82_sum_cry_6_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_9_1_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_9_1_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_9_1_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_9_1_5  (
            .in0(N__23833),
            .in1(N__23746),
            .in2(N__23923),
            .in3(N__23518),
            .lcout(\POWERLED.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_6_c ),
            .carryout(\POWERLED.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_9_1_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_9_1_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_9_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23719),
            .in3(N__23515),
            .lcout(\POWERLED.mult1_un82_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_9_1_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_9_1_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_9_1_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_9_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25618),
            .lcout(\POWERLED.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_2_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_2_0  (
            .in0(_gnd_net_),
            .in1(N__23808),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_2_0_),
            .carryout(\POWERLED.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_9_2_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_9_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_9_2_1  (
            .in0(_gnd_net_),
            .in1(N__23791),
            .in2(N__23736),
            .in3(N__23770),
            .lcout(\POWERLED.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_9_2_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_9_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_9_2_2  (
            .in0(_gnd_net_),
            .in1(N__23732),
            .in2(N__25693),
            .in3(N__23761),
            .lcout(\POWERLED.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_9_2_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_9_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_9_2_3  (
            .in0(_gnd_net_),
            .in1(N__25678),
            .in2(N__25624),
            .in3(N__23749),
            .lcout(\POWERLED.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_9_2_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_9_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_9_2_4  (
            .in0(_gnd_net_),
            .in1(N__25622),
            .in2(N__25666),
            .in3(N__23740),
            .lcout(\POWERLED.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_9_2_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_9_2_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_9_2_5  (
            .in0(N__23695),
            .in1(N__25651),
            .in2(N__23737),
            .in3(N__23710),
            .lcout(\POWERLED.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_9_2_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_9_2_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_9_2_6  (
            .in0(_gnd_net_),
            .in1(N__25639),
            .in2(_gnd_net_),
            .in3(N__23707),
            .lcout(\POWERLED.mult1_un75_sum_s_8 ),
            .ltout(\POWERLED.mult1_un75_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_9_2_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_9_2_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_9_2_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_9_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23926),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_3_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_3_0  (
            .in0(_gnd_net_),
            .in1(N__23905),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_3_0_),
            .carryout(\POWERLED.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_3_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_3_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23884),
            .in3(N__23872),
            .lcout(\POWERLED.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_9_3_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_9_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_9_3_2  (
            .in0(_gnd_net_),
            .in1(N__23932),
            .in2(N__23953),
            .in3(N__23869),
            .lcout(\POWERLED.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_9_3_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_9_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_9_3_3  (
            .in0(_gnd_net_),
            .in1(N__27234),
            .in2(N__24040),
            .in3(N__23866),
            .lcout(\POWERLED.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_9_3_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_9_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_9_3_4  (
            .in0(_gnd_net_),
            .in1(N__27235),
            .in2(N__24019),
            .in3(N__23863),
            .lcout(\POWERLED.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_9_3_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_9_3_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_9_3_5  (
            .in0(N__25904),
            .in1(N__23992),
            .in2(N__23854),
            .in3(N__23860),
            .lcout(\POWERLED.mult1_un61_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_9_3_6 .C_ON=1'b0;
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_9_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_9_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23857),
            .lcout(\POWERLED.mult1_un54_sum_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_3_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_3_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_3_7  (
            .in0(N__23990),
            .in1(N__23991),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_4_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24085),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_4_0_),
            .carryout(\POWERLED.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_9_4_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_9_4_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_9_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24061),
            .in3(N__24052),
            .lcout(\POWERLED.mult1_un47_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_9_4_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_9_4_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_9_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24049),
            .in3(N__24031),
            .lcout(\POWERLED.mult1_un47_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_9_4_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_9_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_9_4_3  (
            .in0(_gnd_net_),
            .in1(N__27236),
            .in2(N__24028),
            .in3(N__24010),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_9_4_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_9_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_9_4_4  (
            .in0(_gnd_net_),
            .in1(N__27237),
            .in2(N__24007),
            .in3(N__23977),
            .lcout(\POWERLED.mult1_un47_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_9_4_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_9_4_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_9_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23974),
            .in3(N__23965),
            .lcout(\POWERLED.mult1_un54_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_9_4_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_9_4_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_9_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25807),
            .lcout(\POWERLED.mult1_un61_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_9_4_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_9_4_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_9_4_7  (
            .in0(N__23948),
            .in1(N__23949),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_9_LC_9_5_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_9_LC_9_5_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_9_LC_9_5_0 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \POWERLED.dutycycle_9_LC_9_5_0  (
            .in0(N__24130),
            .in1(N__24235),
            .in2(N__28175),
            .in3(N__24124),
            .lcout(\POWERLED.dutycycleZ1Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32818),
            .ce(),
            .sr(N__26652));
    defparam \POWERLED.dutycycle_RNIB8VL4_14_LC_9_5_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIB8VL4_14_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIB8VL4_14_LC_9_5_2 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \POWERLED.dutycycle_RNIB8VL4_14_LC_9_5_2  (
            .in0(N__26137),
            .in1(N__26172),
            .in2(N__28174),
            .in3(N__26148),
            .lcout(\POWERLED.dutycycleZ0Z_13 ),
            .ltout(\POWERLED.dutycycleZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_14_LC_9_5_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_9_5_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_14_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24136),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_2293_i ),
            .ltout(\POWERLED.N_2293_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOBHB2_0_1_LC_9_5_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOBHB2_0_1_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOBHB2_0_1_LC_9_5_4 .LUT_INIT=16'b1100110111011101;
    LogicCell40 \POWERLED.func_state_RNIOBHB2_0_1_LC_9_5_4  (
            .in0(N__28486),
            .in1(N__28590),
            .in2(N__24133),
            .in3(N__31102),
            .lcout(\POWERLED.dutycycle_eena_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOBHB2_9_LC_9_5_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOBHB2_9_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOBHB2_9_LC_9_5_5 .LUT_INIT=16'b1100110011101111;
    LogicCell40 \POWERLED.dutycycle_RNIOBHB2_9_LC_9_5_5  (
            .in0(N__29792),
            .in1(N__28589),
            .in2(N__31115),
            .in3(N__28485),
            .lcout(\POWERLED.dutycycle_eena_2 ),
            .ltout(\POWERLED.dutycycle_eena_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJDG64_9_LC_9_5_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJDG64_9_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJDG64_9_LC_9_5_6 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.dutycycle_RNIJDG64_9_LC_9_5_6  (
            .in0(N__28159),
            .in1(N__24123),
            .in2(N__24115),
            .in3(N__24234),
            .lcout(\POWERLED.dutycycleZ0Z_2 ),
            .ltout(\POWERLED.dutycycleZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_11_LC_9_5_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_9_5_7 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_11_LC_9_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24112),
            .in3(N__30157),
            .lcout(\POWERLED.un1_dutycycle_53_7_a0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_13_LC_9_6_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_13_LC_9_6_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_13_LC_9_6_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.dutycycle_13_LC_9_6_0  (
            .in0(N__24109),
            .in1(N__28141),
            .in2(N__28234),
            .in3(N__24525),
            .lcout(\POWERLED.dutycycleZ1Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32921),
            .ce(),
            .sr(N__26631));
    defparam \POWERLED.dutycycle_RNI95UL4_13_LC_9_6_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI95UL4_13_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI95UL4_13_LC_9_6_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.dutycycle_RNI95UL4_13_LC_9_6_1  (
            .in0(N__28140),
            .in1(N__24108),
            .in2(N__24526),
            .in3(N__28230),
            .lcout(\POWERLED.dutycycleZ0Z_9 ),
            .ltout(\POWERLED.dutycycleZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_13_LC_9_6_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_9_6_2 .LUT_INIT=16'b1010000000100000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_13_LC_9_6_2  (
            .in0(N__26208),
            .in1(N__24099),
            .in2(N__24214),
            .in3(N__24193),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_13 ),
            .ltout(\POWERLED.dutycycle_RNI_1Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_14_LC_9_6_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_14_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_14_LC_9_6_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_14_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24211),
            .in3(N__28329),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_7_LC_9_6_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_7_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_7_LC_9_6_4 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_7_LC_9_6_4  (
            .in0(N__31320),
            .in1(N__29102),
            .in2(N__27869),
            .in3(N__29660),
            .lcout(\POWERLED.un1_dutycycle_53_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_14_LC_9_6_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_14_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_14_LC_9_6_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_1_14_LC_9_6_5  (
            .in0(N__28643),
            .in1(N__28328),
            .in2(_gnd_net_),
            .in3(N__24187),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_LC_9_6_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_LC_9_6_6 .LUT_INIT=16'b1011001100110011;
    LogicCell40 \POWERLED.dutycycle_RNI_6_LC_9_6_6  (
            .in0(N__31321),
            .in1(N__24169),
            .in2(N__27870),
            .in3(N__29661),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_57_a0_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_13_LC_9_6_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_13_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_13_LC_9_6_7 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \POWERLED.dutycycle_RNI_3_13_LC_9_6_7  (
            .in0(N__26090),
            .in1(N__28330),
            .in2(N__24160),
            .in3(N__26209),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_1_LC_9_7_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_2_1_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_1_LC_9_7_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_1_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31464),
            .in3(N__31520),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_1 ),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_9_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_9_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__31521),
            .in2(N__24492),
            .in3(N__24142),
            .lcout(\POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__24464),
            .in2(N__26420),
            .in3(N__24139),
            .lcout(\POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(N__28943),
            .in2(N__24493),
            .in3(N__24289),
            .lcout(\POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__24468),
            .in2(N__29292),
            .in3(N__24277),
            .lcout(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__24472),
            .in2(N__30869),
            .in3(N__24274),
            .lcout(\POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_4 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI_LC_9_7_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI_LC_9_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNI_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(N__31349),
            .in2(N__24495),
            .in3(N__24271),
            .lcout(\POWERLED.un1_dutycycle_94_cry_5_c_RNIZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_7_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(N__29129),
            .in2(N__24494),
            .in3(N__24241),
            .lcout(\POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__24500),
            .in2(N__29682),
            .in3(N__24238),
            .lcout(\POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNI3B2U_LC_9_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNI3B2U_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNI3B2U_LC_9_8_1 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_8_c_RNI3B2U_LC_9_8_1  (
            .in0(N__31086),
            .in1(N__29856),
            .in2(N__24507),
            .in3(N__24223),
            .lcout(\POWERLED.un1_dutycycle_94_cry_8_c_RNI3B2UZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_8 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNI4D3U_LC_9_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNI4D3U_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNI4D3U_LC_9_8_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_9_c_RNI4D3U_LC_9_8_2  (
            .in0(N__31094),
            .in1(N__24499),
            .in2(N__30005),
            .in3(N__24220),
            .lcout(\POWERLED.un1_dutycycle_94_cry_9_c_RNI4D3UZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIC0LB1_LC_9_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIC0LB1_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIC0LB1_LC_9_8_3 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_10_c_RNIC0LB1_LC_9_8_3  (
            .in0(N__31087),
            .in1(N__24506),
            .in2(N__30160),
            .in3(N__24217),
            .lcout(\POWERLED.un1_dutycycle_94_cry_10_c_RNIC0LBZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNID2MB1_LC_9_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNID2MB1_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNID2MB1_LC_9_8_4 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_11_c_RNID2MB1_LC_9_8_4  (
            .in0(N__31096),
            .in1(N__24502),
            .in2(N__29477),
            .in3(N__24529),
            .lcout(\POWERLED.un1_dutycycle_94_cry_11_c_RNID2MBZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIE4NB1_LC_9_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIE4NB1_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIE4NB1_LC_9_8_5 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_12_c_RNIE4NB1_LC_9_8_5  (
            .in0(N__31088),
            .in1(N__26098),
            .in2(N__24508),
            .in3(N__24511),
            .lcout(\POWERLED.un1_dutycycle_94_cry_12_c_RNIE4NBZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNIF6OB1_LC_9_8_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNIF6OB1_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNIF6OB1_LC_9_8_6 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_13_c_RNIF6OB1_LC_9_8_6  (
            .in0(N__31095),
            .in1(N__24501),
            .in2(N__28355),
            .in3(N__24427),
            .lcout(\POWERLED.un1_dutycycle_94_cry_13_c_RNIF6OBZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIG8PB1_LC_9_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIG8PB1_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIG8PB1_LC_9_8_7 .LUT_INIT=16'b0001001000100001;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_14_c_RNIG8PB1_LC_9_8_7  (
            .in0(N__30768),
            .in1(N__31097),
            .in2(N__28654),
            .in3(N__24424),
            .lcout(\POWERLED.un1_dutycycle_94_cry_14_c_RNIG8PBZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2MQD_1_LC_9_9_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2MQD_1_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2MQD_1_LC_9_9_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \POWERLED.func_state_RNI2MQD_1_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__30243),
            .in2(_gnd_net_),
            .in3(N__28820),
            .lcout(),
            .ltout(\POWERLED.dutycycle_1_0_iv_i_a3_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIUO1P2_LC_9_9_3 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIUO1P2_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIUO1P2_LC_9_9_3 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNIUO1P2_LC_9_9_3  (
            .in0(N__24412),
            .in1(N__26698),
            .in2(N__24388),
            .in3(N__24385),
            .lcout(\POWERLED.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_LC_9_9_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_LC_9_9_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.dutycycle_RNI_1_LC_9_9_4  (
            .in0(N__31455),
            .in1(N__31533),
            .in2(N__30694),
            .in3(N__28951),
            .lcout(m57_i_o2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIEVTS3_LC_9_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIEVTS3_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIEVTS3_LC_9_9_6 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNIEVTS3_LC_9_9_6  (
            .in0(N__24610),
            .in1(N__28559),
            .in2(N__24355),
            .in3(N__31001),
            .lcout(\POWERLED.un1_dutycycle_94_cry_5_c_RNIEVTSZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNILH0U3_LC_9_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNILH0U3_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNILH0U3_LC_9_9_7 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNILH0U3_LC_9_9_7  (
            .in0(N__31002),
            .in1(N__24325),
            .in2(N__28586),
            .in3(N__24609),
            .lcout(\POWERLED.dutycycle_set_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_6_LC_9_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_6_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_6_LC_9_10_0 .LUT_INIT=16'b1111000011110111;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_6_LC_9_10_0  (
            .in0(N__24740),
            .in1(N__24820),
            .in2(N__24808),
            .in3(N__30683),
            .lcout(\POWERLED.dutycycle_RNI2O4A1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_5_LC_9_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_5_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_5_LC_9_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_5_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__24753),
            .in2(_gnd_net_),
            .in3(N__24739),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_5Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOGRS_0_1_LC_9_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOGRS_0_1_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOGRS_0_1_LC_9_10_2 .LUT_INIT=16'b1111111101010111;
    LogicCell40 \POWERLED.func_state_RNIOGRS_0_1_LC_9_10_2  (
            .in0(N__31892),
            .in1(N__30684),
            .in2(N__24700),
            .in3(N__31082),
            .lcout(),
            .ltout(\POWERLED.func_state_RNIOGRS_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIQ8072_1_LC_9_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIQ8072_1_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIQ8072_1_LC_9_10_3 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \POWERLED.func_state_RNIQ8072_1_LC_9_10_3  (
            .in0(N__30769),
            .in1(N__24697),
            .in2(N__24691),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIR1FD4_1_LC_9_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIR1FD4_1_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIR1FD4_1_LC_9_10_4 .LUT_INIT=16'b1010111110111011;
    LogicCell40 \POWERLED.func_state_RNIR1FD4_1_LC_9_10_4  (
            .in0(N__24683),
            .in1(N__30556),
            .in2(N__24658),
            .in3(N__24934),
            .lcout(\POWERLED.N_379_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIVRVA2_6_LC_9_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIVRVA2_6_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIVRVA2_6_LC_9_10_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \POWERLED.dutycycle_RNIVRVA2_6_LC_9_10_5  (
            .in0(N__24935),
            .in1(N__26686),
            .in2(_gnd_net_),
            .in3(N__28554),
            .lcout(G_22_i_a2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIMJCH1_1_LC_9_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIMJCH1_1_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIMJCH1_1_LC_9_10_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.func_state_RNIMJCH1_1_LC_9_10_7  (
            .in0(N__28857),
            .in1(N__31669),
            .in2(N__31164),
            .in3(N__24631),
            .lcout(\POWERLED.N_564 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_3_LC_9_11_0 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_3_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_3_LC_9_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_3_LC_9_11_0  (
            .in0(N__24601),
            .in1(N__24586),
            .in2(N__24571),
            .in3(N__24555),
            .lcout(),
            .ltout(\VCCIN_PWRGD.un10_outputZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_LC_9_11_1 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_LC_9_11_1 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_LC_9_11_1  (
            .in0(N__24954),
            .in1(_gnd_net_),
            .in2(N__24901),
            .in3(N__25240),
            .lcout(vccin_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_0_LC_9_11_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_0_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_0_LC_9_11_2 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_0_LC_9_11_2  (
            .in0(N__25184),
            .in1(N__25215),
            .in2(_gnd_net_),
            .in3(N__24886),
            .lcout(RSMRST_PWRGD_curr_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32843),
            .ce(N__27385),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNIJVRG6_1_LC_9_11_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNIJVRG6_1_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNIJVRG6_1_LC_9_11_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNIJVRG6_1_LC_9_11_3  (
            .in0(N__25179),
            .in1(N__25239),
            .in2(_gnd_net_),
            .in3(N__26883),
            .lcout(N_323),
            .ltout(N_323_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_12_LC_9_11_4 .C_ON=1'b0;
    defparam \POWERLED.G_12_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_12_LC_9_11_4 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \POWERLED.G_12_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__25212),
            .in2(N__24880),
            .in3(N__27522),
            .lcout(G_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_1_LC_9_11_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_1_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_1_LC_9_11_5 .LUT_INIT=16'b0000010001010100;
    LogicCell40 \RSMRST_PWRGD.curr_state_1_LC_9_11_5  (
            .in0(N__25216),
            .in1(N__25238),
            .in2(N__25186),
            .in3(N__26884),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32843),
            .ce(N__27385),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_9_11_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_9_11_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_9_11_6  (
            .in0(N__25237),
            .in1(N__25180),
            .in2(_gnd_net_),
            .in3(N__25214),
            .lcout(RSMRSTn_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32843),
            .ce(N__27385),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_9_11_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_9_11_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_fast_LC_9_11_7  (
            .in0(N__25213),
            .in1(N__25236),
            .in2(_gnd_net_),
            .in3(N__25185),
            .lcout(RSMRSTn_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32843),
            .ce(N__27385),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNIOAEU1_0_LC_9_12_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNIOAEU1_0_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNIOAEU1_0_LC_9_12_0 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNIOAEU1_0_LC_9_12_0  (
            .in0(N__25235),
            .in1(N__25210),
            .in2(_gnd_net_),
            .in3(N__25177),
            .lcout(\RSMRST_PWRGD.N_445_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PRIMARY_VOLTAGES_EN.un2_v1p8a_en_i_o3_LC_9_12_2 .C_ON=1'b0;
    defparam \PRIMARY_VOLTAGES_EN.un2_v1p8a_en_i_o3_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \PRIMARY_VOLTAGES_EN.un2_v1p8a_en_i_o3_LC_9_12_2 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \PRIMARY_VOLTAGES_EN.un2_v1p8a_en_i_o3_LC_9_12_2  (
            .in0(N__24870),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24838),
            .lcout(),
            .ltout(N_171_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_3_0_a2_LC_9_12_3 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_3_0_a2_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_3_0_a2_LC_9_12_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_3_0_a2_LC_9_12_3  (
            .in0(N__25293),
            .in1(N__25279),
            .in2(N__25258),
            .in3(N__25255),
            .lcout(N_283),
            .ltout(N_283_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_9_12_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_9_12_4 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__25211),
            .in2(N__25189),
            .in3(N__25178),
            .lcout(rsmrstn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32995),
            .ce(N__27389),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI38QU_6_LC_9_12_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI38QU_6_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI38QU_6_LC_9_12_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNI38QU_6_LC_9_12_5  (
            .in0(N__25428),
            .in1(N__25455),
            .in2(_gnd_net_),
            .in3(N__32050),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI38QU_0_6_LC_9_12_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI38QU_0_6_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI38QU_0_6_LC_9_12_6 .LUT_INIT=16'b0001000000010011;
    LogicCell40 \VPP_VDDQ.count_2_RNI38QU_0_6_LC_9_12_6  (
            .in0(N__25456),
            .in1(N__25033),
            .in2(N__32076),
            .in3(N__25429),
            .lcout(),
            .ltout(\VPP_VDDQ.un9_clk_100khz_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIOUR33_1_LC_9_12_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIOUR33_1_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIOUR33_1_LC_9_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIOUR33_1_LC_9_12_7  (
            .in0(N__32137),
            .in1(N__25066),
            .in2(N__25060),
            .in3(N__31585),
            .lcout(\VPP_VDDQ.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_9_13_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_9_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__32194),
            .in2(N__32170),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_9_13_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_9_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__25057),
            .in2(_gnd_net_),
            .in3(N__25039),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_9_13_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_9_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__27678),
            .in2(_gnd_net_),
            .in3(N__25036),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_9_13_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_9_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__25032),
            .in2(_gnd_net_),
            .in3(N__25012),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_9_13_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_9_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__25392),
            .in2(_gnd_net_),
            .in3(N__25369),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_9_13_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_9_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__25366),
            .in2(_gnd_net_),
            .in3(N__25360),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_9_13_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_9_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__32209),
            .in2(_gnd_net_),
            .in3(N__25357),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_9_13_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_9_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__25353),
            .in2(_gnd_net_),
            .in3(N__25321),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_9_14_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_9_14_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31638),
            .in3(N__25318),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_9_14_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_9_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__31599),
            .in2(_gnd_net_),
            .in3(N__25315),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_9_14_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_9_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__31912),
            .in2(_gnd_net_),
            .in3(N__25312),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_9_14_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_9_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__25560),
            .in2(_gnd_net_),
            .in3(N__25309),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_9_14_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_9_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__25527),
            .in2(_gnd_net_),
            .in3(N__25498),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_9_14_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_9_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__25467),
            .in2(_gnd_net_),
            .in3(N__25495),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_9_14_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_9_14_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_9_14_6  (
            .in0(N__25480),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25492),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_15_LC_9_14_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_15_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_15_LC_9_14_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_2_RNI_15_LC_9_14_7  (
            .in0(N__25528),
            .in1(N__25479),
            .in2(N__25471),
            .in3(N__25561),
            .lcout(\VPP_VDDQ.un9_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_9_15_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_9_15_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_9_15_0  (
            .in0(N__33649),
            .in1(N__33264),
            .in2(N__25444),
            .in3(N__33427),
            .lcout(\VPP_VDDQ.count_2_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_6_LC_9_15_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_6_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_6_LC_9_15_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.count_2_6_LC_9_15_1  (
            .in0(N__33268),
            .in1(N__25443),
            .in2(N__33490),
            .in3(N__33656),
            .lcout(\VPP_VDDQ.count_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33039),
            .ce(N__32089),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_9_15_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_9_15_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_9_15_2  (
            .in0(N__33650),
            .in1(N__33265),
            .in2(N__25413),
            .in3(N__33428),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIRP961_9_LC_9_15_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIRP961_9_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIRP961_9_LC_9_15_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIRP961_9_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__25399),
            .in2(N__25417),
            .in3(N__32079),
            .lcout(\VPP_VDDQ.count_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_9_LC_9_15_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_9_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_9_LC_9_15_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_9_LC_9_15_4  (
            .in0(N__33654),
            .in1(N__33269),
            .in2(N__25414),
            .in3(N__33436),
            .lcout(\VPP_VDDQ.count_2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33039),
            .ce(N__32089),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_10_LC_9_15_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_10_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_10_LC_9_15_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.count_2_10_LC_9_15_5  (
            .in0(N__33267),
            .in1(N__33655),
            .in2(N__33489),
            .in3(N__25582),
            .lcout(\VPP_VDDQ.count_2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33039),
            .ce(N__32089),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_9_15_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_9_15_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_9_15_6  (
            .in0(N__25581),
            .in1(N__33266),
            .in2(N__33705),
            .in3(N__33429),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI4TU51_10_LC_9_15_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI4TU51_10_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI4TU51_10_LC_9_15_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNI4TU51_10_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__25573),
            .in2(N__25567),
            .in3(N__32080),
            .lcout(\VPP_VDDQ.count_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_9_16_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_9_16_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_9_16_0  (
            .in0(N__25548),
            .in1(N__33491),
            .in2(N__33718),
            .in3(N__33296),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIFU5C1_12_LC_9_16_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIFU5C1_12_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIFU5C1_12_LC_9_16_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIFU5C1_12_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__32081),
            .in2(N__25564),
            .in3(N__25537),
            .lcout(\VPP_VDDQ.count_2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_12_LC_9_16_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_12_LC_9_16_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_12_LC_9_16_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.count_2_12_LC_9_16_2  (
            .in0(N__25549),
            .in1(N__33492),
            .in2(N__33720),
            .in3(N__33299),
            .lcout(\VPP_VDDQ.count_2_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33040),
            .ce(N__32073),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_9_16_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_9_16_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_9_16_4  (
            .in0(N__33493),
            .in1(N__25515),
            .in2(N__33719),
            .in3(N__33297),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIH17C1_13_LC_9_16_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIH17C1_13_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIH17C1_13_LC_9_16_5 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \VPP_VDDQ.count_2_RNIH17C1_13_LC_9_16_5  (
            .in0(N__25504),
            .in1(N__32082),
            .in2(N__25531),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_13_LC_9_16_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_13_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_13_LC_9_16_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.count_2_13_LC_9_16_6  (
            .in0(N__33494),
            .in1(N__25516),
            .in2(N__33721),
            .in3(N__33300),
            .lcout(\VPP_VDDQ.count_2_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33040),
            .ce(N__32073),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_14_LC_9_16_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_14_LC_9_16_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_14_LC_9_16_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.count_2_14_LC_9_16_7  (
            .in0(N__33298),
            .in1(N__33495),
            .in2(N__25756),
            .in3(N__33684),
            .lcout(\VPP_VDDQ.count_2_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33040),
            .ce(N__32073),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_11_2_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_11_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_11_2_0  (
            .in0(_gnd_net_),
            .in1(N__25726),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_2_0_),
            .carryout(\POWERLED.mult1_un68_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_11_2_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_11_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_11_2_1  (
            .in0(_gnd_net_),
            .in1(N__25705),
            .in2(N__25773),
            .in3(N__25681),
            .lcout(\POWERLED.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_11_2_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_11_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_11_2_2  (
            .in0(_gnd_net_),
            .in1(N__25769),
            .in2(N__25975),
            .in3(N__25669),
            .lcout(\POWERLED.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_11_2_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_11_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_11_2_3  (
            .in0(_gnd_net_),
            .in1(N__25948),
            .in2(N__25803),
            .in3(N__25654),
            .lcout(\POWERLED.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_11_2_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_11_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_11_2_4  (
            .in0(_gnd_net_),
            .in1(N__25799),
            .in2(N__25930),
            .in3(N__25642),
            .lcout(\POWERLED.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_11_2_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_11_2_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_11_2_5  (
            .in0(N__25614),
            .in1(N__25870),
            .in2(N__25774),
            .in3(N__25630),
            .lcout(\POWERLED.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_11_2_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_11_2_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_11_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25834),
            .in3(N__25627),
            .lcout(\POWERLED.mult1_un68_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_11_2_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_11_2_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_11_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25913),
            .lcout(\POWERLED.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_3_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_3_0  (
            .in0(_gnd_net_),
            .in1(N__26008),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(\POWERLED.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_11_3_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_11_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(N__25987),
            .in2(N__25851),
            .in3(N__25966),
            .lcout(\POWERLED.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_11_3_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_11_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__25847),
            .in2(N__25963),
            .in3(N__25942),
            .lcout(\POWERLED.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_11_3_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_11_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_11_3_3  (
            .in0(_gnd_net_),
            .in1(N__25939),
            .in2(N__25918),
            .in3(N__25921),
            .lcout(\POWERLED.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_11_3_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_11_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_11_3_4  (
            .in0(_gnd_net_),
            .in1(N__25917),
            .in2(N__25882),
            .in3(N__25864),
            .lcout(\POWERLED.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_11_3_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_11_3_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_11_3_5  (
            .in0(N__25795),
            .in1(N__25861),
            .in2(N__25852),
            .in3(N__25825),
            .lcout(\POWERLED.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_11_3_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_11_3_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_11_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25822),
            .in3(N__25810),
            .lcout(\POWERLED.mult1_un61_sum_s_8 ),
            .ltout(\POWERLED.mult1_un61_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_3_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_3_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25777),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_14_LC_11_4_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_14_LC_11_4_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_14_LC_11_4_7 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \POWERLED.dutycycle_14_LC_11_4_7  (
            .in0(N__26133),
            .in1(N__26176),
            .in2(N__28177),
            .in3(N__26155),
            .lcout(\POWERLED.dutycycleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32735),
            .ce(),
            .sr(N__26630));
    defparam \POWERLED.dutycycle_RNI_4_12_LC_11_5_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_11_5_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_12_LC_11_5_0  (
            .in0(N__29825),
            .in1(N__29140),
            .in2(N__29485),
            .in3(N__30144),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_8_a3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_9_LC_11_5_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_9_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_9_LC_11_5_1 .LUT_INIT=16'b1111111100110000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_9_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__26041),
            .in2(N__26119),
            .in3(N__26440),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_7_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_13_LC_11_5_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_13_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_13_LC_11_5_2 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \POWERLED.dutycycle_RNI_13_LC_11_5_2  (
            .in0(N__26115),
            .in1(N__26032),
            .in2(N__26059),
            .in3(N__26017),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_9_LC_11_5_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_9_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_9_LC_11_5_3 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \POWERLED.dutycycle_RNI_4_9_LC_11_5_3  (
            .in0(N__29828),
            .in1(N__31360),
            .in2(N__27916),
            .in3(N__29635),
            .lcout(\POWERLED.un1_N_5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_7_LC_11_5_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_7_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_7_LC_11_5_4 .LUT_INIT=16'b1100100011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_2_7_LC_11_5_4  (
            .in0(N__31359),
            .in1(N__29137),
            .in2(N__29667),
            .in3(N__27766),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_8_6_tz_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_7_LC_11_5_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_7_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_7_LC_11_5_5 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_8_7_LC_11_5_5  (
            .in0(N__29138),
            .in1(N__29824),
            .in2(N__26035),
            .in3(N__27914),
            .lcout(\POWERLED.un1_dutycycle_53_8_2_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_10_LC_11_5_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_10_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_10_LC_11_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_10_LC_11_5_6  (
            .in0(N__30004),
            .in1(N__29139),
            .in2(N__31376),
            .in3(N__26016),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_9_LC_11_5_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_9_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_9_LC_11_5_7 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_9_LC_11_5_7  (
            .in0(_gnd_net_),
            .in1(N__29823),
            .in2(N__27915),
            .in3(N__31358),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_8_LC_11_6_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_8_LC_11_6_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_8_LC_11_6_0 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \POWERLED.dutycycle_8_LC_11_6_0  (
            .in0(N__27934),
            .in1(N__26232),
            .in2(N__31104),
            .in3(N__26242),
            .lcout(\POWERLED.dutycycleZ1Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32747),
            .ce(),
            .sr(N__26649));
    defparam \POWERLED.dutycycle_RNI73694_8_LC_11_6_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI73694_8_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI73694_8_LC_11_6_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \POWERLED.dutycycle_RNI73694_8_LC_11_6_1  (
            .in0(N__26241),
            .in1(N__31065),
            .in2(N__26233),
            .in3(N__27933),
            .lcout(\POWERLED.dutycycleZ0Z_1 ),
            .ltout(\POWERLED.dutycycleZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_11_LC_11_6_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_11_6_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \POWERLED.dutycycle_RNI_1_11_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__29872),
            .in2(N__26215),
            .in3(N__30113),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_1Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_12_LC_11_6_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_11_6_3 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_12_LC_11_6_3  (
            .in0(N__30114),
            .in1(N__29465),
            .in2(N__26212),
            .in3(N__29998),
            .lcout(\POWERLED.un1_dutycycle_53_57_a0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_10_LC_11_6_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_10_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_10_LC_11_6_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.dutycycle_RNI_10_10_LC_11_6_4  (
            .in0(N__31369),
            .in1(N__29616),
            .in2(N__30013),
            .in3(N__29273),
            .lcout(\POWERLED.dutycycle_RNI_10Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_LC_11_6_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_LC_11_6_5 .LUT_INIT=16'b1111111010100000;
    LogicCell40 \POWERLED.dutycycle_RNI_10_LC_11_6_5  (
            .in0(N__30115),
            .in1(N__29659),
            .in2(N__29886),
            .in3(N__29997),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_10_LC_11_6_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_10_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_10_LC_11_6_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \POWERLED.dutycycle_RNI_11_10_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(N__27925),
            .in2(N__26197),
            .in3(N__26194),
            .lcout(\POWERLED.dutycycle_RNI_11Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOBHB2_11_LC_11_7_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOBHB2_11_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOBHB2_11_LC_11_7_0 .LUT_INIT=16'b1100110011101111;
    LogicCell40 \POWERLED.dutycycle_RNIOBHB2_11_LC_11_7_0  (
            .in0(N__30117),
            .in1(N__28599),
            .in2(N__31103),
            .in3(N__28461),
            .lcout(\POWERLED.dutycycle_eena_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_10_LC_11_7_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_10_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_10_LC_11_7_1 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \POWERLED.dutycycle_RNI_4_10_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29993),
            .in3(N__30116),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_13_a1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_LC_11_7_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_LC_11_7_2 .LUT_INIT=16'b0010000011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_8_LC_11_7_2  (
            .in0(N__26764),
            .in1(N__29605),
            .in2(N__26314),
            .in3(N__26251),
            .lcout(\POWERLED.un1_dutycycle_53_axb_11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_11_LC_11_7_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_11_LC_11_7_3 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_11_LC_11_7_3 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.dutycycle_11_LC_11_7_3  (
            .in0(N__26311),
            .in1(N__26278),
            .in2(N__28148),
            .in3(N__26298),
            .lcout(\POWERLED.dutycycleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32751),
            .ce(),
            .sr(N__26650));
    defparam \POWERLED.dutycycle_RNI_6_7_LC_11_7_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_7_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_7_LC_11_7_4 .LUT_INIT=16'b0101011111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_6_7_LC_11_7_4  (
            .in0(N__31346),
            .in1(N__29864),
            .in2(N__29155),
            .in3(N__26266),
            .lcout(\POWERLED.dutycycle_RNI_6Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5VRL4_11_LC_11_7_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5VRL4_11_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5VRL4_11_LC_11_7_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.dutycycle_RNI5VRL4_11_LC_11_7_5  (
            .in0(N__28111),
            .in1(N__26310),
            .in2(N__26299),
            .in3(N__26277),
            .lcout(\POWERLED.dutycycleZ0Z_7 ),
            .ltout(\POWERLED.dutycycleZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_10_LC_11_7_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_10_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_10_LC_11_7_6 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_10_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__29604),
            .in2(N__26269),
            .in3(N__29954),
            .lcout(\POWERLED.un1_dutycycle_53_46_a3_1 ),
            .ltout(\POWERLED.un1_dutycycle_53_46_a3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_6_LC_11_7_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_6_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_6_LC_11_7_7 .LUT_INIT=16'b0111111100101010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_6_LC_11_7_7  (
            .in0(N__27905),
            .in1(N__31347),
            .in2(N__26260),
            .in3(N__26257),
            .lcout(\POWERLED.un1_dutycycle_53_46_a3_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOBHB2_12_LC_11_8_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOBHB2_12_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOBHB2_12_LC_11_8_0 .LUT_INIT=16'b1010111010101111;
    LogicCell40 \POWERLED.dutycycle_RNIOBHB2_12_LC_11_8_0  (
            .in0(N__28598),
            .in1(N__29438),
            .in2(N__28483),
            .in3(N__31114),
            .lcout(\POWERLED.dutycycle_eena_9 ),
            .ltout(\POWERLED.dutycycle_eena_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_12_LC_11_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_12_LC_11_8_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_12_LC_11_8_1 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \POWERLED.dutycycle_12_LC_11_8_1  (
            .in0(N__26485),
            .in1(N__26467),
            .in2(N__26245),
            .in3(N__28155),
            .lcout(\POWERLED.dutycycleZ1Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32857),
            .ce(),
            .sr(N__26634));
    defparam \POWERLED.dutycycle_10_LC_11_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_10_LC_11_8_2 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_10_LC_11_8_2 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \POWERLED.dutycycle_10_LC_11_8_2  (
            .in0(N__26518),
            .in1(N__26500),
            .in2(N__28170),
            .in3(N__26512),
            .lcout(\POWERLED.dutycycleZ1Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32857),
            .ce(),
            .sr(N__26634));
    defparam \POWERLED.dutycycle_RNIOBHB2_10_LC_11_8_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOBHB2_10_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOBHB2_10_LC_11_8_3 .LUT_INIT=16'b1010101011101111;
    LogicCell40 \POWERLED.dutycycle_RNIOBHB2_10_LC_11_8_3  (
            .in0(N__28597),
            .in1(N__30003),
            .in2(N__31117),
            .in3(N__28469),
            .lcout(\POWERLED.dutycycle_eena_4 ),
            .ltout(\POWERLED.dutycycle_eena_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNISAA84_10_LC_11_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNISAA84_10_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNISAA84_10_LC_11_8_4 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.dutycycle_RNISAA84_10_LC_11_8_4  (
            .in0(N__28150),
            .in1(N__26511),
            .in2(N__26503),
            .in3(N__26499),
            .lcout(\POWERLED.dutycycleZ0Z_5 ),
            .ltout(\POWERLED.dutycycleZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_12_LC_11_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_11_8_5 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_12_LC_11_8_5  (
            .in0(N__29437),
            .in1(N__29871),
            .in2(N__26488),
            .in3(N__29639),
            .lcout(\POWERLED.un1_dutycycle_53_7_3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI72TL4_12_LC_11_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI72TL4_12_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI72TL4_12_LC_11_8_6 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.dutycycle_RNI72TL4_12_LC_11_8_6  (
            .in0(N__28151),
            .in1(N__26484),
            .in2(N__26476),
            .in3(N__26466),
            .lcout(\POWERLED.dutycycleZ0Z_10 ),
            .ltout(\POWERLED.dutycycleZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_12_LC_11_8_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_11_8_7 .LUT_INIT=16'b1100110111101100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_12_LC_11_8_7  (
            .in0(N__26449),
            .in1(N__27757),
            .in2(N__26443),
            .in3(N__30118),
            .lcout(\POWERLED.un1_dutycycle_53_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_2_LC_11_9_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_2_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_2_LC_11_9_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_2_LC_11_9_0  (
            .in0(N__26427),
            .in1(N__30551),
            .in2(N__30274),
            .in3(N__26940),
            .lcout(\POWERLED.N_414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_6_LC_11_9_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_6_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_6_LC_11_9_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_6_LC_11_9_1  (
            .in0(N__29327),
            .in1(N__26344),
            .in2(_gnd_net_),
            .in3(N__31341),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_6_LC_11_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_6_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_6_LC_11_9_2 .LUT_INIT=16'b0000000010111111;
    LogicCell40 \POWERLED.dutycycle_RNI_4_6_LC_11_9_2  (
            .in0(N__31342),
            .in1(N__26809),
            .in2(N__29334),
            .in3(N__28668),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_172_m2s4_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_6_LC_11_9_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_6_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_6_LC_11_9_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_6_LC_11_9_3  (
            .in0(N__30770),
            .in1(N__30678),
            .in2(N__26317),
            .in3(N__26779),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_172_m2s4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_6_LC_11_9_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_6_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_6_LC_11_9_4 .LUT_INIT=16'b1111000111110001;
    LogicCell40 \POWERLED.dutycycle_RNI_7_6_LC_11_9_4  (
            .in0(N__30679),
            .in1(N__26818),
            .in2(N__26812),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_7Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_3_LC_11_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_3_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_3_LC_11_9_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \POWERLED.dutycycle_RNI_7_3_LC_11_9_5  (
            .in0(N__26808),
            .in1(N__29298),
            .in2(N__28669),
            .in3(N__28950),
            .lcout(\POWERLED.dutycycle_RNI_7Z0Z_3 ),
            .ltout(\POWERLED.dutycycle_RNI_7Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQ8072_2_LC_11_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQ8072_2_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQ8072_2_LC_11_9_6 .LUT_INIT=16'b1100000011001010;
    LogicCell40 \POWERLED.dutycycle_RNIQ8072_2_LC_11_9_6  (
            .in0(N__31897),
            .in1(N__26773),
            .in2(N__26767),
            .in3(N__31072),
            .lcout(POWERLED_g1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_4_LC_11_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_4_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_4_LC_11_9_7 .LUT_INIT=16'b0101011101011111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_4_LC_11_9_7  (
            .in0(N__29136),
            .in1(N__29870),
            .in2(N__31364),
            .in3(N__29297),
            .lcout(\POWERLED.g0_i_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIDNFD1_1_LC_11_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIDNFD1_1_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIDNFD1_1_LC_11_10_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.func_state_RNIDNFD1_1_LC_11_10_2  (
            .in0(N__31749),
            .in1(N__26755),
            .in2(N__26730),
            .in3(N__28856),
            .lcout(\POWERLED.N_462 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_12_LC_11_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_12_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_12_LC_11_10_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_12_LC_11_10_3  (
            .in0(N__29509),
            .in1(N__28270),
            .in2(N__29388),
            .in3(N__29475),
            .lcout(\POWERLED.g1_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_5_LC_11_10_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_5_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_5_LC_11_10_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_1_5_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__28855),
            .in2(_gnd_net_),
            .in3(N__30861),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_52_and_i_0_m3_1_rn_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIV0AS_5_LC_11_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIV0AS_5_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIV0AS_5_LC_11_10_5 .LUT_INIT=16'b1101000101010101;
    LogicCell40 \POWERLED.dutycycle_RNIV0AS_5_LC_11_10_5  (
            .in0(N__26679),
            .in1(N__30218),
            .in2(N__26668),
            .in3(N__26939),
            .lcout(POWERLED_un1_clk_100khz_52_and_i_0_m3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_5_LC_11_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_5_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_5_LC_11_10_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_4_5_LC_11_10_6  (
            .in0(N__28269),
            .in1(N__29381),
            .in2(N__30600),
            .in3(N__29508),
            .lcout(\POWERLED.m69_0_o2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_5_LC_11_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_5_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_5_LC_11_10_7 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_5_LC_11_10_7  (
            .in0(N__30568),
            .in1(N__30596),
            .in2(N__26941),
            .in3(N__30217),
            .lcout(N_110_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_RNIDV4H_15_LC_11_11_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_RNIDV4H_15_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_esr_RNIDV4H_15_LC_11_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.count_esr_RNIDV4H_15_LC_11_11_0  (
            .in0(N__27277),
            .in1(N__27610),
            .in2(N__27169),
            .in3(N__27628),
            .lcout(),
            .ltout(\RSMRST_PWRGD.un4_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIR8OP4_10_LC_11_11_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIR8OP4_10_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIR8OP4_10_LC_11_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIR8OP4_10_LC_11_11_1  (
            .in0(N__26860),
            .in1(N__26866),
            .in2(N__26887),
            .in3(N__26872),
            .lcout(\RSMRST_PWRGD.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI9RLK1_3_LC_11_11_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI9RLK1_3_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI9RLK1_3_LC_11_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.count_RNI9RLK1_3_LC_11_11_2  (
            .in0(N__27021),
            .in1(N__27036),
            .in2(N__27073),
            .in3(N__27006),
            .lcout(\RSMRST_PWRGD.un4_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIQUU91_10_LC_11_11_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIQUU91_10_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIQUU91_10_LC_11_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIQUU91_10_LC_11_11_3  (
            .in0(N__27051),
            .in1(N__27646),
            .in2(N__26974),
            .in3(N__26992),
            .lcout(\RSMRST_PWRGD.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIBFU91_13_LC_11_11_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIBFU91_13_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIBFU91_13_LC_11_11_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \RSMRST_PWRGD.count_RNIBFU91_13_LC_11_11_4  (
            .in0(N__27592),
            .in1(N__27102),
            .in2(N__26836),
            .in3(N__27087),
            .lcout(\RSMRST_PWRGD.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_11_11_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_11_11_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RSMRST_PWRGD.count_esr_RNO_0_15_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__27525),
            .in2(_gnd_net_),
            .in3(N__27127),
            .lcout(\RSMRST_PWRGD.N_42_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_0_LC_11_12_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_0_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_0_LC_11_12_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_0_LC_11_12_0  (
            .in0(N__27559),
            .in1(N__26832),
            .in2(N__26854),
            .in3(N__26853),
            .lcout(\RSMRST_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .clk(N__32957),
            .ce(),
            .sr(N__27137));
    defparam \RSMRST_PWRGD.count_1_LC_11_12_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_1_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_1_LC_11_12_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_1_LC_11_12_1  (
            .in0(N__27548),
            .in1(N__27103),
            .in2(_gnd_net_),
            .in3(N__27091),
            .lcout(\RSMRST_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .clk(N__32957),
            .ce(),
            .sr(N__27137));
    defparam \RSMRST_PWRGD.count_2_LC_11_12_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_2_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_2_LC_11_12_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_2_LC_11_12_2  (
            .in0(N__27560),
            .in1(N__27088),
            .in2(_gnd_net_),
            .in3(N__27076),
            .lcout(\RSMRST_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .clk(N__32957),
            .ce(),
            .sr(N__27137));
    defparam \RSMRST_PWRGD.count_3_LC_11_12_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_3_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_3_LC_11_12_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_3_LC_11_12_3  (
            .in0(N__27549),
            .in1(N__27069),
            .in2(_gnd_net_),
            .in3(N__27055),
            .lcout(\RSMRST_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .clk(N__32957),
            .ce(),
            .sr(N__27137));
    defparam \RSMRST_PWRGD.count_4_LC_11_12_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_4_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_4_LC_11_12_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_4_LC_11_12_4  (
            .in0(N__27561),
            .in1(N__27052),
            .in2(_gnd_net_),
            .in3(N__27040),
            .lcout(\RSMRST_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .clk(N__32957),
            .ce(),
            .sr(N__27137));
    defparam \RSMRST_PWRGD.count_5_LC_11_12_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_5_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_5_LC_11_12_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_5_LC_11_12_5  (
            .in0(N__27550),
            .in1(N__27037),
            .in2(_gnd_net_),
            .in3(N__27025),
            .lcout(\RSMRST_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .clk(N__32957),
            .ce(),
            .sr(N__27137));
    defparam \RSMRST_PWRGD.count_6_LC_11_12_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_6_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_6_LC_11_12_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_6_LC_11_12_6  (
            .in0(N__27562),
            .in1(N__27022),
            .in2(_gnd_net_),
            .in3(N__27010),
            .lcout(\RSMRST_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .clk(N__32957),
            .ce(),
            .sr(N__27137));
    defparam \RSMRST_PWRGD.count_7_LC_11_12_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_7_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_7_LC_11_12_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_7_LC_11_12_7  (
            .in0(N__27551),
            .in1(N__27007),
            .in2(_gnd_net_),
            .in3(N__26995),
            .lcout(\RSMRST_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .clk(N__32957),
            .ce(),
            .sr(N__27137));
    defparam \RSMRST_PWRGD.count_8_LC_11_13_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_8_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_8_LC_11_13_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_8_LC_11_13_0  (
            .in0(N__27555),
            .in1(N__26991),
            .in2(_gnd_net_),
            .in3(N__26977),
            .lcout(\RSMRST_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .clk(N__32961),
            .ce(),
            .sr(N__27139));
    defparam \RSMRST_PWRGD.count_9_LC_11_13_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_9_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_9_LC_11_13_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_9_LC_11_13_1  (
            .in0(N__27547),
            .in1(N__26970),
            .in2(_gnd_net_),
            .in3(N__26956),
            .lcout(\RSMRST_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .clk(N__32961),
            .ce(),
            .sr(N__27139));
    defparam \RSMRST_PWRGD.count_10_LC_11_13_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_10_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_10_LC_11_13_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_10_LC_11_13_2  (
            .in0(N__27552),
            .in1(N__27645),
            .in2(_gnd_net_),
            .in3(N__27631),
            .lcout(\RSMRST_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .clk(N__32961),
            .ce(),
            .sr(N__27139));
    defparam \RSMRST_PWRGD.count_11_LC_11_13_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_11_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_11_LC_11_13_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_11_LC_11_13_3  (
            .in0(N__27545),
            .in1(N__27627),
            .in2(_gnd_net_),
            .in3(N__27613),
            .lcout(\RSMRST_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .clk(N__32961),
            .ce(),
            .sr(N__27139));
    defparam \RSMRST_PWRGD.count_12_LC_11_13_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_12_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_12_LC_11_13_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_12_LC_11_13_4  (
            .in0(N__27553),
            .in1(N__27609),
            .in2(_gnd_net_),
            .in3(N__27595),
            .lcout(\RSMRST_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .clk(N__32961),
            .ce(),
            .sr(N__27139));
    defparam \RSMRST_PWRGD.count_13_LC_11_13_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_13_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_13_LC_11_13_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_13_LC_11_13_5  (
            .in0(N__27546),
            .in1(N__27591),
            .in2(_gnd_net_),
            .in3(N__27577),
            .lcout(\RSMRST_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .clk(N__32961),
            .ce(),
            .sr(N__27139));
    defparam \RSMRST_PWRGD.count_14_LC_11_13_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_14_LC_11_13_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_14_LC_11_13_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_14_LC_11_13_6  (
            .in0(N__27554),
            .in1(N__27276),
            .in2(_gnd_net_),
            .in3(N__27262),
            .lcout(\RSMRST_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .clk(N__32961),
            .ce(),
            .sr(N__27139));
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_13_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__27259),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_15_LC_11_14_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_15_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_esr_15_LC_11_14_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \RSMRST_PWRGD.count_esr_15_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__27165),
            .in2(_gnd_net_),
            .in3(N__27172),
            .lcout(\RSMRST_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33017),
            .ce(N__27151),
            .sr(N__27138));
    defparam \VPP_VDDQ.curr_state_2_0_LC_11_15_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_0_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_0_LC_11_15_3 .LUT_INIT=16'b0100010010100000;
    LogicCell40 \VPP_VDDQ.curr_state_2_0_LC_11_15_3  (
            .in0(N__33203),
            .in1(N__33114),
            .in2(N__33725),
            .in3(N__33391),
            .lcout(\VPP_VDDQ.curr_state_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32962),
            .ce(N__32291),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_i_LC_11_15_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_i_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_i_LC_11_15_4 .LUT_INIT=16'b1111001101011111;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m4_i_LC_11_15_4  (
            .in0(N__33115),
            .in1(N__33700),
            .in2(N__33452),
            .in3(N__33201),
            .lcout(),
            .ltout(\VPP_VDDQ.N_190_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_11_15_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_11_15_5 .LUT_INIT=16'b0000111111001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__27724),
            .in2(N__27718),
            .in3(N__33929),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_11_15_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_11_15_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_11_15_6  (
            .in0(N__27715),
            .in1(N__33701),
            .in2(N__27697),
            .in3(N__33202),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIF7361_3_LC_11_15_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIF7361_3_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIF7361_3_LC_11_15_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIF7361_3_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__27694),
            .in2(N__27682),
            .in3(N__32020),
            .lcout(\VPP_VDDQ.count_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_3_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_3_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27824),
            .lcout(\VPP_VDDQ.N_28_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_1_LC_12_3_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_1_LC_12_3_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_1_LC_12_3_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI8PF7_1_LC_12_3_3  (
            .in0(_gnd_net_),
            .in1(N__33135),
            .in2(_gnd_net_),
            .in3(N__31659),
            .lcout(\VPP_VDDQ.N_537_0 ),
            .ltout(\VPP_VDDQ.N_537_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_12_3_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_12_3_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_12_3_4 .LUT_INIT=16'b1111110011111111;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(N__33519),
            .in2(N__27661),
            .in3(N__33931),
            .lcout(\VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIVBNA1_0_LC_12_3_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIVBNA1_0_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIVBNA1_0_LC_12_3_5 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIVBNA1_0_LC_12_3_5  (
            .in0(N__33520),
            .in1(N__33136),
            .in2(N__27658),
            .in3(N__32318),
            .lcout(\VPP_VDDQ.delayed_vddq_ok_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_12_4_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_12_4_0 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_12_4_0  (
            .in0(N__31660),
            .in1(N__32315),
            .in2(N__27655),
            .in3(N__33497),
            .lcout(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_12_4_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_12_4_4 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_12_4_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_LC_12_4_4  (
            .in0(N__33133),
            .in1(N__27825),
            .in2(N__27810),
            .in3(N__27795),
            .lcout(\VPP_VDDQ.delayed_vddq_okZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32726),
            .ce(),
            .sr(N__27838));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNIEC852_LC_12_4_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNIEC852_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNIEC852_LC_12_4_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNIEC852_LC_12_4_6  (
            .in0(N__33134),
            .in1(N__27826),
            .in2(N__27811),
            .in3(N__27796),
            .lcout(VPP_VDDQ_delayed_vddq_ok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_9_LC_12_5_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_9_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_9_LC_12_5_0 .LUT_INIT=16'b1011001000110010;
    LogicCell40 \POWERLED.dutycycle_RNI_2_9_LC_12_5_0  (
            .in0(N__29615),
            .in1(N__27748),
            .in2(N__31374),
            .in3(N__29826),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_2Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_9_LC_12_5_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_9_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_9_LC_12_5_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_9_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(N__27739),
            .in2(N__27778),
            .in3(N__27912),
            .lcout(\POWERLED.dutycycle_RNI_6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_12_LC_12_5_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_12_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_12_LC_12_5_2 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \POWERLED.dutycycle_RNI_7_12_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(N__29476),
            .in2(N__29868),
            .in3(N__30143),
            .lcout(\POWERLED.un1_dutycycle_53_4_a0_1 ),
            .ltout(\POWERLED.un1_dutycycle_53_4_a0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_7_LC_12_5_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_7_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_7_LC_12_5_3 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_7_LC_12_5_3  (
            .in0(N__29157),
            .in1(N__31350),
            .in2(N__27760),
            .in3(N__29613),
            .lcout(\POWERLED.un1_dutycycle_53_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_7_LC_12_5_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_7_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_7_LC_12_5_4 .LUT_INIT=16'b0000010101011111;
    LogicCell40 \POWERLED.dutycycle_RNI_7_7_LC_12_5_4  (
            .in0(N__29614),
            .in1(_gnd_net_),
            .in2(N__29869),
            .in3(N__29158),
            .lcout(\POWERLED.un1_dutycycle_53_8_1 ),
            .ltout(\POWERLED.un1_dutycycle_53_8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_9_LC_12_5_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_9_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_9_LC_12_5_5 .LUT_INIT=16'b1000111110001110;
    LogicCell40 \POWERLED.dutycycle_RNI_1_9_LC_12_5_5  (
            .in0(N__29631),
            .in1(N__31351),
            .in2(N__27742),
            .in3(N__29822),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_LC_12_5_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_LC_12_5_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNI_5_LC_12_5_6  (
            .in0(N__27913),
            .in1(N__30880),
            .in2(N__31375),
            .in3(N__29827),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOBHB2_1_1_LC_12_5_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOBHB2_1_1_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOBHB2_1_1_LC_12_5_7 .LUT_INIT=16'b1100110011011111;
    LogicCell40 \POWERLED.func_state_RNIOBHB2_1_1_LC_12_5_7  (
            .in0(N__29389),
            .in1(N__28588),
            .in2(N__31116),
            .in3(N__28484),
            .lcout(\POWERLED.dutycycle_eena_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOGRS_8_LC_12_6_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOGRS_8_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOGRS_8_LC_12_6_0 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \POWERLED.dutycycle_RNIOGRS_8_LC_12_6_0  (
            .in0(N__29612),
            .in1(N__31108),
            .in2(_gnd_net_),
            .in3(N__28481),
            .lcout(),
            .ltout(\POWERLED.N_84_f0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIFOI43_8_LC_12_6_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIFOI43_8_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIFOI43_8_LC_12_6_1 .LUT_INIT=16'b1000111100000000;
    LogicCell40 \POWERLED.dutycycle_RNIFOI43_8_LC_12_6_1  (
            .in0(N__31720),
            .in1(N__28216),
            .in2(N__28180),
            .in3(N__28149),
            .lcout(\POWERLED.dutycycle_en_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_11_LC_12_6_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_12_6_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.dutycycle_RNI_2_11_LC_12_6_2  (
            .in0(N__29879),
            .in1(N__29131),
            .in2(N__31377),
            .in3(N__30109),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_10_LC_12_6_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_10_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_10_LC_12_6_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_10_LC_12_6_3  (
            .in0(N__29132),
            .in1(N__29999),
            .in2(N__30146),
            .in3(N__29611),
            .lcout(),
            .ltout(\POWERLED.N_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_4_LC_12_6_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_4_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_4_LC_12_6_4 .LUT_INIT=16'b1111100011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_9_4_LC_12_6_4  (
            .in0(N__27844),
            .in1(N__28372),
            .in2(N__27919),
            .in3(N__28240),
            .lcout(\POWERLED.g0_i_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_3_LC_12_6_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_12_6_5 .LUT_INIT=16'b1111100011100000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_3_LC_12_6_5  (
            .in0(N__29130),
            .in1(N__28962),
            .in2(N__29295),
            .in3(N__29609),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_3_LC_12_6_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_12_6_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_3_LC_12_6_6  (
            .in0(N__28963),
            .in1(_gnd_net_),
            .in2(N__28366),
            .in3(N__27880),
            .lcout(\POWERLED.un1_dutycycle_53_25_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_4_LC_12_6_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_4_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_4_LC_12_6_7 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_4_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(N__31365),
            .in2(N__29296),
            .in3(N__29610),
            .lcout(\POWERLED.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_15_LC_12_7_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_15_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_15_LC_12_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_1_15_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28653),
            .lcout(\POWERLED.N_2191_i ),
            .ltout(\POWERLED.N_2191_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOBHB2_1_LC_12_7_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOBHB2_1_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOBHB2_1_LC_12_7_1 .LUT_INIT=16'b1100110011011111;
    LogicCell40 \POWERLED.func_state_RNIOBHB2_1_LC_12_7_1  (
            .in0(N__31098),
            .in1(N__28600),
            .in2(N__28489),
            .in3(N__28482),
            .lcout(\POWERLED.dutycycle_eena_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_10_LC_12_7_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_10_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_10_LC_12_7_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_10_LC_12_7_2  (
            .in0(N__29965),
            .in1(N__29145),
            .in2(N__29884),
            .in3(N__30104),
            .lcout(\POWERLED.g0_i_i_a6_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_4_LC_12_7_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_4_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_4_LC_12_7_3 .LUT_INIT=16'b0001011100011111;
    LogicCell40 \POWERLED.dutycycle_RNI_4_4_LC_12_7_3  (
            .in0(N__29607),
            .in1(N__31348),
            .in2(N__29156),
            .in3(N__29294),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_LC_12_7_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_LC_12_7_4 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \POWERLED.dutycycle_RNI_4_LC_12_7_4  (
            .in0(N__29293),
            .in1(N__29141),
            .in2(N__29883),
            .in3(N__29606),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_14_LC_12_7_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_14_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_14_LC_12_7_5 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \POWERLED.dutycycle_RNI_2_14_LC_12_7_5  (
            .in0(N__28356),
            .in1(N__30166),
            .in2(N__28303),
            .in3(N__28294),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_10_LC_12_7_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_10_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_10_LC_12_7_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \POWERLED.dutycycle_RNI_5_10_LC_12_7_6  (
            .in0(N__29967),
            .in1(N__28268),
            .in2(_gnd_net_),
            .in3(N__30108),
            .lcout(\POWERLED.un2_count_clk_17_0_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_10_LC_12_7_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_10_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_10_LC_12_7_7 .LUT_INIT=16'b1110001101111100;
    LogicCell40 \POWERLED.dutycycle_RNI_1_10_LC_12_7_7  (
            .in0(N__29608),
            .in1(N__29863),
            .in2(N__30145),
            .in3(N__29966),
            .lcout(\POWERLED.un1_dutycycle_53_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_4_LC_12_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_4_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_4_LC_12_8_1 .LUT_INIT=16'b0001001100011111;
    LogicCell40 \POWERLED.dutycycle_RNI_6_4_LC_12_8_1  (
            .in0(N__29307),
            .in1(N__29151),
            .in2(N__31378),
            .in3(N__29671),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_6Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_3_LC_12_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_12_8_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_3_LC_12_8_2  (
            .in0(N__28953),
            .in1(_gnd_net_),
            .in2(N__30178),
            .in3(N__30175),
            .lcout(),
            .ltout(\POWERLED.o2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_10_LC_12_8_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_10_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_10_LC_12_8_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_10_LC_12_8_3  (
            .in0(N__29880),
            .in1(N__29971),
            .in2(N__30169),
            .in3(N__30119),
            .lcout(\POWERLED.dutycycle_RNI_7Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_10_LC_12_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_10_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_10_LC_12_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.dutycycle_RNI_9_10_LC_12_8_4  (
            .in0(N__29673),
            .in1(N__29882),
            .in2(N__30147),
            .in3(N__29978),
            .lcout(\POWERLED.g1_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_9_LC_12_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_9_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_9_LC_12_8_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_9_LC_12_8_5  (
            .in0(N__29881),
            .in1(N__29672),
            .in2(N__29502),
            .in3(N__31405),
            .lcout(),
            .ltout(\POWERLED.un2_count_clk_17_0_0_a2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_12_LC_12_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_12_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_12_LC_12_8_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_12_LC_12_8_6  (
            .in0(N__29453),
            .in1(N__29377),
            .in2(N__29347),
            .in3(N__29344),
            .lcout(\POWERLED.N_501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_3_LC_12_8_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_12_8_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.dutycycle_RNI_6_3_LC_12_8_7  (
            .in0(N__29308),
            .in1(N__29152),
            .in2(_gnd_net_),
            .in3(N__28952),
            .lcout(\POWERLED.N_493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_LC_12_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_LC_12_9_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \POWERLED.func_state_RNI_1_LC_12_9_3  (
            .in0(N__30676),
            .in1(N__31896),
            .in2(_gnd_net_),
            .in3(N__28819),
            .lcout(\POWERLED.un2_count_clk_17_0_1 ),
            .ltout(\POWERLED.un2_count_clk_17_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_6_LC_12_9_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_6_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_6_LC_12_9_4 .LUT_INIT=16'b0111011101110000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_6_LC_12_9_4  (
            .in0(N__30771),
            .in1(N__30677),
            .in2(N__28657),
            .in3(N__31189),
            .lcout(N_46),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_1_LC_12_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_1_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_1_LC_12_9_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_1_LC_12_9_6  (
            .in0(N__31549),
            .in1(N__31479),
            .in2(_gnd_net_),
            .in3(N__31404),
            .lcout(),
            .ltout(\POWERLED.g1_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_6_LC_12_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_6_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_6_LC_12_9_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_6_LC_12_9_7  (
            .in0(N__31393),
            .in1(N__31387),
            .in2(N__31381),
            .in3(N__31373),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIOGRS_LC_12_10_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIOGRS_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIOGRS_LC_12_10_0 .LUT_INIT=16'b1110110011100100;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_fast_RNIOGRS_LC_12_10_0  (
            .in0(N__30613),
            .in1(N__30577),
            .in2(N__30878),
            .in3(N__31182),
            .lcout(),
            .ltout(\RSMRST_PWRGD.N_8_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIG1NP1_LC_12_10_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIG1NP1_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIG1NP1_LC_12_10_1 .LUT_INIT=16'b0000111100101111;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_fast_RNIG1NP1_LC_12_10_1  (
            .in0(N__31883),
            .in1(N__30612),
            .in2(N__31120),
            .in3(N__31110),
            .lcout(),
            .ltout(\RSMRST_PWRGD.N_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIAAN04_LC_12_10_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIAAN04_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_RNIAAN04_LC_12_10_2 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_fast_RNIAAN04_LC_12_10_2  (
            .in0(N__30865),
            .in1(N__30796),
            .in2(N__30790),
            .in3(N__30787),
            .lcout(\RSMRST_PWRGD.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_2_1_LC_12_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_2_1_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_2_1_LC_12_10_4 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \POWERLED.func_state_RNI_2_1_LC_12_10_4  (
            .in0(N__30772),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30700),
            .lcout(N_22_0),
            .ltout(N_22_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_S4n_RNI5DLR_LC_12_10_5.C_ON=1'b0;
    defparam SLP_S4n_RNI5DLR_LC_12_10_5.SEQ_MODE=4'b0000;
    defparam SLP_S4n_RNI5DLR_LC_12_10_5.LUT_INIT=16'b0010000000101111;
    LogicCell40 SLP_S4n_RNI5DLR_LC_12_10_5 (
            .in0(N__30570),
            .in1(N__30276),
            .in2(N__30604),
            .in3(N__30601),
            .lcout(g0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8H551_0_LC_12_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8H551_0_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8H551_0_LC_12_10_7 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \POWERLED.func_state_RNI8H551_0_LC_12_10_7  (
            .in0(N__30569),
            .in1(N__30275),
            .in2(N__31895),
            .in3(N__31748),
            .lcout(\POWERLED.dutycycle_1_0_iv_i_a2_sx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_12_12_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_12_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_1_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33232),
            .lcout(\VPP_VDDQ.N_2112_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_12_13_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_12_13_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_12_13_0  (
            .in0(N__33234),
            .in1(N__31560),
            .in2(N__33459),
            .in3(N__33715),
            .lcout(\VPP_VDDQ.count_2_1_7 ),
            .ltout(\VPP_VDDQ.count_2_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINJ761_0_7_LC_12_13_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINJ761_0_7_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINJ761_0_7_LC_12_13_1 .LUT_INIT=16'b0000010100010001;
    LogicCell40 \VPP_VDDQ.count_2_RNINJ761_0_7_LC_12_13_1  (
            .in0(N__31642),
            .in1(N__32224),
            .in2(N__31621),
            .in3(N__32078),
            .lcout(),
            .ltout(\VPP_VDDQ.un9_clk_100khz_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINJ761_1_7_LC_12_13_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINJ761_1_7_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINJ761_1_7_LC_12_13_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.count_2_RNINJ761_1_7_LC_12_13_2  (
            .in0(N__31618),
            .in1(N__31606),
            .in2(N__31588),
            .in3(N__31908),
            .lcout(\VPP_VDDQ.un9_clk_100khz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_0_LC_12_13_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_0_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_0_LC_12_13_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \VPP_VDDQ.count_2_RNI_0_LC_12_13_3  (
            .in0(N__33714),
            .in1(N__33401),
            .in2(N__32169),
            .in3(N__33233),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIT1QU_0_LC_12_13_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIT1QU_0_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIT1QU_0_LC_12_13_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIT1QU_0_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__31567),
            .in2(N__31573),
            .in3(N__31987),
            .lcout(\VPP_VDDQ.count_2Z0Z_0 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_0_LC_12_13_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_0_LC_12_13_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_0_LC_12_13_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \VPP_VDDQ.count_2_0_LC_12_13_5  (
            .in0(N__33716),
            .in1(N__33405),
            .in2(N__31570),
            .in3(N__33236),
            .lcout(\VPP_VDDQ.count_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33038),
            .ce(N__32077),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_7_LC_12_13_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_7_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_7_LC_12_13_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.count_2_7_LC_12_13_6  (
            .in0(N__33235),
            .in1(N__31561),
            .in2(N__33460),
            .in3(N__33717),
            .lcout(\VPP_VDDQ.count_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33038),
            .ce(N__32077),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINJ761_7_LC_12_13_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINJ761_7_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINJ761_7_LC_12_13_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_2_RNINJ761_7_LC_12_13_7  (
            .in0(N__31988),
            .in1(N__32223),
            .in2(_gnd_net_),
            .in3(N__32215),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_1_LC_12_14_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_12_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \VPP_VDDQ.count_2_RNI_1_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__32158),
            .in2(_gnd_net_),
            .in3(N__32190),
            .lcout(\VPP_VDDQ.count_2_RNIZ0Z_1 ),
            .ltout(\VPP_VDDQ.count_2_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_14_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_14_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_14_1  (
            .in0(N__33184),
            .in1(N__33706),
            .in2(N__32200),
            .in3(N__33363),
            .lcout(\VPP_VDDQ.count_2_1_1 ),
            .ltout(\VPP_VDDQ.count_2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIU2QU_1_LC_12_14_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIU2QU_1_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIU2QU_1_LC_12_14_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNIU2QU_1_LC_12_14_2  (
            .in0(N__32118),
            .in1(_gnd_net_),
            .in2(N__32197),
            .in3(N__31986),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_12_14_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_12_14_3 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_12_14_3  (
            .in0(N__32176),
            .in1(N__32119),
            .in2(N__32168),
            .in3(N__32034),
            .lcout(\VPP_VDDQ.un9_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_1_LC_12_14_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_1_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_1_LC_12_14_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.count_2_1_LC_12_14_4  (
            .in0(N__33364),
            .in1(N__33188),
            .in2(N__33726),
            .in3(N__32125),
            .lcout(\VPP_VDDQ.count_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33015),
            .ce(N__32032),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_11_LC_12_14_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_11_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_11_LC_12_14_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.count_2_11_LC_12_14_5  (
            .in0(N__32109),
            .in1(N__33710),
            .in2(N__33231),
            .in3(N__33365),
            .lcout(\VPP_VDDQ.count_2_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33015),
            .ce(N__32032),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_14_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_14_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_14_6  (
            .in0(N__33366),
            .in1(N__32110),
            .in2(N__33727),
            .in3(N__33183),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIDR4C1_11_LC_12_14_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIDR4C1_11_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIDR4C1_11_LC_12_14_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIDR4C1_11_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__32098),
            .in2(N__32092),
            .in3(N__32033),
            .lcout(\VPP_VDDQ.count_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_12_15_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_12_15_1 .LUT_INIT=16'b1111101011110011;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_12_15_1  (
            .in0(N__33724),
            .in1(N__33088),
            .in2(N__33496),
            .in3(N__33230),
            .lcout(),
            .ltout(\VPP_VDDQ.N_178_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_12_15_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_12_15_2 .LUT_INIT=16'b0000111111001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__33070),
            .in2(N__34030),
            .in3(N__33928),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_1_LC_12_16_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_1_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_1_LC_12_16_5 .LUT_INIT=16'b0001001100010000;
    LogicCell40 \VPP_VDDQ.curr_state_2_1_LC_12_16_5  (
            .in0(N__33723),
            .in1(N__33395),
            .in2(N__33281),
            .in3(N__33116),
            .lcout(\VPP_VDDQ.curr_state_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33016),
            .ce(N__32292),
            .sr(_gnd_net_));
endmodule // TOP
