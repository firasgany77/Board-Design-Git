// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 13 2022 11:36:22

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VR_READY_VCCINAUX,
    V33A_ENn,
    V1P8A_EN,
    VDDQ_EN,
    VCCST_OVERRIDE_3V3,
    V5S_OK,
    SLP_S3n,
    SLP_S0n,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    GPIO_FPGA_SoC_2,
    VCCIN_VR_PROCHOT_FPGA,
    SLP_SUSn,
    CPU_C10_GATE_N,
    VCCST_EN,
    V33DSW_OK,
    TPM_GPIO,
    SUSWARN_N,
    PLTRSTn,
    GPIO_FPGA_SoC_4,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    FPGA_OSC,
    VCCST_PWRGD,
    SYS_PWROK,
    SPI_FP_IO2,
    SATAXPCIE1_FPGA,
    GPIO_FPGA_EXP_1,
    VCCINAUX_VR_PROCHOT_FPGA,
    VCCINAUX_VR_PE,
    HDA_SDO_ATP,
    GPIO_FPGA_EXP_2,
    VPP_EN,
    VDDQ_OK,
    SUSACK_N,
    SLP_S4n,
    VCCST_CPU_OK,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    GPIO_FPGA_SoC_1,
    DSW_PWROK,
    V5A_EN,
    GPIO_FPGA_SoC_3,
    VR_PROCHOT_FPGA_OUT_N,
    VPP_OK,
    VCCIN_VR_PE,
    VCCIN_EN,
    SOC_SPKR,
    SLP_S5n,
    V12_MAIN_MON,
    SPI_FP_IO3,
    SATAXPCIE0_FPGA,
    V33A_OK,
    PCH_PWROK,
    FPGA_SLP_WLAN_N);

    input VR_READY_VCCINAUX;
    output V33A_ENn;
    output V1P8A_EN;
    output VDDQ_EN;
    input VCCST_OVERRIDE_3V3;
    input V5S_OK;
    input SLP_S3n;
    input SLP_S0n;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input GPIO_FPGA_SoC_2;
    input VCCIN_VR_PROCHOT_FPGA;
    input SLP_SUSn;
    input CPU_C10_GATE_N;
    output VCCST_EN;
    input V33DSW_OK;
    input TPM_GPIO;
    input SUSWARN_N;
    input PLTRSTn;
    input GPIO_FPGA_SoC_4;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output SYS_PWROK;
    input SPI_FP_IO2;
    input SATAXPCIE1_FPGA;
    input GPIO_FPGA_EXP_1;
    input VCCINAUX_VR_PROCHOT_FPGA;
    output VCCINAUX_VR_PE;
    output HDA_SDO_ATP;
    input GPIO_FPGA_EXP_2;
    output VPP_EN;
    input VDDQ_OK;
    input SUSACK_N;
    input SLP_S4n;
    input VCCST_CPU_OK;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input GPIO_FPGA_SoC_1;
    output DSW_PWROK;
    output V5A_EN;
    input GPIO_FPGA_SoC_3;
    input VR_PROCHOT_FPGA_OUT_N;
    input VPP_OK;
    output VCCIN_VR_PE;
    output VCCIN_EN;
    input SOC_SPKR;
    input SLP_S5n;
    input V12_MAIN_MON;
    input SPI_FP_IO3;
    input SATAXPCIE0_FPGA;
    input V33A_OK;
    output PCH_PWROK;
    input FPGA_SLP_WLAN_N;

    wire N__33702;
    wire N__33701;
    wire N__33700;
    wire N__33693;
    wire N__33692;
    wire N__33691;
    wire N__33684;
    wire N__33683;
    wire N__33682;
    wire N__33675;
    wire N__33674;
    wire N__33673;
    wire N__33666;
    wire N__33665;
    wire N__33664;
    wire N__33657;
    wire N__33656;
    wire N__33655;
    wire N__33648;
    wire N__33647;
    wire N__33646;
    wire N__33639;
    wire N__33638;
    wire N__33637;
    wire N__33630;
    wire N__33629;
    wire N__33628;
    wire N__33621;
    wire N__33620;
    wire N__33619;
    wire N__33612;
    wire N__33611;
    wire N__33610;
    wire N__33603;
    wire N__33602;
    wire N__33601;
    wire N__33594;
    wire N__33593;
    wire N__33592;
    wire N__33585;
    wire N__33584;
    wire N__33583;
    wire N__33576;
    wire N__33575;
    wire N__33574;
    wire N__33567;
    wire N__33566;
    wire N__33565;
    wire N__33558;
    wire N__33557;
    wire N__33556;
    wire N__33549;
    wire N__33548;
    wire N__33547;
    wire N__33540;
    wire N__33539;
    wire N__33538;
    wire N__33531;
    wire N__33530;
    wire N__33529;
    wire N__33522;
    wire N__33521;
    wire N__33520;
    wire N__33513;
    wire N__33512;
    wire N__33511;
    wire N__33504;
    wire N__33503;
    wire N__33502;
    wire N__33495;
    wire N__33494;
    wire N__33493;
    wire N__33486;
    wire N__33485;
    wire N__33484;
    wire N__33477;
    wire N__33476;
    wire N__33475;
    wire N__33468;
    wire N__33467;
    wire N__33466;
    wire N__33459;
    wire N__33458;
    wire N__33457;
    wire N__33450;
    wire N__33449;
    wire N__33448;
    wire N__33441;
    wire N__33440;
    wire N__33439;
    wire N__33432;
    wire N__33431;
    wire N__33430;
    wire N__33423;
    wire N__33422;
    wire N__33421;
    wire N__33414;
    wire N__33413;
    wire N__33412;
    wire N__33405;
    wire N__33404;
    wire N__33403;
    wire N__33396;
    wire N__33395;
    wire N__33394;
    wire N__33387;
    wire N__33386;
    wire N__33385;
    wire N__33378;
    wire N__33377;
    wire N__33376;
    wire N__33369;
    wire N__33368;
    wire N__33367;
    wire N__33360;
    wire N__33359;
    wire N__33358;
    wire N__33351;
    wire N__33350;
    wire N__33349;
    wire N__33342;
    wire N__33341;
    wire N__33340;
    wire N__33333;
    wire N__33332;
    wire N__33331;
    wire N__33324;
    wire N__33323;
    wire N__33322;
    wire N__33315;
    wire N__33314;
    wire N__33313;
    wire N__33306;
    wire N__33305;
    wire N__33304;
    wire N__33297;
    wire N__33296;
    wire N__33295;
    wire N__33288;
    wire N__33287;
    wire N__33286;
    wire N__33279;
    wire N__33278;
    wire N__33277;
    wire N__33270;
    wire N__33269;
    wire N__33268;
    wire N__33261;
    wire N__33260;
    wire N__33259;
    wire N__33252;
    wire N__33251;
    wire N__33250;
    wire N__33243;
    wire N__33242;
    wire N__33241;
    wire N__33234;
    wire N__33233;
    wire N__33232;
    wire N__33225;
    wire N__33224;
    wire N__33223;
    wire N__33216;
    wire N__33215;
    wire N__33214;
    wire N__33207;
    wire N__33206;
    wire N__33205;
    wire N__33198;
    wire N__33197;
    wire N__33196;
    wire N__33189;
    wire N__33188;
    wire N__33187;
    wire N__33180;
    wire N__33179;
    wire N__33178;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33152;
    wire N__33149;
    wire N__33146;
    wire N__33145;
    wire N__33144;
    wire N__33141;
    wire N__33136;
    wire N__33131;
    wire N__33130;
    wire N__33129;
    wire N__33128;
    wire N__33127;
    wire N__33124;
    wire N__33123;
    wire N__33120;
    wire N__33117;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33101;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33087;
    wire N__33086;
    wire N__33085;
    wire N__33084;
    wire N__33081;
    wire N__33078;
    wire N__33077;
    wire N__33074;
    wire N__33069;
    wire N__33068;
    wire N__33067;
    wire N__33064;
    wire N__33063;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33049;
    wire N__33044;
    wire N__33039;
    wire N__33026;
    wire N__33023;
    wire N__33020;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32987;
    wire N__32984;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32956;
    wire N__32955;
    wire N__32954;
    wire N__32953;
    wire N__32950;
    wire N__32949;
    wire N__32948;
    wire N__32945;
    wire N__32944;
    wire N__32941;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32913;
    wire N__32910;
    wire N__32905;
    wire N__32902;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32890;
    wire N__32887;
    wire N__32880;
    wire N__32875;
    wire N__32864;
    wire N__32861;
    wire N__32858;
    wire N__32855;
    wire N__32852;
    wire N__32849;
    wire N__32846;
    wire N__32843;
    wire N__32842;
    wire N__32837;
    wire N__32836;
    wire N__32835;
    wire N__32834;
    wire N__32833;
    wire N__32832;
    wire N__32831;
    wire N__32828;
    wire N__32827;
    wire N__32826;
    wire N__32825;
    wire N__32822;
    wire N__32821;
    wire N__32816;
    wire N__32815;
    wire N__32814;
    wire N__32813;
    wire N__32812;
    wire N__32811;
    wire N__32806;
    wire N__32803;
    wire N__32800;
    wire N__32797;
    wire N__32794;
    wire N__32793;
    wire N__32792;
    wire N__32789;
    wire N__32784;
    wire N__32783;
    wire N__32780;
    wire N__32775;
    wire N__32772;
    wire N__32769;
    wire N__32768;
    wire N__32765;
    wire N__32754;
    wire N__32749;
    wire N__32746;
    wire N__32745;
    wire N__32744;
    wire N__32741;
    wire N__32740;
    wire N__32737;
    wire N__32732;
    wire N__32727;
    wire N__32724;
    wire N__32715;
    wire N__32712;
    wire N__32709;
    wire N__32706;
    wire N__32703;
    wire N__32698;
    wire N__32691;
    wire N__32678;
    wire N__32675;
    wire N__32674;
    wire N__32673;
    wire N__32672;
    wire N__32671;
    wire N__32670;
    wire N__32669;
    wire N__32668;
    wire N__32667;
    wire N__32664;
    wire N__32661;
    wire N__32656;
    wire N__32653;
    wire N__32650;
    wire N__32647;
    wire N__32646;
    wire N__32645;
    wire N__32644;
    wire N__32641;
    wire N__32640;
    wire N__32639;
    wire N__32638;
    wire N__32637;
    wire N__32634;
    wire N__32631;
    wire N__32630;
    wire N__32629;
    wire N__32628;
    wire N__32627;
    wire N__32626;
    wire N__32621;
    wire N__32614;
    wire N__32611;
    wire N__32608;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32594;
    wire N__32593;
    wire N__32590;
    wire N__32587;
    wire N__32584;
    wire N__32579;
    wire N__32576;
    wire N__32575;
    wire N__32570;
    wire N__32567;
    wire N__32562;
    wire N__32559;
    wire N__32556;
    wire N__32553;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32534;
    wire N__32529;
    wire N__32522;
    wire N__32515;
    wire N__32510;
    wire N__32507;
    wire N__32492;
    wire N__32489;
    wire N__32488;
    wire N__32483;
    wire N__32480;
    wire N__32479;
    wire N__32476;
    wire N__32473;
    wire N__32472;
    wire N__32471;
    wire N__32470;
    wire N__32469;
    wire N__32468;
    wire N__32467;
    wire N__32466;
    wire N__32465;
    wire N__32464;
    wire N__32463;
    wire N__32462;
    wire N__32461;
    wire N__32460;
    wire N__32459;
    wire N__32454;
    wire N__32451;
    wire N__32450;
    wire N__32449;
    wire N__32446;
    wire N__32443;
    wire N__32440;
    wire N__32437;
    wire N__32436;
    wire N__32435;
    wire N__32432;
    wire N__32431;
    wire N__32430;
    wire N__32427;
    wire N__32424;
    wire N__32423;
    wire N__32420;
    wire N__32419;
    wire N__32416;
    wire N__32413;
    wire N__32412;
    wire N__32411;
    wire N__32408;
    wire N__32407;
    wire N__32406;
    wire N__32403;
    wire N__32402;
    wire N__32401;
    wire N__32398;
    wire N__32397;
    wire N__32392;
    wire N__32389;
    wire N__32386;
    wire N__32385;
    wire N__32384;
    wire N__32381;
    wire N__32380;
    wire N__32377;
    wire N__32372;
    wire N__32369;
    wire N__32366;
    wire N__32363;
    wire N__32360;
    wire N__32357;
    wire N__32356;
    wire N__32355;
    wire N__32354;
    wire N__32351;
    wire N__32350;
    wire N__32349;
    wire N__32346;
    wire N__32343;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32335;
    wire N__32334;
    wire N__32333;
    wire N__32332;
    wire N__32329;
    wire N__32326;
    wire N__32323;
    wire N__32322;
    wire N__32319;
    wire N__32318;
    wire N__32317;
    wire N__32316;
    wire N__32313;
    wire N__32310;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32299;
    wire N__32296;
    wire N__32293;
    wire N__32290;
    wire N__32285;
    wire N__32284;
    wire N__32283;
    wire N__32282;
    wire N__32281;
    wire N__32280;
    wire N__32279;
    wire N__32276;
    wire N__32273;
    wire N__32270;
    wire N__32269;
    wire N__32266;
    wire N__32265;
    wire N__32262;
    wire N__32261;
    wire N__32252;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32236;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32228;
    wire N__32227;
    wire N__32226;
    wire N__32225;
    wire N__32224;
    wire N__32221;
    wire N__32220;
    wire N__32215;
    wire N__32212;
    wire N__32207;
    wire N__32206;
    wire N__32205;
    wire N__32202;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32184;
    wire N__32181;
    wire N__32180;
    wire N__32179;
    wire N__32176;
    wire N__32173;
    wire N__32170;
    wire N__32167;
    wire N__32166;
    wire N__32161;
    wire N__32158;
    wire N__32155;
    wire N__32150;
    wire N__32147;
    wire N__32144;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32127;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32112;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32083;
    wire N__32080;
    wire N__32075;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32060;
    wire N__32057;
    wire N__32054;
    wire N__32053;
    wire N__32052;
    wire N__32047;
    wire N__32046;
    wire N__32045;
    wire N__32042;
    wire N__32039;
    wire N__32036;
    wire N__32033;
    wire N__32030;
    wire N__32025;
    wire N__32022;
    wire N__32017;
    wire N__32014;
    wire N__32011;
    wire N__32008;
    wire N__32003;
    wire N__32000;
    wire N__31997;
    wire N__31994;
    wire N__31991;
    wire N__31988;
    wire N__31981;
    wire N__31968;
    wire N__31965;
    wire N__31958;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31936;
    wire N__31925;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31906;
    wire N__31903;
    wire N__31896;
    wire N__31891;
    wire N__31886;
    wire N__31877;
    wire N__31868;
    wire N__31863;
    wire N__31856;
    wire N__31851;
    wire N__31846;
    wire N__31837;
    wire N__31836;
    wire N__31833;
    wire N__31826;
    wire N__31821;
    wire N__31814;
    wire N__31807;
    wire N__31802;
    wire N__31799;
    wire N__31794;
    wire N__31781;
    wire N__31780;
    wire N__31777;
    wire N__31774;
    wire N__31773;
    wire N__31772;
    wire N__31771;
    wire N__31768;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31757;
    wire N__31756;
    wire N__31755;
    wire N__31754;
    wire N__31751;
    wire N__31750;
    wire N__31747;
    wire N__31744;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31722;
    wire N__31721;
    wire N__31718;
    wire N__31715;
    wire N__31710;
    wire N__31707;
    wire N__31700;
    wire N__31697;
    wire N__31694;
    wire N__31691;
    wire N__31688;
    wire N__31685;
    wire N__31680;
    wire N__31677;
    wire N__31672;
    wire N__31669;
    wire N__31664;
    wire N__31657;
    wire N__31654;
    wire N__31651;
    wire N__31644;
    wire N__31637;
    wire N__31634;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31622;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31603;
    wire N__31600;
    wire N__31595;
    wire N__31592;
    wire N__31591;
    wire N__31590;
    wire N__31589;
    wire N__31588;
    wire N__31587;
    wire N__31586;
    wire N__31585;
    wire N__31584;
    wire N__31583;
    wire N__31582;
    wire N__31581;
    wire N__31580;
    wire N__31579;
    wire N__31576;
    wire N__31575;
    wire N__31572;
    wire N__31569;
    wire N__31568;
    wire N__31567;
    wire N__31566;
    wire N__31565;
    wire N__31564;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31545;
    wire N__31540;
    wire N__31535;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31508;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31498;
    wire N__31497;
    wire N__31488;
    wire N__31479;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31460;
    wire N__31453;
    wire N__31442;
    wire N__31439;
    wire N__31436;
    wire N__31435;
    wire N__31434;
    wire N__31433;
    wire N__31432;
    wire N__31431;
    wire N__31430;
    wire N__31427;
    wire N__31426;
    wire N__31425;
    wire N__31424;
    wire N__31423;
    wire N__31422;
    wire N__31421;
    wire N__31418;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31406;
    wire N__31405;
    wire N__31402;
    wire N__31401;
    wire N__31400;
    wire N__31399;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31385;
    wire N__31380;
    wire N__31377;
    wire N__31374;
    wire N__31369;
    wire N__31358;
    wire N__31353;
    wire N__31348;
    wire N__31345;
    wire N__31340;
    wire N__31337;
    wire N__31322;
    wire N__31321;
    wire N__31318;
    wire N__31315;
    wire N__31314;
    wire N__31311;
    wire N__31310;
    wire N__31309;
    wire N__31308;
    wire N__31307;
    wire N__31306;
    wire N__31305;
    wire N__31302;
    wire N__31299;
    wire N__31298;
    wire N__31297;
    wire N__31294;
    wire N__31291;
    wire N__31288;
    wire N__31285;
    wire N__31282;
    wire N__31277;
    wire N__31276;
    wire N__31273;
    wire N__31270;
    wire N__31265;
    wire N__31264;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31252;
    wire N__31249;
    wire N__31248;
    wire N__31247;
    wire N__31244;
    wire N__31241;
    wire N__31238;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31222;
    wire N__31217;
    wire N__31212;
    wire N__31199;
    wire N__31190;
    wire N__31187;
    wire N__31186;
    wire N__31183;
    wire N__31180;
    wire N__31177;
    wire N__31174;
    wire N__31169;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31153;
    wire N__31152;
    wire N__31151;
    wire N__31150;
    wire N__31149;
    wire N__31148;
    wire N__31147;
    wire N__31146;
    wire N__31145;
    wire N__31144;
    wire N__31141;
    wire N__31140;
    wire N__31133;
    wire N__31128;
    wire N__31123;
    wire N__31122;
    wire N__31119;
    wire N__31116;
    wire N__31109;
    wire N__31106;
    wire N__31105;
    wire N__31104;
    wire N__31103;
    wire N__31102;
    wire N__31097;
    wire N__31094;
    wire N__31091;
    wire N__31090;
    wire N__31089;
    wire N__31088;
    wire N__31087;
    wire N__31084;
    wire N__31079;
    wire N__31076;
    wire N__31069;
    wire N__31064;
    wire N__31061;
    wire N__31056;
    wire N__31051;
    wire N__31046;
    wire N__31039;
    wire N__31028;
    wire N__31025;
    wire N__31024;
    wire N__31023;
    wire N__31022;
    wire N__31021;
    wire N__31020;
    wire N__31019;
    wire N__31018;
    wire N__31015;
    wire N__31014;
    wire N__31013;
    wire N__31010;
    wire N__31007;
    wire N__31004;
    wire N__31003;
    wire N__31002;
    wire N__30999;
    wire N__30994;
    wire N__30991;
    wire N__30988;
    wire N__30983;
    wire N__30982;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30968;
    wire N__30963;
    wire N__30960;
    wire N__30955;
    wire N__30950;
    wire N__30945;
    wire N__30938;
    wire N__30929;
    wire N__30928;
    wire N__30927;
    wire N__30926;
    wire N__30925;
    wire N__30924;
    wire N__30921;
    wire N__30920;
    wire N__30919;
    wire N__30918;
    wire N__30917;
    wire N__30916;
    wire N__30913;
    wire N__30906;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30893;
    wire N__30886;
    wire N__30883;
    wire N__30880;
    wire N__30875;
    wire N__30872;
    wire N__30867;
    wire N__30864;
    wire N__30857;
    wire N__30848;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30836;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30824;
    wire N__30821;
    wire N__30818;
    wire N__30815;
    wire N__30812;
    wire N__30811;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30799;
    wire N__30796;
    wire N__30793;
    wire N__30788;
    wire N__30785;
    wire N__30784;
    wire N__30783;
    wire N__30782;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30770;
    wire N__30769;
    wire N__30766;
    wire N__30759;
    wire N__30756;
    wire N__30751;
    wire N__30748;
    wire N__30745;
    wire N__30740;
    wire N__30739;
    wire N__30738;
    wire N__30737;
    wire N__30736;
    wire N__30735;
    wire N__30734;
    wire N__30733;
    wire N__30732;
    wire N__30729;
    wire N__30728;
    wire N__30727;
    wire N__30724;
    wire N__30723;
    wire N__30722;
    wire N__30721;
    wire N__30720;
    wire N__30713;
    wire N__30710;
    wire N__30709;
    wire N__30708;
    wire N__30707;
    wire N__30706;
    wire N__30705;
    wire N__30700;
    wire N__30697;
    wire N__30696;
    wire N__30695;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30676;
    wire N__30673;
    wire N__30672;
    wire N__30671;
    wire N__30670;
    wire N__30667;
    wire N__30666;
    wire N__30665;
    wire N__30664;
    wire N__30659;
    wire N__30656;
    wire N__30647;
    wire N__30642;
    wire N__30639;
    wire N__30634;
    wire N__30629;
    wire N__30626;
    wire N__30619;
    wire N__30612;
    wire N__30609;
    wire N__30606;
    wire N__30603;
    wire N__30602;
    wire N__30599;
    wire N__30598;
    wire N__30595;
    wire N__30588;
    wire N__30581;
    wire N__30580;
    wire N__30579;
    wire N__30578;
    wire N__30577;
    wire N__30576;
    wire N__30575;
    wire N__30572;
    wire N__30569;
    wire N__30564;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30550;
    wire N__30545;
    wire N__30540;
    wire N__30533;
    wire N__30526;
    wire N__30521;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30501;
    wire N__30498;
    wire N__30493;
    wire N__30488;
    wire N__30485;
    wire N__30482;
    wire N__30477;
    wire N__30470;
    wire N__30469;
    wire N__30464;
    wire N__30461;
    wire N__30458;
    wire N__30455;
    wire N__30452;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30442;
    wire N__30437;
    wire N__30434;
    wire N__30433;
    wire N__30428;
    wire N__30425;
    wire N__30422;
    wire N__30421;
    wire N__30420;
    wire N__30417;
    wire N__30416;
    wire N__30415;
    wire N__30414;
    wire N__30413;
    wire N__30412;
    wire N__30411;
    wire N__30410;
    wire N__30409;
    wire N__30402;
    wire N__30395;
    wire N__30390;
    wire N__30389;
    wire N__30388;
    wire N__30387;
    wire N__30384;
    wire N__30381;
    wire N__30378;
    wire N__30377;
    wire N__30374;
    wire N__30369;
    wire N__30364;
    wire N__30355;
    wire N__30354;
    wire N__30353;
    wire N__30352;
    wire N__30349;
    wire N__30348;
    wire N__30347;
    wire N__30346;
    wire N__30337;
    wire N__30332;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30318;
    wire N__30317;
    wire N__30316;
    wire N__30315;
    wire N__30314;
    wire N__30311;
    wire N__30306;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30289;
    wire N__30288;
    wire N__30285;
    wire N__30284;
    wire N__30281;
    wire N__30274;
    wire N__30267;
    wire N__30266;
    wire N__30265;
    wire N__30264;
    wire N__30259;
    wire N__30258;
    wire N__30255;
    wire N__30248;
    wire N__30245;
    wire N__30244;
    wire N__30243;
    wire N__30240;
    wire N__30239;
    wire N__30236;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30228;
    wire N__30227;
    wire N__30224;
    wire N__30221;
    wire N__30218;
    wire N__30213;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30197;
    wire N__30192;
    wire N__30189;
    wire N__30186;
    wire N__30177;
    wire N__30174;
    wire N__30169;
    wire N__30158;
    wire N__30157;
    wire N__30154;
    wire N__30153;
    wire N__30152;
    wire N__30151;
    wire N__30150;
    wire N__30149;
    wire N__30148;
    wire N__30147;
    wire N__30146;
    wire N__30145;
    wire N__30144;
    wire N__30143;
    wire N__30134;
    wire N__30129;
    wire N__30126;
    wire N__30125;
    wire N__30124;
    wire N__30123;
    wire N__30122;
    wire N__30119;
    wire N__30118;
    wire N__30117;
    wire N__30116;
    wire N__30115;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30096;
    wire N__30091;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30079;
    wire N__30076;
    wire N__30075;
    wire N__30074;
    wire N__30073;
    wire N__30070;
    wire N__30065;
    wire N__30062;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30050;
    wire N__30049;
    wire N__30046;
    wire N__30037;
    wire N__30032;
    wire N__30029;
    wire N__30026;
    wire N__30023;
    wire N__30022;
    wire N__30019;
    wire N__30018;
    wire N__30015;
    wire N__30014;
    wire N__30013;
    wire N__30012;
    wire N__30005;
    wire N__30002;
    wire N__29997;
    wire N__29994;
    wire N__29991;
    wire N__29982;
    wire N__29981;
    wire N__29980;
    wire N__29977;
    wire N__29974;
    wire N__29969;
    wire N__29966;
    wire N__29963;
    wire N__29960;
    wire N__29955;
    wire N__29946;
    wire N__29941;
    wire N__29936;
    wire N__29915;
    wire N__29914;
    wire N__29913;
    wire N__29912;
    wire N__29909;
    wire N__29904;
    wire N__29901;
    wire N__29900;
    wire N__29899;
    wire N__29898;
    wire N__29897;
    wire N__29896;
    wire N__29895;
    wire N__29894;
    wire N__29893;
    wire N__29892;
    wire N__29889;
    wire N__29886;
    wire N__29881;
    wire N__29876;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29862;
    wire N__29859;
    wire N__29848;
    wire N__29845;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29833;
    wire N__29830;
    wire N__29827;
    wire N__29820;
    wire N__29813;
    wire N__29812;
    wire N__29809;
    wire N__29806;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29780;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29765;
    wire N__29762;
    wire N__29759;
    wire N__29758;
    wire N__29757;
    wire N__29754;
    wire N__29749;
    wire N__29748;
    wire N__29745;
    wire N__29744;
    wire N__29743;
    wire N__29742;
    wire N__29739;
    wire N__29736;
    wire N__29733;
    wire N__29730;
    wire N__29727;
    wire N__29726;
    wire N__29725;
    wire N__29722;
    wire N__29717;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29699;
    wire N__29694;
    wire N__29691;
    wire N__29688;
    wire N__29683;
    wire N__29680;
    wire N__29669;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29656;
    wire N__29655;
    wire N__29654;
    wire N__29651;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29626;
    wire N__29623;
    wire N__29620;
    wire N__29619;
    wire N__29618;
    wire N__29617;
    wire N__29614;
    wire N__29611;
    wire N__29610;
    wire N__29609;
    wire N__29608;
    wire N__29605;
    wire N__29604;
    wire N__29601;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29586;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29573;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29559;
    wire N__29558;
    wire N__29557;
    wire N__29554;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29537;
    wire N__29536;
    wire N__29533;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29521;
    wire N__29518;
    wire N__29511;
    wire N__29506;
    wire N__29489;
    wire N__29486;
    wire N__29485;
    wire N__29484;
    wire N__29481;
    wire N__29476;
    wire N__29471;
    wire N__29470;
    wire N__29467;
    wire N__29462;
    wire N__29459;
    wire N__29456;
    wire N__29455;
    wire N__29452;
    wire N__29449;
    wire N__29446;
    wire N__29443;
    wire N__29442;
    wire N__29437;
    wire N__29434;
    wire N__29429;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29408;
    wire N__29405;
    wire N__29402;
    wire N__29399;
    wire N__29396;
    wire N__29395;
    wire N__29390;
    wire N__29389;
    wire N__29388;
    wire N__29385;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29369;
    wire N__29366;
    wire N__29365;
    wire N__29364;
    wire N__29361;
    wire N__29356;
    wire N__29355;
    wire N__29352;
    wire N__29349;
    wire N__29346;
    wire N__29339;
    wire N__29336;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29317;
    wire N__29312;
    wire N__29309;
    wire N__29308;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29293;
    wire N__29292;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29276;
    wire N__29275;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29267;
    wire N__29264;
    wire N__29261;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29240;
    wire N__29231;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29223;
    wire N__29222;
    wire N__29219;
    wire N__29216;
    wire N__29213;
    wire N__29210;
    wire N__29209;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29187;
    wire N__29180;
    wire N__29177;
    wire N__29174;
    wire N__29173;
    wire N__29170;
    wire N__29167;
    wire N__29162;
    wire N__29161;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29135;
    wire N__29134;
    wire N__29133;
    wire N__29126;
    wire N__29123;
    wire N__29120;
    wire N__29119;
    wire N__29118;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29110;
    wire N__29107;
    wire N__29106;
    wire N__29105;
    wire N__29104;
    wire N__29103;
    wire N__29100;
    wire N__29099;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29082;
    wire N__29081;
    wire N__29080;
    wire N__29077;
    wire N__29076;
    wire N__29075;
    wire N__29074;
    wire N__29071;
    wire N__29070;
    wire N__29069;
    wire N__29066;
    wire N__29063;
    wire N__29062;
    wire N__29061;
    wire N__29060;
    wire N__29057;
    wire N__29052;
    wire N__29047;
    wire N__29040;
    wire N__29039;
    wire N__29038;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29007;
    wire N__29000;
    wire N__28997;
    wire N__28992;
    wire N__28991;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28977;
    wire N__28970;
    wire N__28961;
    wire N__28956;
    wire N__28943;
    wire N__28940;
    wire N__28939;
    wire N__28934;
    wire N__28931;
    wire N__28928;
    wire N__28925;
    wire N__28924;
    wire N__28923;
    wire N__28920;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28885;
    wire N__28882;
    wire N__28877;
    wire N__28874;
    wire N__28873;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28849;
    wire N__28848;
    wire N__28847;
    wire N__28846;
    wire N__28845;
    wire N__28844;
    wire N__28843;
    wire N__28842;
    wire N__28841;
    wire N__28836;
    wire N__28833;
    wire N__28832;
    wire N__28829;
    wire N__28824;
    wire N__28817;
    wire N__28816;
    wire N__28815;
    wire N__28814;
    wire N__28813;
    wire N__28810;
    wire N__28805;
    wire N__28802;
    wire N__28801;
    wire N__28800;
    wire N__28797;
    wire N__28792;
    wire N__28791;
    wire N__28790;
    wire N__28787;
    wire N__28782;
    wire N__28779;
    wire N__28772;
    wire N__28767;
    wire N__28762;
    wire N__28757;
    wire N__28754;
    wire N__28739;
    wire N__28736;
    wire N__28733;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28717;
    wire N__28716;
    wire N__28715;
    wire N__28714;
    wire N__28711;
    wire N__28702;
    wire N__28697;
    wire N__28696;
    wire N__28695;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28681;
    wire N__28676;
    wire N__28673;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28648;
    wire N__28645;
    wire N__28642;
    wire N__28637;
    wire N__28634;
    wire N__28631;
    wire N__28628;
    wire N__28625;
    wire N__28624;
    wire N__28623;
    wire N__28618;
    wire N__28615;
    wire N__28612;
    wire N__28609;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28597;
    wire N__28594;
    wire N__28591;
    wire N__28590;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28574;
    wire N__28571;
    wire N__28568;
    wire N__28565;
    wire N__28562;
    wire N__28559;
    wire N__28556;
    wire N__28553;
    wire N__28552;
    wire N__28551;
    wire N__28550;
    wire N__28549;
    wire N__28548;
    wire N__28547;
    wire N__28546;
    wire N__28545;
    wire N__28544;
    wire N__28543;
    wire N__28542;
    wire N__28541;
    wire N__28540;
    wire N__28533;
    wire N__28524;
    wire N__28523;
    wire N__28522;
    wire N__28521;
    wire N__28520;
    wire N__28517;
    wire N__28516;
    wire N__28509;
    wire N__28502;
    wire N__28497;
    wire N__28484;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28466;
    wire N__28463;
    wire N__28460;
    wire N__28459;
    wire N__28456;
    wire N__28453;
    wire N__28448;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28429;
    wire N__28428;
    wire N__28425;
    wire N__28420;
    wire N__28415;
    wire N__28414;
    wire N__28409;
    wire N__28406;
    wire N__28403;
    wire N__28400;
    wire N__28397;
    wire N__28394;
    wire N__28393;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28381;
    wire N__28378;
    wire N__28377;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28358;
    wire N__28357;
    wire N__28352;
    wire N__28349;
    wire N__28346;
    wire N__28345;
    wire N__28344;
    wire N__28339;
    wire N__28336;
    wire N__28331;
    wire N__28330;
    wire N__28325;
    wire N__28322;
    wire N__28319;
    wire N__28318;
    wire N__28315;
    wire N__28314;
    wire N__28311;
    wire N__28310;
    wire N__28307;
    wire N__28304;
    wire N__28301;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28277;
    wire N__28274;
    wire N__28265;
    wire N__28264;
    wire N__28259;
    wire N__28256;
    wire N__28253;
    wire N__28250;
    wire N__28247;
    wire N__28246;
    wire N__28245;
    wire N__28242;
    wire N__28237;
    wire N__28234;
    wire N__28229;
    wire N__28228;
    wire N__28223;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28213;
    wire N__28210;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28193;
    wire N__28190;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28178;
    wire N__28175;
    wire N__28172;
    wire N__28169;
    wire N__28168;
    wire N__28163;
    wire N__28160;
    wire N__28157;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28147;
    wire N__28142;
    wire N__28139;
    wire N__28136;
    wire N__28133;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28120;
    wire N__28117;
    wire N__28112;
    wire N__28111;
    wire N__28110;
    wire N__28107;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28091;
    wire N__28088;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28075;
    wire N__28072;
    wire N__28071;
    wire N__28070;
    wire N__28067;
    wire N__28064;
    wire N__28059;
    wire N__28056;
    wire N__28049;
    wire N__28046;
    wire N__28045;
    wire N__28044;
    wire N__28041;
    wire N__28036;
    wire N__28033;
    wire N__28028;
    wire N__28027;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__28003;
    wire N__28002;
    wire N__27995;
    wire N__27992;
    wire N__27989;
    wire N__27988;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27961;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27938;
    wire N__27935;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27913;
    wire N__27908;
    wire N__27905;
    wire N__27902;
    wire N__27901;
    wire N__27898;
    wire N__27897;
    wire N__27894;
    wire N__27893;
    wire N__27892;
    wire N__27891;
    wire N__27886;
    wire N__27881;
    wire N__27880;
    wire N__27879;
    wire N__27878;
    wire N__27875;
    wire N__27872;
    wire N__27867;
    wire N__27862;
    wire N__27861;
    wire N__27856;
    wire N__27849;
    wire N__27846;
    wire N__27841;
    wire N__27836;
    wire N__27835;
    wire N__27834;
    wire N__27833;
    wire N__27832;
    wire N__27831;
    wire N__27826;
    wire N__27825;
    wire N__27820;
    wire N__27819;
    wire N__27814;
    wire N__27811;
    wire N__27810;
    wire N__27807;
    wire N__27804;
    wire N__27801;
    wire N__27798;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27779;
    wire N__27770;
    wire N__27769;
    wire N__27768;
    wire N__27767;
    wire N__27764;
    wire N__27763;
    wire N__27756;
    wire N__27755;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27747;
    wire N__27746;
    wire N__27745;
    wire N__27744;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27726;
    wire N__27721;
    wire N__27716;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27692;
    wire N__27689;
    wire N__27688;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27677;
    wire N__27674;
    wire N__27673;
    wire N__27672;
    wire N__27667;
    wire N__27666;
    wire N__27665;
    wire N__27664;
    wire N__27663;
    wire N__27660;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27644;
    wire N__27641;
    wire N__27640;
    wire N__27637;
    wire N__27634;
    wire N__27631;
    wire N__27626;
    wire N__27625;
    wire N__27624;
    wire N__27623;
    wire N__27622;
    wire N__27621;
    wire N__27618;
    wire N__27617;
    wire N__27612;
    wire N__27609;
    wire N__27600;
    wire N__27595;
    wire N__27590;
    wire N__27583;
    wire N__27582;
    wire N__27579;
    wire N__27576;
    wire N__27575;
    wire N__27574;
    wire N__27569;
    wire N__27566;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27546;
    wire N__27543;
    wire N__27538;
    wire N__27535;
    wire N__27524;
    wire N__27521;
    wire N__27520;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27512;
    wire N__27511;
    wire N__27510;
    wire N__27507;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27497;
    wire N__27492;
    wire N__27487;
    wire N__27476;
    wire N__27475;
    wire N__27472;
    wire N__27467;
    wire N__27464;
    wire N__27461;
    wire N__27460;
    wire N__27459;
    wire N__27458;
    wire N__27457;
    wire N__27456;
    wire N__27453;
    wire N__27452;
    wire N__27451;
    wire N__27446;
    wire N__27443;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27401;
    wire N__27396;
    wire N__27391;
    wire N__27388;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27376;
    wire N__27375;
    wire N__27374;
    wire N__27373;
    wire N__27372;
    wire N__27371;
    wire N__27370;
    wire N__27369;
    wire N__27368;
    wire N__27365;
    wire N__27364;
    wire N__27361;
    wire N__27360;
    wire N__27359;
    wire N__27356;
    wire N__27355;
    wire N__27354;
    wire N__27347;
    wire N__27346;
    wire N__27345;
    wire N__27344;
    wire N__27343;
    wire N__27342;
    wire N__27341;
    wire N__27340;
    wire N__27337;
    wire N__27328;
    wire N__27325;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27307;
    wire N__27302;
    wire N__27299;
    wire N__27290;
    wire N__27287;
    wire N__27280;
    wire N__27275;
    wire N__27260;
    wire N__27257;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27247;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27235;
    wire N__27234;
    wire N__27229;
    wire N__27228;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27206;
    wire N__27205;
    wire N__27202;
    wire N__27197;
    wire N__27192;
    wire N__27185;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27177;
    wire N__27176;
    wire N__27175;
    wire N__27174;
    wire N__27173;
    wire N__27172;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27160;
    wire N__27157;
    wire N__27152;
    wire N__27151;
    wire N__27146;
    wire N__27141;
    wire N__27138;
    wire N__27133;
    wire N__27130;
    wire N__27127;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27107;
    wire N__27106;
    wire N__27105;
    wire N__27104;
    wire N__27103;
    wire N__27100;
    wire N__27099;
    wire N__27098;
    wire N__27097;
    wire N__27096;
    wire N__27093;
    wire N__27090;
    wire N__27089;
    wire N__27086;
    wire N__27085;
    wire N__27082;
    wire N__27079;
    wire N__27076;
    wire N__27075;
    wire N__27074;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27066;
    wire N__27065;
    wire N__27058;
    wire N__27051;
    wire N__27046;
    wire N__27043;
    wire N__27040;
    wire N__27033;
    wire N__27028;
    wire N__27025;
    wire N__27020;
    wire N__27015;
    wire N__27004;
    wire N__26999;
    wire N__26996;
    wire N__26993;
    wire N__26992;
    wire N__26989;
    wire N__26986;
    wire N__26981;
    wire N__26978;
    wire N__26977;
    wire N__26976;
    wire N__26975;
    wire N__26974;
    wire N__26973;
    wire N__26970;
    wire N__26969;
    wire N__26968;
    wire N__26967;
    wire N__26964;
    wire N__26963;
    wire N__26956;
    wire N__26953;
    wire N__26952;
    wire N__26949;
    wire N__26942;
    wire N__26939;
    wire N__26936;
    wire N__26931;
    wire N__26928;
    wire N__26923;
    wire N__26920;
    wire N__26909;
    wire N__26906;
    wire N__26903;
    wire N__26900;
    wire N__26897;
    wire N__26894;
    wire N__26891;
    wire N__26888;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26870;
    wire N__26869;
    wire N__26864;
    wire N__26861;
    wire N__26858;
    wire N__26855;
    wire N__26852;
    wire N__26851;
    wire N__26846;
    wire N__26843;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26824;
    wire N__26823;
    wire N__26822;
    wire N__26821;
    wire N__26820;
    wire N__26817;
    wire N__26806;
    wire N__26805;
    wire N__26804;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26770;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26755;
    wire N__26754;
    wire N__26753;
    wire N__26752;
    wire N__26749;
    wire N__26748;
    wire N__26747;
    wire N__26746;
    wire N__26745;
    wire N__26744;
    wire N__26743;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26735;
    wire N__26734;
    wire N__26731;
    wire N__26728;
    wire N__26721;
    wire N__26718;
    wire N__26715;
    wire N__26710;
    wire N__26709;
    wire N__26708;
    wire N__26707;
    wire N__26704;
    wire N__26701;
    wire N__26694;
    wire N__26691;
    wire N__26682;
    wire N__26679;
    wire N__26676;
    wire N__26671;
    wire N__26668;
    wire N__26663;
    wire N__26658;
    wire N__26651;
    wire N__26648;
    wire N__26645;
    wire N__26640;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26585;
    wire N__26582;
    wire N__26579;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26557;
    wire N__26554;
    wire N__26553;
    wire N__26552;
    wire N__26549;
    wire N__26548;
    wire N__26547;
    wire N__26544;
    wire N__26541;
    wire N__26540;
    wire N__26537;
    wire N__26532;
    wire N__26529;
    wire N__26526;
    wire N__26523;
    wire N__26522;
    wire N__26519;
    wire N__26516;
    wire N__26513;
    wire N__26510;
    wire N__26509;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26489;
    wire N__26484;
    wire N__26471;
    wire N__26470;
    wire N__26467;
    wire N__26462;
    wire N__26459;
    wire N__26458;
    wire N__26457;
    wire N__26456;
    wire N__26455;
    wire N__26454;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26446;
    wire N__26441;
    wire N__26436;
    wire N__26431;
    wire N__26426;
    wire N__26425;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26405;
    wire N__26404;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26386;
    wire N__26385;
    wire N__26384;
    wire N__26383;
    wire N__26380;
    wire N__26377;
    wire N__26372;
    wire N__26371;
    wire N__26368;
    wire N__26367;
    wire N__26366;
    wire N__26365;
    wire N__26358;
    wire N__26353;
    wire N__26350;
    wire N__26349;
    wire N__26346;
    wire N__26343;
    wire N__26342;
    wire N__26339;
    wire N__26334;
    wire N__26331;
    wire N__26328;
    wire N__26325;
    wire N__26322;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26293;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26281;
    wire N__26280;
    wire N__26277;
    wire N__26276;
    wire N__26275;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26261;
    wire N__26256;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26240;
    wire N__26239;
    wire N__26236;
    wire N__26235;
    wire N__26232;
    wire N__26231;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26210;
    wire N__26205;
    wire N__26200;
    wire N__26197;
    wire N__26192;
    wire N__26191;
    wire N__26186;
    wire N__26183;
    wire N__26180;
    wire N__26179;
    wire N__26176;
    wire N__26175;
    wire N__26174;
    wire N__26171;
    wire N__26164;
    wire N__26161;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26147;
    wire N__26144;
    wire N__26141;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26131;
    wire N__26130;
    wire N__26129;
    wire N__26128;
    wire N__26127;
    wire N__26126;
    wire N__26125;
    wire N__26124;
    wire N__26123;
    wire N__26122;
    wire N__26121;
    wire N__26120;
    wire N__26119;
    wire N__26114;
    wire N__26107;
    wire N__26102;
    wire N__26101;
    wire N__26100;
    wire N__26099;
    wire N__26098;
    wire N__26097;
    wire N__26096;
    wire N__26087;
    wire N__26080;
    wire N__26077;
    wire N__26072;
    wire N__26059;
    wire N__26056;
    wire N__26053;
    wire N__26046;
    wire N__26041;
    wire N__26038;
    wire N__26033;
    wire N__26030;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26020;
    wire N__26015;
    wire N__26014;
    wire N__26011;
    wire N__26010;
    wire N__26007;
    wire N__26004;
    wire N__25999;
    wire N__25996;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25978;
    wire N__25973;
    wire N__25970;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25960;
    wire N__25957;
    wire N__25954;
    wire N__25951;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25925;
    wire N__25922;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25892;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25873;
    wire N__25872;
    wire N__25871;
    wire N__25868;
    wire N__25867;
    wire N__25866;
    wire N__25865;
    wire N__25864;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25847;
    wire N__25844;
    wire N__25839;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25823;
    wire N__25820;
    wire N__25817;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25801;
    wire N__25800;
    wire N__25797;
    wire N__25794;
    wire N__25791;
    wire N__25786;
    wire N__25783;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25756;
    wire N__25755;
    wire N__25754;
    wire N__25753;
    wire N__25752;
    wire N__25751;
    wire N__25750;
    wire N__25749;
    wire N__25748;
    wire N__25747;
    wire N__25746;
    wire N__25745;
    wire N__25744;
    wire N__25743;
    wire N__25742;
    wire N__25741;
    wire N__25740;
    wire N__25739;
    wire N__25738;
    wire N__25737;
    wire N__25736;
    wire N__25735;
    wire N__25734;
    wire N__25733;
    wire N__25732;
    wire N__25727;
    wire N__25718;
    wire N__25709;
    wire N__25702;
    wire N__25699;
    wire N__25698;
    wire N__25697;
    wire N__25694;
    wire N__25687;
    wire N__25684;
    wire N__25673;
    wire N__25668;
    wire N__25659;
    wire N__25658;
    wire N__25657;
    wire N__25656;
    wire N__25655;
    wire N__25648;
    wire N__25635;
    wire N__25634;
    wire N__25631;
    wire N__25624;
    wire N__25621;
    wire N__25620;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25605;
    wire N__25600;
    wire N__25595;
    wire N__25586;
    wire N__25583;
    wire N__25582;
    wire N__25581;
    wire N__25580;
    wire N__25579;
    wire N__25578;
    wire N__25577;
    wire N__25574;
    wire N__25569;
    wire N__25566;
    wire N__25561;
    wire N__25558;
    wire N__25553;
    wire N__25544;
    wire N__25543;
    wire N__25540;
    wire N__25537;
    wire N__25534;
    wire N__25529;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25516;
    wire N__25513;
    wire N__25510;
    wire N__25507;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25478;
    wire N__25475;
    wire N__25472;
    wire N__25471;
    wire N__25468;
    wire N__25465;
    wire N__25462;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25450;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25436;
    wire N__25433;
    wire N__25432;
    wire N__25431;
    wire N__25430;
    wire N__25429;
    wire N__25428;
    wire N__25427;
    wire N__25426;
    wire N__25425;
    wire N__25424;
    wire N__25423;
    wire N__25422;
    wire N__25421;
    wire N__25420;
    wire N__25419;
    wire N__25418;
    wire N__25417;
    wire N__25416;
    wire N__25415;
    wire N__25414;
    wire N__25413;
    wire N__25412;
    wire N__25411;
    wire N__25410;
    wire N__25409;
    wire N__25408;
    wire N__25407;
    wire N__25406;
    wire N__25405;
    wire N__25404;
    wire N__25403;
    wire N__25402;
    wire N__25401;
    wire N__25400;
    wire N__25399;
    wire N__25390;
    wire N__25381;
    wire N__25372;
    wire N__25363;
    wire N__25356;
    wire N__25347;
    wire N__25340;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25320;
    wire N__25317;
    wire N__25316;
    wire N__25315;
    wire N__25314;
    wire N__25313;
    wire N__25312;
    wire N__25311;
    wire N__25310;
    wire N__25309;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25287;
    wire N__25284;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25272;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25213;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25195;
    wire N__25194;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25183;
    wire N__25182;
    wire N__25181;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25113;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25097;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25069;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25055;
    wire N__25052;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25042;
    wire N__25037;
    wire N__25034;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25024;
    wire N__25019;
    wire N__25016;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25001;
    wire N__24998;
    wire N__24997;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24983;
    wire N__24980;
    wire N__24979;
    wire N__24976;
    wire N__24973;
    wire N__24970;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24944;
    wire N__24941;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24926;
    wire N__24923;
    wire N__24920;
    wire N__24919;
    wire N__24914;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24904;
    wire N__24899;
    wire N__24896;
    wire N__24893;
    wire N__24890;
    wire N__24887;
    wire N__24886;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24859;
    wire N__24858;
    wire N__24857;
    wire N__24856;
    wire N__24853;
    wire N__24850;
    wire N__24843;
    wire N__24840;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24814;
    wire N__24813;
    wire N__24810;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24796;
    wire N__24795;
    wire N__24794;
    wire N__24793;
    wire N__24790;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24778;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24768;
    wire N__24767;
    wire N__24762;
    wire N__24757;
    wire N__24750;
    wire N__24749;
    wire N__24748;
    wire N__24747;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24732;
    wire N__24729;
    wire N__24720;
    wire N__24707;
    wire N__24706;
    wire N__24705;
    wire N__24704;
    wire N__24703;
    wire N__24702;
    wire N__24701;
    wire N__24700;
    wire N__24697;
    wire N__24696;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24682;
    wire N__24679;
    wire N__24678;
    wire N__24677;
    wire N__24676;
    wire N__24673;
    wire N__24670;
    wire N__24665;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24649;
    wire N__24646;
    wire N__24637;
    wire N__24634;
    wire N__24623;
    wire N__24620;
    wire N__24619;
    wire N__24618;
    wire N__24615;
    wire N__24614;
    wire N__24613;
    wire N__24612;
    wire N__24609;
    wire N__24608;
    wire N__24607;
    wire N__24606;
    wire N__24605;
    wire N__24604;
    wire N__24603;
    wire N__24600;
    wire N__24599;
    wire N__24596;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24582;
    wire N__24579;
    wire N__24574;
    wire N__24569;
    wire N__24564;
    wire N__24557;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24512;
    wire N__24509;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24499;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24476;
    wire N__24473;
    wire N__24472;
    wire N__24469;
    wire N__24468;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24456;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24442;
    wire N__24441;
    wire N__24438;
    wire N__24435;
    wire N__24434;
    wire N__24431;
    wire N__24428;
    wire N__24427;
    wire N__24426;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24397;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24376;
    wire N__24371;
    wire N__24368;
    wire N__24365;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24353;
    wire N__24350;
    wire N__24349;
    wire N__24348;
    wire N__24345;
    wire N__24340;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24314;
    wire N__24313;
    wire N__24310;
    wire N__24307;
    wire N__24302;
    wire N__24299;
    wire N__24298;
    wire N__24295;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24281;
    wire N__24278;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24224;
    wire N__24223;
    wire N__24222;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24187;
    wire N__24182;
    wire N__24179;
    wire N__24176;
    wire N__24175;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24163;
    wire N__24158;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24136;
    wire N__24131;
    wire N__24128;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24116;
    wire N__24115;
    wire N__24114;
    wire N__24113;
    wire N__24112;
    wire N__24111;
    wire N__24108;
    wire N__24103;
    wire N__24098;
    wire N__24095;
    wire N__24094;
    wire N__24093;
    wire N__24090;
    wire N__24085;
    wire N__24082;
    wire N__24079;
    wire N__24076;
    wire N__24071;
    wire N__24062;
    wire N__24061;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24047;
    wire N__24044;
    wire N__24043;
    wire N__24042;
    wire N__24041;
    wire N__24040;
    wire N__24039;
    wire N__24038;
    wire N__24037;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24022;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24014;
    wire N__24011;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__23999;
    wire N__23994;
    wire N__23983;
    wire N__23972;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23956;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23936;
    wire N__23935;
    wire N__23932;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23848;
    wire N__23843;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23816;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23786;
    wire N__23783;
    wire N__23780;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23728;
    wire N__23723;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23677;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23656;
    wire N__23655;
    wire N__23654;
    wire N__23649;
    wire N__23644;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23593;
    wire N__23588;
    wire N__23587;
    wire N__23584;
    wire N__23581;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23563;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23545;
    wire N__23544;
    wire N__23543;
    wire N__23542;
    wire N__23541;
    wire N__23540;
    wire N__23539;
    wire N__23538;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23522;
    wire N__23521;
    wire N__23520;
    wire N__23519;
    wire N__23518;
    wire N__23515;
    wire N__23512;
    wire N__23511;
    wire N__23508;
    wire N__23505;
    wire N__23502;
    wire N__23499;
    wire N__23496;
    wire N__23491;
    wire N__23490;
    wire N__23489;
    wire N__23488;
    wire N__23487;
    wire N__23486;
    wire N__23485;
    wire N__23484;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23469;
    wire N__23466;
    wire N__23461;
    wire N__23456;
    wire N__23453;
    wire N__23442;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23424;
    wire N__23415;
    wire N__23410;
    wire N__23403;
    wire N__23396;
    wire N__23393;
    wire N__23392;
    wire N__23391;
    wire N__23388;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23359;
    wire N__23356;
    wire N__23353;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23341;
    wire N__23340;
    wire N__23339;
    wire N__23338;
    wire N__23335;
    wire N__23326;
    wire N__23323;
    wire N__23320;
    wire N__23315;
    wire N__23312;
    wire N__23311;
    wire N__23306;
    wire N__23303;
    wire N__23302;
    wire N__23301;
    wire N__23298;
    wire N__23297;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23274;
    wire N__23267;
    wire N__23264;
    wire N__23261;
    wire N__23258;
    wire N__23255;
    wire N__23254;
    wire N__23253;
    wire N__23252;
    wire N__23251;
    wire N__23248;
    wire N__23239;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23224;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23167;
    wire N__23164;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23095;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23050;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23020;
    wire N__23017;
    wire N__23012;
    wire N__23009;
    wire N__23008;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22955;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22942;
    wire N__22937;
    wire N__22934;
    wire N__22931;
    wire N__22930;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22915;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22877;
    wire N__22874;
    wire N__22871;
    wire N__22870;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22841;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22813;
    wire N__22812;
    wire N__22811;
    wire N__22808;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22790;
    wire N__22789;
    wire N__22786;
    wire N__22785;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22768;
    wire N__22763;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22744;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22724;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22666;
    wire N__22665;
    wire N__22660;
    wire N__22657;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22636;
    wire N__22633;
    wire N__22632;
    wire N__22627;
    wire N__22624;
    wire N__22619;
    wire N__22616;
    wire N__22615;
    wire N__22612;
    wire N__22611;
    wire N__22608;
    wire N__22601;
    wire N__22598;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22558;
    wire N__22553;
    wire N__22550;
    wire N__22549;
    wire N__22548;
    wire N__22547;
    wire N__22544;
    wire N__22543;
    wire N__22540;
    wire N__22539;
    wire N__22538;
    wire N__22537;
    wire N__22528;
    wire N__22525;
    wire N__22524;
    wire N__22523;
    wire N__22522;
    wire N__22521;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22504;
    wire N__22503;
    wire N__22500;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22486;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22453;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22396;
    wire N__22391;
    wire N__22388;
    wire N__22387;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22351;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22333;
    wire N__22332;
    wire N__22331;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22323;
    wire N__22322;
    wire N__22319;
    wire N__22312;
    wire N__22305;
    wire N__22302;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22264;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22252;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22237;
    wire N__22234;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22153;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22138;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22106;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22094;
    wire N__22091;
    wire N__22090;
    wire N__22089;
    wire N__22086;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22074;
    wire N__22071;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22037;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21928;
    wire N__21923;
    wire N__21920;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21908;
    wire N__21907;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21853;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21778;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21743;
    wire N__21740;
    wire N__21739;
    wire N__21736;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21719;
    wire N__21716;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21688;
    wire N__21685;
    wire N__21682;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21625;
    wire N__21622;
    wire N__21617;
    wire N__21616;
    wire N__21615;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21603;
    wire N__21596;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21569;
    wire N__21566;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21545;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21512;
    wire N__21509;
    wire N__21506;
    wire N__21503;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21425;
    wire N__21422;
    wire N__21419;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21331;
    wire N__21326;
    wire N__21323;
    wire N__21320;
    wire N__21317;
    wire N__21314;
    wire N__21311;
    wire N__21308;
    wire N__21305;
    wire N__21302;
    wire N__21299;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21280;
    wire N__21275;
    wire N__21272;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21241;
    wire N__21236;
    wire N__21233;
    wire N__21230;
    wire N__21229;
    wire N__21226;
    wire N__21221;
    wire N__21218;
    wire N__21217;
    wire N__21216;
    wire N__21215;
    wire N__21214;
    wire N__21213;
    wire N__21208;
    wire N__21199;
    wire N__21198;
    wire N__21197;
    wire N__21196;
    wire N__21195;
    wire N__21190;
    wire N__21183;
    wire N__21180;
    wire N__21173;
    wire N__21170;
    wire N__21169;
    wire N__21168;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21156;
    wire N__21153;
    wire N__21152;
    wire N__21151;
    wire N__21150;
    wire N__21149;
    wire N__21148;
    wire N__21145;
    wire N__21140;
    wire N__21129;
    wire N__21124;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21097;
    wire N__21094;
    wire N__21091;
    wire N__21088;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21062;
    wire N__21061;
    wire N__21058;
    wire N__21055;
    wire N__21050;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21035;
    wire N__21034;
    wire N__21031;
    wire N__21028;
    wire N__21023;
    wire N__21022;
    wire N__21019;
    wire N__21016;
    wire N__21011;
    wire N__21010;
    wire N__21007;
    wire N__21004;
    wire N__20999;
    wire N__20998;
    wire N__20995;
    wire N__20992;
    wire N__20989;
    wire N__20984;
    wire N__20983;
    wire N__20980;
    wire N__20977;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20959;
    wire N__20956;
    wire N__20955;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20945;
    wire N__20942;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20926;
    wire N__20921;
    wire N__20918;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20910;
    wire N__20907;
    wire N__20902;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20872;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20854;
    wire N__20851;
    wire N__20848;
    wire N__20845;
    wire N__20840;
    wire N__20839;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20815;
    wire N__20810;
    wire N__20809;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20794;
    wire N__20791;
    wire N__20788;
    wire N__20785;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20743;
    wire N__20742;
    wire N__20739;
    wire N__20738;
    wire N__20735;
    wire N__20730;
    wire N__20727;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20695;
    wire N__20692;
    wire N__20691;
    wire N__20688;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20653;
    wire N__20650;
    wire N__20649;
    wire N__20648;
    wire N__20647;
    wire N__20642;
    wire N__20639;
    wire N__20634;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20599;
    wire N__20596;
    wire N__20595;
    wire N__20592;
    wire N__20591;
    wire N__20588;
    wire N__20583;
    wire N__20580;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20554;
    wire N__20551;
    wire N__20550;
    wire N__20547;
    wire N__20540;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20516;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20461;
    wire N__20458;
    wire N__20457;
    wire N__20454;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20300;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20288;
    wire N__20285;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20259;
    wire N__20258;
    wire N__20257;
    wire N__20254;
    wire N__20247;
    wire N__20244;
    wire N__20237;
    wire N__20236;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20228;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20216;
    wire N__20213;
    wire N__20204;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20196;
    wire N__20193;
    wire N__20188;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20133;
    wire N__20132;
    wire N__20129;
    wire N__20124;
    wire N__20121;
    wire N__20114;
    wire N__20111;
    wire N__20110;
    wire N__20107;
    wire N__20106;
    wire N__20099;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20071;
    wire N__20068;
    wire N__20067;
    wire N__20064;
    wire N__20063;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20051;
    wire N__20048;
    wire N__20039;
    wire N__20038;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20020;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19917;
    wire N__19916;
    wire N__19913;
    wire N__19908;
    wire N__19905;
    wire N__19898;
    wire N__19895;
    wire N__19894;
    wire N__19891;
    wire N__19890;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19867;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19852;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19840;
    wire N__19839;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19810;
    wire N__19805;
    wire N__19802;
    wire N__19801;
    wire N__19800;
    wire N__19799;
    wire N__19798;
    wire N__19789;
    wire N__19786;
    wire N__19785;
    wire N__19784;
    wire N__19783;
    wire N__19782;
    wire N__19781;
    wire N__19780;
    wire N__19779;
    wire N__19778;
    wire N__19777;
    wire N__19776;
    wire N__19775;
    wire N__19774;
    wire N__19773;
    wire N__19772;
    wire N__19767;
    wire N__19766;
    wire N__19765;
    wire N__19764;
    wire N__19763;
    wire N__19754;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19738;
    wire N__19729;
    wire N__19726;
    wire N__19717;
    wire N__19714;
    wire N__19711;
    wire N__19706;
    wire N__19701;
    wire N__19694;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19672;
    wire N__19669;
    wire N__19666;
    wire N__19661;
    wire N__19658;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19592;
    wire N__19589;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19577;
    wire N__19574;
    wire N__19573;
    wire N__19570;
    wire N__19567;
    wire N__19564;
    wire N__19559;
    wire N__19556;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19523;
    wire N__19520;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19505;
    wire N__19502;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19466;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19454;
    wire N__19451;
    wire N__19450;
    wire N__19447;
    wire N__19444;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19414;
    wire N__19411;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19373;
    wire N__19370;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19358;
    wire N__19355;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19343;
    wire N__19340;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19325;
    wire N__19322;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19310;
    wire N__19307;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19297;
    wire N__19292;
    wire N__19289;
    wire N__19288;
    wire N__19285;
    wire N__19282;
    wire N__19277;
    wire N__19274;
    wire N__19273;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19259;
    wire N__19258;
    wire N__19255;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19243;
    wire N__19240;
    wire N__19235;
    wire N__19234;
    wire N__19231;
    wire N__19228;
    wire N__19225;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19213;
    wire N__19212;
    wire N__19211;
    wire N__19210;
    wire N__19209;
    wire N__19208;
    wire N__19207;
    wire N__19202;
    wire N__19199;
    wire N__19198;
    wire N__19197;
    wire N__19186;
    wire N__19183;
    wire N__19180;
    wire N__19175;
    wire N__19170;
    wire N__19163;
    wire N__19162;
    wire N__19161;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19150;
    wire N__19147;
    wire N__19146;
    wire N__19145;
    wire N__19144;
    wire N__19141;
    wire N__19140;
    wire N__19135;
    wire N__19132;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19106;
    wire N__19099;
    wire N__19096;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19075;
    wire N__19074;
    wire N__19071;
    wire N__19066;
    wire N__19061;
    wire N__19060;
    wire N__19059;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19047;
    wire N__19040;
    wire N__19039;
    wire N__19038;
    wire N__19035;
    wire N__19032;
    wire N__19029;
    wire N__19026;
    wire N__19023;
    wire N__19016;
    wire N__19015;
    wire N__19014;
    wire N__19011;
    wire N__19008;
    wire N__19003;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18985;
    wire N__18984;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18958;
    wire N__18957;
    wire N__18954;
    wire N__18949;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18934;
    wire N__18933;
    wire N__18930;
    wire N__18925;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18910;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18895;
    wire N__18890;
    wire N__18889;
    wire N__18886;
    wire N__18883;
    wire N__18878;
    wire N__18875;
    wire N__18874;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18864;
    wire N__18861;
    wire N__18854;
    wire N__18853;
    wire N__18850;
    wire N__18847;
    wire N__18842;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18830;
    wire N__18829;
    wire N__18826;
    wire N__18823;
    wire N__18818;
    wire N__18815;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18803;
    wire N__18802;
    wire N__18799;
    wire N__18796;
    wire N__18791;
    wire N__18790;
    wire N__18787;
    wire N__18784;
    wire N__18783;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18767;
    wire N__18766;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18719;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18707;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18692;
    wire N__18691;
    wire N__18688;
    wire N__18685;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18637;
    wire N__18636;
    wire N__18633;
    wire N__18632;
    wire N__18629;
    wire N__18624;
    wire N__18621;
    wire N__18614;
    wire N__18611;
    wire N__18610;
    wire N__18607;
    wire N__18606;
    wire N__18603;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18583;
    wire N__18580;
    wire N__18579;
    wire N__18576;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18508;
    wire N__18505;
    wire N__18504;
    wire N__18501;
    wire N__18500;
    wire N__18499;
    wire N__18496;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18427;
    wire N__18424;
    wire N__18423;
    wire N__18420;
    wire N__18413;
    wire N__18410;
    wire N__18409;
    wire N__18408;
    wire N__18405;
    wire N__18404;
    wire N__18401;
    wire N__18396;
    wire N__18393;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18373;
    wire N__18372;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18361;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18347;
    wire N__18344;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18310;
    wire N__18307;
    wire N__18306;
    wire N__18303;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18275;
    wire N__18272;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18262;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18249;
    wire N__18244;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18221;
    wire N__18218;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18206;
    wire N__18205;
    wire N__18204;
    wire N__18203;
    wire N__18202;
    wire N__18201;
    wire N__18200;
    wire N__18199;
    wire N__18198;
    wire N__18197;
    wire N__18196;
    wire N__18195;
    wire N__18194;
    wire N__18193;
    wire N__18186;
    wire N__18179;
    wire N__18170;
    wire N__18161;
    wire N__18160;
    wire N__18155;
    wire N__18150;
    wire N__18149;
    wire N__18146;
    wire N__18145;
    wire N__18142;
    wire N__18139;
    wire N__18132;
    wire N__18125;
    wire N__18122;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18049;
    wire N__18044;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18032;
    wire N__18029;
    wire N__18028;
    wire N__18025;
    wire N__18022;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18004;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17986;
    wire N__17983;
    wire N__17980;
    wire N__17975;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17965;
    wire N__17960;
    wire N__17957;
    wire N__17956;
    wire N__17953;
    wire N__17950;
    wire N__17947;
    wire N__17944;
    wire N__17939;
    wire N__17938;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17924;
    wire N__17923;
    wire N__17920;
    wire N__17917;
    wire N__17912;
    wire N__17911;
    wire N__17906;
    wire N__17903;
    wire N__17900;
    wire N__17899;
    wire N__17896;
    wire N__17893;
    wire N__17890;
    wire N__17885;
    wire N__17884;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17872;
    wire N__17869;
    wire N__17866;
    wire N__17861;
    wire N__17860;
    wire N__17855;
    wire N__17852;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17821;
    wire N__17820;
    wire N__17817;
    wire N__17816;
    wire N__17815;
    wire N__17810;
    wire N__17807;
    wire N__17802;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17788;
    wire N__17787;
    wire N__17784;
    wire N__17779;
    wire N__17776;
    wire N__17771;
    wire N__17768;
    wire N__17767;
    wire N__17764;
    wire N__17761;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17749;
    wire N__17746;
    wire N__17743;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17644;
    wire N__17641;
    wire N__17640;
    wire N__17637;
    wire N__17634;
    wire N__17631;
    wire N__17628;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17608;
    wire N__17607;
    wire N__17604;
    wire N__17603;
    wire N__17598;
    wire N__17595;
    wire N__17592;
    wire N__17589;
    wire N__17586;
    wire N__17583;
    wire N__17580;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17530;
    wire N__17527;
    wire N__17526;
    wire N__17523;
    wire N__17520;
    wire N__17517;
    wire N__17514;
    wire N__17507;
    wire N__17504;
    wire N__17501;
    wire N__17498;
    wire N__17497;
    wire N__17494;
    wire N__17493;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17465;
    wire N__17464;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17454;
    wire N__17451;
    wire N__17448;
    wire N__17445;
    wire N__17442;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17410;
    wire N__17407;
    wire N__17404;
    wire N__17403;
    wire N__17400;
    wire N__17397;
    wire N__17394;
    wire N__17389;
    wire N__17384;
    wire N__17381;
    wire N__17378;
    wire N__17375;
    wire N__17372;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17364;
    wire N__17361;
    wire N__17358;
    wire N__17355;
    wire N__17350;
    wire N__17345;
    wire N__17342;
    wire N__17339;
    wire N__17336;
    wire N__17333;
    wire N__17330;
    wire N__17329;
    wire N__17328;
    wire N__17325;
    wire N__17322;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17294;
    wire N__17293;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire N__17283;
    wire N__17280;
    wire N__17277;
    wire N__17274;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17254;
    wire N__17253;
    wire N__17252;
    wire N__17251;
    wire N__17248;
    wire N__17241;
    wire N__17238;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17218;
    wire N__17215;
    wire N__17214;
    wire N__17211;
    wire N__17208;
    wire N__17205;
    wire N__17202;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17186;
    wire N__17183;
    wire N__17180;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17169;
    wire N__17166;
    wire N__17163;
    wire N__17160;
    wire N__17157;
    wire N__17150;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17130;
    wire N__17127;
    wire N__17124;
    wire N__17121;
    wire N__17118;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17098;
    wire N__17095;
    wire N__17094;
    wire N__17091;
    wire N__17088;
    wire N__17085;
    wire N__17082;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17063;
    wire N__17060;
    wire N__17059;
    wire N__17058;
    wire N__17055;
    wire N__17052;
    wire N__17049;
    wire N__17046;
    wire N__17043;
    wire N__17040;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17020;
    wire N__17019;
    wire N__17016;
    wire N__17013;
    wire N__17010;
    wire N__17007;
    wire N__17004;
    wire N__17001;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16975;
    wire N__16974;
    wire N__16971;
    wire N__16968;
    wire N__16965;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16876;
    wire N__16873;
    wire N__16872;
    wire N__16869;
    wire N__16862;
    wire N__16859;
    wire N__16858;
    wire N__16855;
    wire N__16854;
    wire N__16851;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16789;
    wire N__16786;
    wire N__16783;
    wire N__16782;
    wire N__16781;
    wire N__16778;
    wire N__16773;
    wire N__16770;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16750;
    wire N__16747;
    wire N__16744;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16715;
    wire N__16712;
    wire N__16711;
    wire N__16706;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16684;
    wire N__16683;
    wire N__16682;
    wire N__16679;
    wire N__16674;
    wire N__16671;
    wire N__16670;
    wire N__16669;
    wire N__16668;
    wire N__16665;
    wire N__16662;
    wire N__16655;
    wire N__16652;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16570;
    wire N__16569;
    wire N__16568;
    wire N__16567;
    wire N__16566;
    wire N__16565;
    wire N__16564;
    wire N__16561;
    wire N__16556;
    wire N__16551;
    wire N__16544;
    wire N__16539;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16525;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16495;
    wire N__16494;
    wire N__16493;
    wire N__16492;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16473;
    wire N__16470;
    wire N__16469;
    wire N__16468;
    wire N__16467;
    wire N__16466;
    wire N__16465;
    wire N__16464;
    wire N__16463;
    wire N__16462;
    wire N__16461;
    wire N__16458;
    wire N__16455;
    wire N__16452;
    wire N__16449;
    wire N__16446;
    wire N__16415;
    wire N__16412;
    wire N__16409;
    wire N__16406;
    wire N__16403;
    wire N__16402;
    wire N__16401;
    wire N__16400;
    wire N__16397;
    wire N__16390;
    wire N__16385;
    wire N__16384;
    wire N__16381;
    wire N__16380;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16370;
    wire N__16369;
    wire N__16368;
    wire N__16367;
    wire N__16364;
    wire N__16361;
    wire N__16350;
    wire N__16347;
    wire N__16340;
    wire N__16337;
    wire N__16334;
    wire N__16331;
    wire N__16330;
    wire N__16329;
    wire N__16326;
    wire N__16321;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16307;
    wire N__16304;
    wire N__16301;
    wire N__16298;
    wire N__16297;
    wire N__16292;
    wire N__16289;
    wire N__16286;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16268;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16258;
    wire N__16255;
    wire N__16252;
    wire N__16249;
    wire N__16246;
    wire N__16243;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16226;
    wire N__16225;
    wire N__16222;
    wire N__16221;
    wire N__16218;
    wire N__16215;
    wire N__16212;
    wire N__16209;
    wire N__16206;
    wire N__16203;
    wire N__16200;
    wire N__16195;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16181;
    wire N__16178;
    wire N__16177;
    wire N__16174;
    wire N__16171;
    wire N__16168;
    wire N__16165;
    wire N__16162;
    wire N__16159;
    wire N__16156;
    wire N__16153;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16141;
    wire N__16138;
    wire N__16135;
    wire N__16132;
    wire N__16127;
    wire N__16124;
    wire N__16121;
    wire N__16118;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16108;
    wire N__16103;
    wire N__16102;
    wire N__16099;
    wire N__16096;
    wire N__16093;
    wire N__16088;
    wire N__16087;
    wire N__16084;
    wire N__16083;
    wire N__16080;
    wire N__16077;
    wire N__16074;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16049;
    wire N__16046;
    wire N__16045;
    wire N__16040;
    wire N__16037;
    wire N__16034;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16009;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15992;
    wire N__15989;
    wire N__15986;
    wire N__15983;
    wire N__15982;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15970;
    wire N__15969;
    wire N__15966;
    wire N__15963;
    wire N__15960;
    wire N__15953;
    wire N__15952;
    wire N__15951;
    wire N__15950;
    wire N__15949;
    wire N__15938;
    wire N__15935;
    wire N__15934;
    wire N__15933;
    wire N__15932;
    wire N__15927;
    wire N__15924;
    wire N__15921;
    wire N__15920;
    wire N__15917;
    wire N__15910;
    wire N__15905;
    wire N__15904;
    wire N__15901;
    wire N__15898;
    wire N__15893;
    wire N__15890;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15863;
    wire N__15862;
    wire N__15859;
    wire N__15856;
    wire N__15853;
    wire N__15850;
    wire N__15845;
    wire N__15842;
    wire N__15841;
    wire N__15840;
    wire N__15839;
    wire N__15836;
    wire N__15835;
    wire N__15828;
    wire N__15825;
    wire N__15822;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15806;
    wire N__15805;
    wire N__15802;
    wire N__15799;
    wire N__15798;
    wire N__15793;
    wire N__15790;
    wire N__15787;
    wire N__15782;
    wire N__15779;
    wire N__15778;
    wire N__15775;
    wire N__15772;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15754;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15736;
    wire N__15731;
    wire N__15728;
    wire N__15725;
    wire N__15722;
    wire N__15721;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15707;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15697;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15668;
    wire N__15665;
    wire N__15664;
    wire N__15659;
    wire N__15656;
    wire N__15653;
    wire N__15650;
    wire N__15649;
    wire N__15644;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15634;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15619;
    wire N__15614;
    wire N__15611;
    wire N__15608;
    wire N__15605;
    wire N__15602;
    wire N__15601;
    wire N__15596;
    wire N__15593;
    wire N__15590;
    wire N__15587;
    wire N__15584;
    wire N__15581;
    wire N__15578;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15553;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15538;
    wire N__15533;
    wire N__15530;
    wire N__15527;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15503;
    wire N__15500;
    wire N__15499;
    wire N__15498;
    wire N__15493;
    wire N__15490;
    wire N__15485;
    wire N__15484;
    wire N__15481;
    wire N__15476;
    wire N__15473;
    wire N__15472;
    wire N__15467;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15427;
    wire N__15424;
    wire N__15421;
    wire N__15418;
    wire N__15413;
    wire N__15410;
    wire N__15407;
    wire N__15406;
    wire N__15403;
    wire N__15400;
    wire N__15395;
    wire N__15392;
    wire N__15391;
    wire N__15390;
    wire N__15383;
    wire N__15380;
    wire N__15379;
    wire N__15376;
    wire N__15375;
    wire N__15374;
    wire N__15373;
    wire N__15370;
    wire N__15361;
    wire N__15356;
    wire N__15355;
    wire N__15354;
    wire N__15353;
    wire N__15352;
    wire N__15351;
    wire N__15350;
    wire N__15349;
    wire N__15340;
    wire N__15337;
    wire N__15336;
    wire N__15335;
    wire N__15334;
    wire N__15331;
    wire N__15330;
    wire N__15329;
    wire N__15328;
    wire N__15325;
    wire N__15324;
    wire N__15323;
    wire N__15320;
    wire N__15319;
    wire N__15316;
    wire N__15307;
    wire N__15304;
    wire N__15299;
    wire N__15296;
    wire N__15285;
    wire N__15280;
    wire N__15269;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15229;
    wire N__15228;
    wire N__15225;
    wire N__15220;
    wire N__15215;
    wire N__15214;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15199;
    wire N__15198;
    wire N__15191;
    wire N__15188;
    wire N__15187;
    wire N__15182;
    wire N__15179;
    wire N__15178;
    wire N__15175;
    wire N__15174;
    wire N__15171;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15155;
    wire N__15152;
    wire N__15151;
    wire N__15148;
    wire N__15145;
    wire N__15140;
    wire N__15139;
    wire N__15138;
    wire N__15137;
    wire N__15136;
    wire N__15133;
    wire N__15132;
    wire N__15131;
    wire N__15130;
    wire N__15127;
    wire N__15124;
    wire N__15119;
    wire N__15116;
    wire N__15113;
    wire N__15108;
    wire N__15103;
    wire N__15102;
    wire N__15101;
    wire N__15100;
    wire N__15099;
    wire N__15098;
    wire N__15095;
    wire N__15090;
    wire N__15089;
    wire N__15088;
    wire N__15085;
    wire N__15082;
    wire N__15073;
    wire N__15072;
    wire N__15071;
    wire N__15070;
    wire N__15069;
    wire N__15068;
    wire N__15067;
    wire N__15066;
    wire N__15065;
    wire N__15064;
    wire N__15061;
    wire N__15056;
    wire N__15055;
    wire N__15054;
    wire N__15053;
    wire N__15048;
    wire N__15041;
    wire N__15036;
    wire N__15033;
    wire N__15026;
    wire N__15019;
    wire N__15018;
    wire N__15017;
    wire N__15016;
    wire N__15013;
    wire N__15010;
    wire N__15003;
    wire N__14998;
    wire N__14989;
    wire N__14984;
    wire N__14981;
    wire N__14966;
    wire N__14965;
    wire N__14962;
    wire N__14961;
    wire N__14960;
    wire N__14959;
    wire N__14958;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14941;
    wire N__14940;
    wire N__14939;
    wire N__14938;
    wire N__14937;
    wire N__14936;
    wire N__14935;
    wire N__14934;
    wire N__14933;
    wire N__14932;
    wire N__14931;
    wire N__14930;
    wire N__14929;
    wire N__14928;
    wire N__14927;
    wire N__14926;
    wire N__14925;
    wire N__14924;
    wire N__14923;
    wire N__14918;
    wire N__14917;
    wire N__14916;
    wire N__14913;
    wire N__14908;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14885;
    wire N__14876;
    wire N__14871;
    wire N__14864;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14850;
    wire N__14849;
    wire N__14848;
    wire N__14847;
    wire N__14846;
    wire N__14845;
    wire N__14844;
    wire N__14841;
    wire N__14836;
    wire N__14833;
    wire N__14822;
    wire N__14811;
    wire N__14800;
    wire N__14795;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14758;
    wire N__14753;
    wire N__14750;
    wire N__14749;
    wire N__14748;
    wire N__14745;
    wire N__14742;
    wire N__14739;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14675;
    wire N__14674;
    wire N__14671;
    wire N__14670;
    wire N__14669;
    wire N__14668;
    wire N__14667;
    wire N__14664;
    wire N__14661;
    wire N__14658;
    wire N__14653;
    wire N__14650;
    wire N__14647;
    wire N__14640;
    wire N__14637;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14609;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14596;
    wire N__14593;
    wire N__14590;
    wire N__14585;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14573;
    wire N__14570;
    wire N__14567;
    wire N__14564;
    wire N__14561;
    wire N__14558;
    wire N__14555;
    wire N__14552;
    wire N__14549;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14530;
    wire N__14527;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14513;
    wire N__14510;
    wire N__14509;
    wire N__14508;
    wire N__14507;
    wire N__14504;
    wire N__14501;
    wire N__14498;
    wire N__14495;
    wire N__14490;
    wire N__14487;
    wire N__14482;
    wire N__14477;
    wire N__14474;
    wire N__14473;
    wire N__14470;
    wire N__14467;
    wire N__14462;
    wire N__14461;
    wire N__14458;
    wire N__14455;
    wire N__14452;
    wire N__14447;
    wire N__14444;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14432;
    wire N__14429;
    wire N__14428;
    wire N__14425;
    wire N__14422;
    wire N__14417;
    wire N__14414;
    wire N__14413;
    wire N__14410;
    wire N__14407;
    wire N__14402;
    wire N__14399;
    wire N__14396;
    wire N__14393;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14378;
    wire N__14375;
    wire N__14372;
    wire N__14371;
    wire N__14366;
    wire N__14363;
    wire N__14360;
    wire N__14359;
    wire N__14356;
    wire N__14353;
    wire N__14348;
    wire N__14347;
    wire N__14344;
    wire N__14341;
    wire N__14336;
    wire N__14333;
    wire N__14332;
    wire N__14329;
    wire N__14326;
    wire N__14321;
    wire N__14318;
    wire N__14315;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14305;
    wire N__14300;
    wire N__14297;
    wire N__14296;
    wire N__14293;
    wire N__14290;
    wire N__14285;
    wire N__14282;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14270;
    wire N__14267;
    wire N__14266;
    wire N__14263;
    wire N__14260;
    wire N__14255;
    wire N__14252;
    wire N__14251;
    wire N__14248;
    wire N__14245;
    wire N__14240;
    wire N__14237;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14222;
    wire N__14219;
    wire N__14218;
    wire N__14215;
    wire N__14212;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14200;
    wire N__14199;
    wire N__14198;
    wire N__14197;
    wire N__14196;
    wire N__14195;
    wire N__14194;
    wire N__14193;
    wire N__14192;
    wire N__14191;
    wire N__14190;
    wire N__14189;
    wire N__14188;
    wire N__14187;
    wire N__14186;
    wire N__14185;
    wire N__14184;
    wire N__14177;
    wire N__14168;
    wire N__14159;
    wire N__14150;
    wire N__14143;
    wire N__14140;
    wire N__14137;
    wire N__14134;
    wire N__14123;
    wire N__14120;
    wire N__14117;
    wire N__14114;
    wire N__14113;
    wire N__14110;
    wire N__14107;
    wire N__14102;
    wire N__14099;
    wire N__14096;
    wire N__14093;
    wire N__14090;
    wire N__14087;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14075;
    wire N__14072;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14060;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14048;
    wire N__14045;
    wire N__14044;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14030;
    wire N__14027;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14000;
    wire N__13997;
    wire N__13994;
    wire N__13991;
    wire N__13988;
    wire N__13985;
    wire N__13984;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13969;
    wire N__13964;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13937;
    wire N__13936;
    wire N__13931;
    wire N__13928;
    wire N__13925;
    wire N__13922;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13891;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13844;
    wire N__13843;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13826;
    wire N__13823;
    wire N__13820;
    wire N__13819;
    wire N__13816;
    wire N__13813;
    wire N__13810;
    wire N__13805;
    wire N__13804;
    wire N__13799;
    wire N__13796;
    wire N__13793;
    wire N__13792;
    wire N__13787;
    wire N__13784;
    wire N__13783;
    wire N__13780;
    wire N__13777;
    wire N__13772;
    wire N__13769;
    wire N__13766;
    wire N__13763;
    wire N__13760;
    wire N__13757;
    wire N__13754;
    wire N__13751;
    wire N__13750;
    wire N__13749;
    wire N__13744;
    wire N__13741;
    wire N__13738;
    wire N__13733;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13721;
    wire N__13718;
    wire N__13715;
    wire N__13714;
    wire N__13711;
    wire N__13706;
    wire N__13703;
    wire N__13702;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13688;
    wire N__13685;
    wire N__13684;
    wire N__13683;
    wire N__13680;
    wire N__13677;
    wire N__13674;
    wire N__13671;
    wire N__13664;
    wire N__13663;
    wire N__13660;
    wire N__13657;
    wire N__13654;
    wire N__13651;
    wire N__13646;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13633;
    wire N__13630;
    wire N__13627;
    wire N__13624;
    wire N__13621;
    wire N__13616;
    wire N__13615;
    wire N__13610;
    wire N__13607;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13595;
    wire N__13592;
    wire N__13589;
    wire N__13586;
    wire N__13583;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13573;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13555;
    wire N__13554;
    wire N__13553;
    wire N__13548;
    wire N__13545;
    wire N__13542;
    wire N__13535;
    wire N__13534;
    wire N__13531;
    wire N__13528;
    wire N__13523;
    wire N__13520;
    wire N__13517;
    wire N__13516;
    wire N__13513;
    wire N__13510;
    wire N__13505;
    wire N__13504;
    wire N__13499;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13477;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire VCCG0;
    wire \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_10_cascade_ ;
    wire \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_11 ;
    wire \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_0_cascade_ ;
    wire \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_12 ;
    wire \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_9 ;
    wire \PCH_PWRGD.count_rst_5_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_9_cascade_ ;
    wire \PCH_PWRGD.count_0_8 ;
    wire \PCH_PWRGD.count_rst_6_cascade_ ;
    wire \PCH_PWRGD.count_0_9 ;
    wire \PCH_PWRGD.countZ0Z_8_cascade_ ;
    wire \PCH_PWRGD.count_rst_5 ;
    wire \PCH_PWRGD.count_rst_11_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_4_cascade_ ;
    wire \PCH_PWRGD.count_0_3 ;
    wire \PCH_PWRGD.count_rst_10 ;
    wire \PCH_PWRGD.count_0_4 ;
    wire \PCH_PWRGD.count_rst_10_cascade_ ;
    wire bfn_1_5_0_;
    wire \PCH_PWRGD.un2_count_1_cry_1 ;
    wire \PCH_PWRGD.countZ0Z_3 ;
    wire \PCH_PWRGD.un2_count_1_cry_2_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_2 ;
    wire \PCH_PWRGD.un2_count_1_axb_4 ;
    wire \PCH_PWRGD.un2_count_1_cry_3_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_3 ;
    wire \PCH_PWRGD.un2_count_1_cry_4 ;
    wire \PCH_PWRGD.un2_count_1_cry_5 ;
    wire \PCH_PWRGD.un2_count_1_cry_6 ;
    wire \PCH_PWRGD.countZ0Z_8 ;
    wire \PCH_PWRGD.un2_count_1_cry_7_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_7 ;
    wire \PCH_PWRGD.un2_count_1_cry_8 ;
    wire \PCH_PWRGD.un2_count_1_axb_9 ;
    wire \PCH_PWRGD.un2_count_1_cry_8_THRU_CO ;
    wire bfn_1_6_0_;
    wire \PCH_PWRGD.un2_count_1_cry_9 ;
    wire \PCH_PWRGD.un2_count_1_cry_10 ;
    wire \PCH_PWRGD.un2_count_1_cry_11 ;
    wire \PCH_PWRGD.un2_count_1_cry_12 ;
    wire \PCH_PWRGD.un2_count_1_cry_13 ;
    wire \PCH_PWRGD.un2_count_1_cry_14 ;
    wire \PCH_PWRGD.un2_count_1_axb_2 ;
    wire \PCH_PWRGD.count_rst_12 ;
    wire \PCH_PWRGD.count_0_2 ;
    wire \PCH_PWRGD.count_0_14 ;
    wire \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7 ;
    wire \PCH_PWRGD.countZ0Z_14 ;
    wire \PCH_PWRGD.count_0_6 ;
    wire \PCH_PWRGD.curr_state_RNISDK72Z0Z_0_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0 ;
    wire \PCH_PWRGD.un2_count_1_axb_1_cascade_ ;
    wire \PCH_PWRGD.N_2284_i_cascade_ ;
    wire \PCH_PWRGD.N_655_cascade_ ;
    wire \PCH_PWRGD.count_0_sqmuxa_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_1 ;
    wire \PCH_PWRGD.count_0_1 ;
    wire \PCH_PWRGD.count_rst_13 ;
    wire vr_ready_vccin;
    wire \PCH_PWRGD.N_2284_i ;
    wire \POWERLED.count_0_2 ;
    wire G_12;
    wire \POWERLED.count_0_11 ;
    wire \POWERLED.count_0_3 ;
    wire \POWERLED.count_0_0 ;
    wire \POWERLED.count_1_0_cascade_ ;
    wire \POWERLED.countZ0Z_0_cascade_ ;
    wire \POWERLED.count_1_1_cascade_ ;
    wire \POWERLED.countZ0Z_1_cascade_ ;
    wire \POWERLED.count_0_1 ;
    wire \POWERLED.count_0_4 ;
    wire bfn_1_11_0_;
    wire \POWERLED.count_1_2 ;
    wire \POWERLED.un1_count_cry_1 ;
    wire \POWERLED.count_1_3 ;
    wire \POWERLED.un1_count_cry_2_cZ0 ;
    wire \POWERLED.count_1_4 ;
    wire \POWERLED.un1_count_cry_3_cZ0 ;
    wire \POWERLED.un1_count_cry_4_cZ0 ;
    wire \POWERLED.un1_count_cry_5 ;
    wire \POWERLED.un1_count_cry_6 ;
    wire \POWERLED.un1_count_cry_7 ;
    wire \POWERLED.un1_count_cry_8 ;
    wire bfn_1_12_0_;
    wire \POWERLED.un1_count_cry_9 ;
    wire \POWERLED.count_1_11 ;
    wire \POWERLED.un1_count_cry_10 ;
    wire \POWERLED.un1_count_cry_11 ;
    wire \POWERLED.un1_count_cry_12 ;
    wire \POWERLED.un1_count_cry_13 ;
    wire \POWERLED.un1_count_cry_14 ;
    wire \POWERLED.count_1_12 ;
    wire \POWERLED.count_0_12 ;
    wire \POWERLED.N_437_cascade_ ;
    wire \POWERLED.N_2305_i_cascade_ ;
    wire \POWERLED.N_660_cascade_ ;
    wire \POWERLED.count_0_sqmuxa_i ;
    wire \POWERLED.pwm_out_1_sqmuxa_0 ;
    wire \POWERLED.pwm_out_en_cascade_ ;
    wire \POWERLED.pwm_outZ0 ;
    wire pwrbtn_led;
    wire vpp_ok;
    wire vddq_en;
    wire \RSMRST_PWRGD.countZ0Z_0 ;
    wire bfn_2_1_0_;
    wire \RSMRST_PWRGD.countZ0Z_1 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_0 ;
    wire \RSMRST_PWRGD.countZ0Z_2 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_1 ;
    wire \RSMRST_PWRGD.countZ0Z_3 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_2 ;
    wire \RSMRST_PWRGD.countZ0Z_4 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_3 ;
    wire \RSMRST_PWRGD.countZ0Z_5 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_4 ;
    wire \RSMRST_PWRGD.countZ0Z_6 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_5 ;
    wire \RSMRST_PWRGD.countZ0Z_7 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_6 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_7 ;
    wire \RSMRST_PWRGD.countZ0Z_8 ;
    wire bfn_2_2_0_;
    wire \RSMRST_PWRGD.countZ0Z_9 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_8 ;
    wire \RSMRST_PWRGD.countZ0Z_10 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_9 ;
    wire \RSMRST_PWRGD.countZ0Z_11 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_10 ;
    wire \RSMRST_PWRGD.countZ0Z_12 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_11 ;
    wire \RSMRST_PWRGD.countZ0Z_13 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_12 ;
    wire \RSMRST_PWRGD.countZ0Z_14 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_13 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_2_3_0_;
    wire \RSMRST_PWRGD.countZ0Z_15 ;
    wire \PCH_PWRGD.count_0_12 ;
    wire \PCH_PWRGD.count_rst_2 ;
    wire \PCH_PWRGD.un2_count_1_cry_4_THRU_CO ;
    wire \PCH_PWRGD.count_0_5 ;
    wire \PCH_PWRGD.count_rst_9_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_10 ;
    wire \PCH_PWRGD.un2_count_1_cry_10_THRU_CO ;
    wire \PCH_PWRGD.N_386_cascade_ ;
    wire \PCH_PWRGD.count_0_11 ;
    wire \PCH_PWRGD.count_rst_3_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_11 ;
    wire \PCH_PWRGD.count_rst_7_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_7 ;
    wire \PCH_PWRGD.un2_count_1_cry_6_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_axb_7_cascade_ ;
    wire \PCH_PWRGD.count_rst_14_cascade_ ;
    wire \PCH_PWRGD.count_rst_7 ;
    wire \PCH_PWRGD.count_0_7 ;
    wire \PCH_PWRGD.countZ0Z_5 ;
    wire \PCH_PWRGD.count_1_i_a2_6_0 ;
    wire \PCH_PWRGD.count_1_i_a2_4_0 ;
    wire \PCH_PWRGD.count_1_i_a2_5_0_cascade_ ;
    wire \PCH_PWRGD.count_1_i_a2_3_0 ;
    wire \PCH_PWRGD.count_1_i_a2_12_0 ;
    wire \PCH_PWRGD.countZ0Z_0 ;
    wire \PCH_PWRGD.count_1_i_a2_12_0_cascade_ ;
    wire \PCH_PWRGD.count_0_0 ;
    wire \PCH_PWRGD.countZ0Z_15 ;
    wire \PCH_PWRGD.countZ0Z_15_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_13 ;
    wire \PCH_PWRGD.countZ0Z_6 ;
    wire \PCH_PWRGD.countZ0Z_12 ;
    wire \PCH_PWRGD.count_1_i_a2_1_0 ;
    wire \PCH_PWRGD.count_1_i_a2_0_0_cascade_ ;
    wire \PCH_PWRGD.count_1_i_a2_2_0 ;
    wire \PCH_PWRGD.count_1_i_a2_11_0 ;
    wire \PCH_PWRGD.count_rst ;
    wire \PCH_PWRGD.count_0_15 ;
    wire \PCH_PWRGD.count_rst_1 ;
    wire \PCH_PWRGD.count_0_13 ;
    wire \PCH_PWRGD.count_rst_4 ;
    wire \PCH_PWRGD.count_0_10 ;
    wire \PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ;
    wire \PCH_PWRGD.count_0_sqmuxa ;
    wire \PCH_PWRGD.N_2266_i_cascade_ ;
    wire \PCH_PWRGD.curr_state_0_1 ;
    wire \PCH_PWRGD.m6_i_i_a2_cascade_ ;
    wire \PCH_PWRGD.curr_state_7_0 ;
    wire \PCH_PWRGD.curr_stateZ0Z_0 ;
    wire \PCH_PWRGD.curr_stateZ0Z_0_cascade_ ;
    wire \PCH_PWRGD.N_655 ;
    wire \PCH_PWRGD.curr_stateZ0Z_1 ;
    wire \PCH_PWRGD.N_386 ;
    wire \PCH_PWRGD.curr_state_0_sqmuxa_cascade_ ;
    wire \PCH_PWRGD.curr_state_0_0 ;
    wire \VPP_VDDQ.N_53_cascade_ ;
    wire \VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ;
    wire \VPP_VDDQ.curr_state_2_0_1 ;
    wire \VPP_VDDQ.curr_state_2_0_0 ;
    wire \VPP_VDDQ.m4_0_0_cascade_ ;
    wire \VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.N_60_cascade_ ;
    wire \VPP_VDDQ.N_60_i ;
    wire \VPP_VDDQ.N_60 ;
    wire \VPP_VDDQ.delayed_vddq_okZ0 ;
    wire \VPP_VDDQ.delayed_vddq_ok_en ;
    wire VPP_VDDQ_delayed_vddq_ok_cascade_;
    wire vccst_pwrgd;
    wire \VPP_VDDQ.curr_state_2_RNIZ0Z_1_cascade_ ;
    wire pch_pwrok;
    wire \POWERLED.pwm_out_1_sqmuxa ;
    wire \POWERLED.un79_clk_100khzlt6 ;
    wire \POWERLED.un79_clk_100khzlto15_5_cascade_ ;
    wire \POWERLED.un79_clk_100khzlto15_4 ;
    wire \POWERLED.un79_clk_100khzlto15_7_cascade_ ;
    wire \POWERLED.un79_clk_100khz ;
    wire \POWERLED.un79_clk_100khz_cascade_ ;
    wire \POWERLED.g0_2_1 ;
    wire \POWERLED.un1_count_cry_14_c_RNIDQ1DZ0 ;
    wire \POWERLED.count_0_15 ;
    wire \POWERLED.count_1_7 ;
    wire \POWERLED.count_0_7 ;
    wire \POWERLED.count_1_8 ;
    wire \POWERLED.count_0_8 ;
    wire \POWERLED.count_1_9 ;
    wire \POWERLED.count_0_9 ;
    wire \POWERLED.count_1_13 ;
    wire \POWERLED.count_0_13 ;
    wire \POWERLED.count_1_5 ;
    wire \POWERLED.count_0_5 ;
    wire \POWERLED.count_1_14 ;
    wire \POWERLED.count_0_14 ;
    wire \POWERLED.count_1_6 ;
    wire \POWERLED.count_0_6 ;
    wire \POWERLED.count_1_10 ;
    wire \POWERLED.count_0_10 ;
    wire v33a_enn;
    wire \HDA_STRAP.N_16_cascade_ ;
    wire \PCH_PWRGD.delayed_vccin_okZ0_cascade_ ;
    wire N_428_cascade_;
    wire gpio_fpga_soc_1;
    wire \HDA_STRAP.m14_i_0_cascade_ ;
    wire N_428;
    wire \HDA_STRAP.curr_stateZ0Z_1 ;
    wire \HDA_STRAP.curr_stateZ0Z_0 ;
    wire \HDA_STRAP.curr_stateZ0Z_2 ;
    wire \HDA_STRAP.HDA_SDO_ATP_3_0 ;
    wire \HDA_STRAP.HDA_SDO_ATP_3_0_cascade_ ;
    wire hda_sdo_atp;
    wire \PCH_PWRGD.N_670 ;
    wire \PCH_PWRGD.N_2266_i ;
    wire \PCH_PWRGD.N_38_f0 ;
    wire \PCH_PWRGD.curr_state_0_sqmuxa ;
    wire \PCH_PWRGD.N_38_f0_cascade_ ;
    wire \PCH_PWRGD.delayed_vccin_ok_0 ;
    wire \VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_ ;
    wire \VPP_VDDQ.count_2_1_sqmuxa_cascade_ ;
    wire \VPP_VDDQ.count_2_1_0_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2_0_0 ;
    wire \VPP_VDDQ.count_2_1_1 ;
    wire \VPP_VDDQ.count_2Z0Z_1 ;
    wire \VPP_VDDQ.count_2_1_1_cascade_ ;
    wire slp_susn;
    wire v5a_ok;
    wire v33a_ok;
    wire v1p8a_ok;
    wire rsmrst_pwrgd_signal_cascade_;
    wire \RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_ ;
    wire \RSMRST_PWRGD.N_264_i ;
    wire \VPP_VDDQ.un9_clk_100khz_1 ;
    wire \VPP_VDDQ.un9_clk_100khz_13_cascade_ ;
    wire \VPP_VDDQ.N_1_i ;
    wire \VPP_VDDQ.curr_state_2Z0Z_1 ;
    wire \VPP_VDDQ.N_1_i_cascade_ ;
    wire \VPP_VDDQ.N_664 ;
    wire N_639;
    wire \VPP_VDDQ.curr_state_2Z0Z_0 ;
    wire \VPP_VDDQ.curr_state_2_RNIZ0Z_1 ;
    wire \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2_0_9 ;
    wire \VPP_VDDQ.count_2Z0Z_9_cascade_ ;
    wire \VPP_VDDQ.un9_clk_100khz_7 ;
    wire \VPP_VDDQ.count_2Z0Z_7 ;
    wire \VPP_VDDQ.count_2_0_11 ;
    wire \VPP_VDDQ.un9_clk_100khz_10 ;
    wire \VPP_VDDQ.count_2_0_12 ;
    wire \VPP_VDDQ.count_2_0_13 ;
    wire \VPP_VDDQ.count_2_0_14 ;
    wire \POWERLED.N_2305_i ;
    wire \POWERLED.N_660 ;
    wire \POWERLED.curr_state_1_0 ;
    wire N_557_g;
    wire bfn_4_10_0_;
    wire \POWERLED.mult1_un117_sum_i ;
    wire \POWERLED.mult1_un117_sum_i_0_8 ;
    wire \POWERLED.mult1_un124_sum_cry_2 ;
    wire \POWERLED.mult1_un124_sum_axb_4_l_fx ;
    wire \POWERLED.mult1_un124_sum_cry_3 ;
    wire \POWERLED.mult1_un124_sum_cry_4 ;
    wire \POWERLED.mult1_un124_sum_cry_5 ;
    wire \POWERLED.mult1_un124_sum_cry_6 ;
    wire \POWERLED.mult1_un124_sum_cry_7 ;
    wire \POWERLED.mult1_un124_sum_axb_7_l_fx ;
    wire bfn_4_11_0_;
    wire \POWERLED.mult1_un117_sum_cry_3_s ;
    wire \POWERLED.mult1_un117_sum_cry_2 ;
    wire \POWERLED.mult1_un117_sum_cry_4_s ;
    wire \POWERLED.mult1_un117_sum_cry_3 ;
    wire \POWERLED.mult1_un117_sum_cry_5_s ;
    wire \POWERLED.mult1_un117_sum_cry_4 ;
    wire \POWERLED.mult1_un117_sum_cry_6_s ;
    wire \POWERLED.mult1_un117_sum_cry_5 ;
    wire \POWERLED.mult1_un124_sum_axb_8 ;
    wire \POWERLED.mult1_un117_sum_cry_6 ;
    wire \POWERLED.mult1_un117_sum_cry_7 ;
    wire \POWERLED.mult1_un117_sum_s_8 ;
    wire \POWERLED.mult1_un110_sum_i_0_8 ;
    wire bfn_4_12_0_;
    wire \POWERLED.mult1_un110_sum_cry_3_s ;
    wire \POWERLED.mult1_un110_sum_cry_2 ;
    wire \POWERLED.mult1_un110_sum_cry_4_s ;
    wire \POWERLED.mult1_un110_sum_cry_3 ;
    wire \POWERLED.mult1_un110_sum_cry_5_s ;
    wire \POWERLED.mult1_un110_sum_cry_4 ;
    wire \POWERLED.mult1_un110_sum_cry_6_s ;
    wire \POWERLED.mult1_un110_sum_cry_5 ;
    wire \POWERLED.mult1_un117_sum_axb_8 ;
    wire \POWERLED.mult1_un110_sum_cry_6 ;
    wire \POWERLED.mult1_un110_sum_cry_7 ;
    wire \POWERLED.mult1_un110_sum_s_8 ;
    wire \POWERLED.mult1_un110_sum_s_8_cascade_ ;
    wire bfn_4_13_0_;
    wire \POWERLED.mult1_un103_sum_cry_3_s ;
    wire \POWERLED.mult1_un103_sum_cry_2 ;
    wire \POWERLED.mult1_un103_sum_cry_4_s ;
    wire \POWERLED.mult1_un103_sum_cry_3 ;
    wire \POWERLED.mult1_un103_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_cry_4 ;
    wire \POWERLED.mult1_un103_sum_cry_6_s ;
    wire \POWERLED.mult1_un103_sum_cry_5 ;
    wire \POWERLED.mult1_un110_sum_axb_8 ;
    wire \POWERLED.mult1_un103_sum_cry_6 ;
    wire \POWERLED.mult1_un103_sum_cry_7 ;
    wire \POWERLED.mult1_un103_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un103_sum_i_0_8 ;
    wire \POWERLED.countZ0Z_0 ;
    wire \POWERLED.un1_count_cry_0_i ;
    wire bfn_4_14_0_;
    wire \POWERLED.countZ0Z_1 ;
    wire \POWERLED.N_5036_i ;
    wire \POWERLED.un85_clk_100khz_cry_0 ;
    wire \POWERLED.countZ0Z_2 ;
    wire \POWERLED.N_5037_i ;
    wire \POWERLED.un85_clk_100khz_cry_1 ;
    wire \POWERLED.countZ0Z_3 ;
    wire \POWERLED.N_5038_i ;
    wire \POWERLED.un85_clk_100khz_cry_2 ;
    wire \POWERLED.countZ0Z_4 ;
    wire \POWERLED.N_5039_i ;
    wire \POWERLED.un85_clk_100khz_cry_3 ;
    wire \POWERLED.countZ0Z_5 ;
    wire \POWERLED.N_5040_i ;
    wire \POWERLED.un85_clk_100khz_cry_4 ;
    wire \POWERLED.countZ0Z_6 ;
    wire \POWERLED.N_5041_i ;
    wire \POWERLED.un85_clk_100khz_cry_5 ;
    wire \POWERLED.countZ0Z_7 ;
    wire \POWERLED.mult1_un117_sum_i_8 ;
    wire \POWERLED.N_5042_i ;
    wire \POWERLED.un85_clk_100khz_cry_6 ;
    wire \POWERLED.un85_clk_100khz_cry_7 ;
    wire \POWERLED.mult1_un110_sum_i_8 ;
    wire \POWERLED.countZ0Z_8 ;
    wire \POWERLED.N_5043_i ;
    wire bfn_4_15_0_;
    wire \POWERLED.countZ0Z_9 ;
    wire \POWERLED.N_5044_i ;
    wire \POWERLED.un85_clk_100khz_cry_8 ;
    wire \POWERLED.countZ0Z_10 ;
    wire \POWERLED.mult1_un96_sum_i_8 ;
    wire \POWERLED.N_5045_i ;
    wire \POWERLED.un85_clk_100khz_cry_9 ;
    wire \POWERLED.countZ0Z_11 ;
    wire \POWERLED.N_5046_i ;
    wire \POWERLED.un85_clk_100khz_cry_10 ;
    wire \POWERLED.countZ0Z_12 ;
    wire \POWERLED.N_5047_i ;
    wire \POWERLED.un85_clk_100khz_cry_11 ;
    wire \POWERLED.countZ0Z_13 ;
    wire \POWERLED.N_5048_i ;
    wire \POWERLED.un85_clk_100khz_cry_12 ;
    wire \POWERLED.countZ0Z_14 ;
    wire \POWERLED.N_5049_i ;
    wire \POWERLED.un85_clk_100khz_cry_13 ;
    wire \POWERLED.countZ0Z_15 ;
    wire \POWERLED.N_5050_i ;
    wire \POWERLED.un85_clk_100khz_cry_14 ;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0 ;
    wire bfn_4_16_0_;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ;
    wire \POWERLED.mult1_un89_sum_i_8 ;
    wire \POWERLED.mult1_un68_sum_i_8 ;
    wire bfn_5_1_0_;
    wire \HDA_STRAP.un1_count_1_cry_0 ;
    wire \HDA_STRAP.un1_count_1_cry_1 ;
    wire \HDA_STRAP.un1_count_1_cry_2 ;
    wire \HDA_STRAP.un1_count_1_cry_3 ;
    wire \HDA_STRAP.un1_count_1_cry_4 ;
    wire \HDA_STRAP.un1_count_1_cry_5_THRU_CO ;
    wire \HDA_STRAP.un1_count_1_cry_5 ;
    wire \HDA_STRAP.un1_count_1_cry_6 ;
    wire \HDA_STRAP.un1_count_1_cry_7 ;
    wire \HDA_STRAP.un1_count_1_cry_7_THRU_CO ;
    wire bfn_5_2_0_;
    wire \HDA_STRAP.un1_count_1_cry_8 ;
    wire \HDA_STRAP.un1_count_1_cry_9_THRU_CO ;
    wire \HDA_STRAP.un1_count_1_cry_9 ;
    wire \HDA_STRAP.un1_count_1_cry_10_THRU_CO ;
    wire \HDA_STRAP.un1_count_1_cry_10 ;
    wire \HDA_STRAP.un1_count_1_cry_11 ;
    wire \HDA_STRAP.un1_count_1_cry_12 ;
    wire \HDA_STRAP.un1_count_1_cry_13 ;
    wire \HDA_STRAP.un1_count_1_cry_14 ;
    wire \HDA_STRAP.un1_count_1_cry_15 ;
    wire bfn_5_3_0_;
    wire \HDA_STRAP.un1_count_1_cry_16 ;
    wire \RSMRST_PWRGD.N_92_1 ;
    wire \VPP_VDDQ.count_2_0_3 ;
    wire \VPP_VDDQ.count_2_0_5 ;
    wire \VPP_VDDQ.count_2_0_8 ;
    wire \VPP_VDDQ.count_2_0_10 ;
    wire \VPP_VDDQ.count_2Z0Z_0 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_1 ;
    wire bfn_5_8_0_;
    wire \VPP_VDDQ.un1_count_2_1_cry_1 ;
    wire \VPP_VDDQ.count_2_1_3 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_2 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_3 ;
    wire \VPP_VDDQ.count_2_1_5 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_4 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_5 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_7 ;
    wire \VPP_VDDQ.count_2_1_7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_6 ;
    wire \VPP_VDDQ.count_2_1_8 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_8 ;
    wire \VPP_VDDQ.count_2Z0Z_9 ;
    wire \VPP_VDDQ.count_2_1_9 ;
    wire bfn_5_9_0_;
    wire \VPP_VDDQ.count_2Z0Z_10 ;
    wire \VPP_VDDQ.count_2_1_10 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_9 ;
    wire \VPP_VDDQ.count_2Z0Z_11 ;
    wire \VPP_VDDQ.count_2_1_11 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_10 ;
    wire \VPP_VDDQ.count_2Z0Z_12 ;
    wire \VPP_VDDQ.count_2_1_12 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_11 ;
    wire \VPP_VDDQ.count_2Z0Z_13 ;
    wire \VPP_VDDQ.count_2_1_13 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_12 ;
    wire \VPP_VDDQ.count_2Z0Z_14 ;
    wire \VPP_VDDQ.count_2_1_14 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_13 ;
    wire \VPP_VDDQ.count_2Z0Z_15 ;
    wire \VPP_VDDQ.count_2_1_sqmuxa ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ;
    wire \VPP_VDDQ.count_2_0_15 ;
    wire bfn_5_10_0_;
    wire \POWERLED.mult1_un131_sum_cry_2 ;
    wire \POWERLED.mult1_un124_sum_cry_3_s ;
    wire \POWERLED.mult1_un131_sum_cry_3 ;
    wire \POWERLED.mult1_un124_sum_cry_4_s ;
    wire \POWERLED.mult1_un131_sum_cry_4 ;
    wire \POWERLED.mult1_un124_sum_cry_5_s ;
    wire \POWERLED.mult1_un131_sum_cry_5 ;
    wire \POWERLED.mult1_un124_sum_cry_6_s ;
    wire \POWERLED.mult1_un131_sum_cry_6 ;
    wire \POWERLED.mult1_un131_sum_axb_8 ;
    wire \POWERLED.mult1_un131_sum_cry_7 ;
    wire \POWERLED.mult1_un124_sum_i_0_8 ;
    wire bfn_5_11_0_;
    wire \POWERLED.mult1_un145_sum_cry_2_c ;
    wire \POWERLED.mult1_un145_sum_cry_3_c ;
    wire \POWERLED.mult1_un145_sum_cry_4_c ;
    wire \POWERLED.mult1_un145_sum_cry_5_c ;
    wire \POWERLED.mult1_un145_sum_cry_6_c ;
    wire \POWERLED.mult1_un145_sum_cry_7 ;
    wire \POWERLED.mult1_un145_sum_s_8_cascade_ ;
    wire bfn_5_12_0_;
    wire \POWERLED.mult1_un166_sum_cry_0 ;
    wire \POWERLED.mult1_un166_sum_cry_1 ;
    wire \POWERLED.mult1_un166_sum_cry_2 ;
    wire \POWERLED.mult1_un166_sum_cry_3 ;
    wire G_2150;
    wire \POWERLED.mult1_un166_sum_cry_4 ;
    wire \POWERLED.mult1_un166_sum_cry_5 ;
    wire \POWERLED.un85_clk_100khz_0 ;
    wire \POWERLED.un85_clk_100khz_2 ;
    wire \POWERLED.un85_clk_100khz_3 ;
    wire \POWERLED.mult1_un138_sum_i_8 ;
    wire \POWERLED.un85_clk_100khz_1 ;
    wire \POWERLED.mult1_un96_sum_i ;
    wire \POWERLED.mult1_un96_sum_i_0_8 ;
    wire \POWERLED.mult1_un103_sum_s_8 ;
    wire \POWERLED.mult1_un103_sum_i_8 ;
    wire \POWERLED.mult1_un124_sum_s_8 ;
    wire \POWERLED.mult1_un124_sum_i_8 ;
    wire bfn_5_14_0_;
    wire \POWERLED.mult1_un96_sum_cry_3_s ;
    wire \POWERLED.mult1_un96_sum_cry_2 ;
    wire \POWERLED.mult1_un96_sum_cry_4_s ;
    wire \POWERLED.mult1_un96_sum_cry_3 ;
    wire \POWERLED.mult1_un96_sum_cry_5_s ;
    wire \POWERLED.mult1_un96_sum_cry_4 ;
    wire \POWERLED.mult1_un96_sum_cry_6_s ;
    wire \POWERLED.mult1_un96_sum_cry_5 ;
    wire \POWERLED.mult1_un103_sum_axb_8 ;
    wire \POWERLED.mult1_un96_sum_cry_6 ;
    wire \POWERLED.mult1_un96_sum_cry_7 ;
    wire \POWERLED.mult1_un96_sum_s_8 ;
    wire \POWERLED.mult1_un131_sum_i_8 ;
    wire bfn_5_15_0_;
    wire \POWERLED.mult1_un89_sum_cry_3_s ;
    wire \POWERLED.mult1_un89_sum_cry_2 ;
    wire \POWERLED.mult1_un89_sum_cry_4_s ;
    wire \POWERLED.mult1_un89_sum_cry_3 ;
    wire \POWERLED.mult1_un89_sum_cry_5_s ;
    wire \POWERLED.mult1_un89_sum_cry_4 ;
    wire \POWERLED.mult1_un89_sum_cry_6_s ;
    wire \POWERLED.mult1_un89_sum_cry_5 ;
    wire \POWERLED.mult1_un96_sum_axb_8 ;
    wire \POWERLED.mult1_un89_sum_cry_6 ;
    wire \POWERLED.mult1_un89_sum_cry_7 ;
    wire \POWERLED.mult1_un89_sum_s_8 ;
    wire \POWERLED.mult1_un89_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un89_sum_i_0_8 ;
    wire \POWERLED.mult1_un75_sum_i_8 ;
    wire \POWERLED.mult1_un82_sum_i_0_8 ;
    wire \POWERLED.mult1_un89_sum_i ;
    wire \POWERLED.mult1_un82_sum_i_8 ;
    wire \HDA_STRAP.countZ0Z_8 ;
    wire \HDA_STRAP.countZ0Z_14 ;
    wire \HDA_STRAP.countZ0Z_6 ;
    wire \HDA_STRAP.countZ0Z_15 ;
    wire \HDA_STRAP.countZ0Z_4 ;
    wire \HDA_STRAP.countZ0Z_2 ;
    wire \HDA_STRAP.countZ0Z_3 ;
    wire \HDA_STRAP.countZ0Z_5 ;
    wire \HDA_STRAP.countZ0Z_11 ;
    wire \HDA_STRAP.countZ0Z_10 ;
    wire \HDA_STRAP.un4_count_12 ;
    wire \HDA_STRAP.un4_count_13_cascade_ ;
    wire \HDA_STRAP.un4_count_10 ;
    wire \HDA_STRAP.countZ0Z_9 ;
    wire \HDA_STRAP.countZ0Z_12 ;
    wire \HDA_STRAP.countZ0Z_13 ;
    wire \HDA_STRAP.countZ0Z_7 ;
    wire \HDA_STRAP.un4_count_11 ;
    wire \HDA_STRAP.countZ0Z_1 ;
    wire \HDA_STRAP.countZ0Z_0 ;
    wire \HDA_STRAP.countZ0Z_17 ;
    wire \HDA_STRAP.un4_count_9 ;
    wire \HDA_STRAP.un4_count ;
    wire \HDA_STRAP.curr_state_RNIH91AZ0Z_0 ;
    wire \HDA_STRAP.un1_count_1_cry_15_THRU_CO ;
    wire \HDA_STRAP.countZ0Z_16 ;
    wire \COUNTER.counterZ0Z_0 ;
    wire \COUNTER.counterZ0Z_1 ;
    wire bfn_6_4_0_;
    wire \COUNTER.counterZ0Z_2 ;
    wire \COUNTER.counter_1_cry_1_THRU_CO ;
    wire \COUNTER.counter_1_cry_1 ;
    wire \COUNTER.counterZ0Z_3 ;
    wire \COUNTER.counter_1_cry_2_THRU_CO ;
    wire \COUNTER.counter_1_cry_2 ;
    wire \COUNTER.counterZ0Z_4 ;
    wire \COUNTER.counter_1_cry_3_THRU_CO ;
    wire \COUNTER.counter_1_cry_3 ;
    wire \COUNTER.counterZ0Z_5 ;
    wire \COUNTER.counter_1_cry_4_THRU_CO ;
    wire \COUNTER.counter_1_cry_4 ;
    wire \COUNTER.counterZ0Z_6 ;
    wire \COUNTER.counter_1_cry_5_THRU_CO ;
    wire \COUNTER.counter_1_cry_5 ;
    wire \COUNTER.counterZ0Z_7 ;
    wire \COUNTER.counter_1_cry_6 ;
    wire \COUNTER.counterZ0Z_8 ;
    wire \COUNTER.counter_1_cry_7 ;
    wire \COUNTER.counter_1_cry_8 ;
    wire \COUNTER.counterZ0Z_9 ;
    wire bfn_6_5_0_;
    wire \COUNTER.counterZ0Z_10 ;
    wire \COUNTER.counter_1_cry_9 ;
    wire \COUNTER.counterZ0Z_11 ;
    wire \COUNTER.counter_1_cry_10 ;
    wire \COUNTER.counterZ0Z_12 ;
    wire \COUNTER.counter_1_cry_11 ;
    wire \COUNTER.counterZ0Z_13 ;
    wire \COUNTER.counter_1_cry_12 ;
    wire \COUNTER.counterZ0Z_14 ;
    wire \COUNTER.counter_1_cry_13 ;
    wire \COUNTER.counterZ0Z_15 ;
    wire \COUNTER.counter_1_cry_14 ;
    wire \COUNTER.counter_1_cry_15 ;
    wire \COUNTER.counter_1_cry_16 ;
    wire bfn_6_6_0_;
    wire \COUNTER.counter_1_cry_17 ;
    wire \COUNTER.counter_1_cry_18 ;
    wire \COUNTER.counter_1_cry_19 ;
    wire \COUNTER.counter_1_cry_20 ;
    wire \COUNTER.counter_1_cry_21 ;
    wire \COUNTER.counter_1_cry_22 ;
    wire \COUNTER.counterZ0Z_24 ;
    wire \COUNTER.counter_1_cry_23 ;
    wire \COUNTER.counter_1_cry_24 ;
    wire \COUNTER.counterZ0Z_25 ;
    wire bfn_6_7_0_;
    wire \COUNTER.counterZ0Z_26 ;
    wire \COUNTER.counter_1_cry_25 ;
    wire \COUNTER.counterZ0Z_27 ;
    wire \COUNTER.counter_1_cry_26 ;
    wire \COUNTER.counterZ0Z_28 ;
    wire \COUNTER.counter_1_cry_27 ;
    wire \COUNTER.counterZ0Z_29 ;
    wire \COUNTER.counter_1_cry_28 ;
    wire \COUNTER.counterZ0Z_30 ;
    wire \COUNTER.counter_1_cry_29 ;
    wire \COUNTER.counter_1_cry_30 ;
    wire \COUNTER.counterZ0Z_31 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_6 ;
    wire \VPP_VDDQ.count_2_0_4 ;
    wire \VPP_VDDQ.count_2_1_4 ;
    wire \VPP_VDDQ.count_2Z0Z_4 ;
    wire \VPP_VDDQ.count_2Z0Z_6 ;
    wire \VPP_VDDQ.count_2Z0Z_4_cascade_ ;
    wire \VPP_VDDQ.count_2_1_6 ;
    wire \VPP_VDDQ.un9_clk_100khz_0 ;
    wire \VPP_VDDQ.count_2_0_2 ;
    wire \VPP_VDDQ.count_2_1_2 ;
    wire \VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0 ;
    wire \VPP_VDDQ.count_2Z0Z_2 ;
    wire \VPP_VDDQ.count_2Z0Z_5 ;
    wire \VPP_VDDQ.count_2Z0Z_8 ;
    wire \VPP_VDDQ.count_2Z0Z_2_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_3 ;
    wire \VPP_VDDQ.un9_clk_100khz_9 ;
    wire bfn_6_10_0_;
    wire \POWERLED.mult1_un138_sum_cry_3_s ;
    wire \POWERLED.mult1_un138_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_cry_3_s ;
    wire \POWERLED.mult1_un138_sum_cry_4_s ;
    wire \POWERLED.mult1_un138_sum_cry_3 ;
    wire \POWERLED.mult1_un131_sum_cry_4_s ;
    wire \POWERLED.mult1_un138_sum_cry_5_s ;
    wire \POWERLED.mult1_un138_sum_cry_4 ;
    wire \POWERLED.mult1_un131_sum_cry_5_s ;
    wire \POWERLED.mult1_un138_sum_cry_6_s ;
    wire \POWERLED.mult1_un138_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_cry_6_s ;
    wire \POWERLED.mult1_un145_sum_axb_8 ;
    wire \POWERLED.mult1_un138_sum_cry_6 ;
    wire \POWERLED.mult1_un138_sum_axb_8 ;
    wire \POWERLED.mult1_un138_sum_cry_7 ;
    wire \POWERLED.mult1_un138_sum_s_8 ;
    wire \POWERLED.mult1_un138_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un138_sum_i_0_8 ;
    wire bfn_6_11_0_;
    wire \POWERLED.mult1_un152_sum_cry_2 ;
    wire \POWERLED.mult1_un145_sum_cry_3_s ;
    wire \POWERLED.mult1_un152_sum_cry_3 ;
    wire \POWERLED.mult1_un145_sum_cry_4_s ;
    wire \POWERLED.mult1_un152_sum_cry_4 ;
    wire \POWERLED.mult1_un145_sum_cry_5_s ;
    wire \POWERLED.mult1_un145_sum_s_8 ;
    wire \POWERLED.mult1_un152_sum_cry_5 ;
    wire \POWERLED.mult1_un145_sum_i_0_8 ;
    wire \POWERLED.mult1_un145_sum_cry_6_s ;
    wire \POWERLED.mult1_un152_sum_cry_6 ;
    wire \POWERLED.mult1_un152_sum_axb_8 ;
    wire \POWERLED.mult1_un152_sum_cry_7 ;
    wire \POWERLED.mult1_un131_sum_s_8 ;
    wire \POWERLED.mult1_un131_sum_i_0_8 ;
    wire bfn_6_12_0_;
    wire \POWERLED.mult1_un159_sum_cry_2_s ;
    wire \POWERLED.mult1_un159_sum_cry_1 ;
    wire \POWERLED.mult1_un152_sum_cry_3_s ;
    wire \POWERLED.mult1_un159_sum_cry_3_s ;
    wire \POWERLED.mult1_un159_sum_cry_2 ;
    wire \POWERLED.mult1_un152_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_cry_3 ;
    wire \POWERLED.mult1_un152_sum_cry_5_s ;
    wire \POWERLED.mult1_un159_sum_cry_5_s ;
    wire \POWERLED.mult1_un159_sum_cry_4 ;
    wire \POWERLED.mult1_un152_sum_cry_6_s ;
    wire \POWERLED.mult1_un166_sum_axb_6 ;
    wire \POWERLED.mult1_un159_sum_cry_5 ;
    wire \POWERLED.mult1_un159_sum_axb_7 ;
    wire \POWERLED.mult1_un159_sum_cry_6 ;
    wire \POWERLED.mult1_un159_sum_s_7 ;
    wire \POWERLED.mult1_un152_sum_s_8 ;
    wire \POWERLED.mult1_un152_sum_i_0_8 ;
    wire \POWERLED.mult1_un138_sum_i ;
    wire \POWERLED.mult1_un131_sum_i ;
    wire \POWERLED.mult1_un145_sum_i ;
    wire \POWERLED.mult1_un103_sum_i ;
    wire \POWERLED.mult1_un124_sum_i ;
    wire \POWERLED.mult1_un110_sum_i ;
    wire \POWERLED.mult1_un61_sum_i_8 ;
    wire bfn_6_14_0_;
    wire \POWERLED.mult1_un68_sum_cry_2 ;
    wire \POWERLED.mult1_un68_sum_cry_3 ;
    wire \POWERLED.mult1_un68_sum_cry_4 ;
    wire \POWERLED.mult1_un68_sum_cry_5 ;
    wire \POWERLED.mult1_un61_sum_i_0_8 ;
    wire \POWERLED.mult1_un68_sum_cry_6 ;
    wire \POWERLED.mult1_un68_sum_cry_7 ;
    wire \POWERLED.mult1_un68_sum_s_8_cascade_ ;
    wire bfn_6_15_0_;
    wire \POWERLED.mult1_un75_sum_cry_2 ;
    wire \POWERLED.mult1_un68_sum_cry_3_s ;
    wire \POWERLED.mult1_un75_sum_cry_3 ;
    wire \POWERLED.mult1_un68_sum_cry_4_s ;
    wire \POWERLED.mult1_un75_sum_cry_4 ;
    wire \POWERLED.mult1_un68_sum_s_8 ;
    wire \POWERLED.mult1_un68_sum_cry_5_s ;
    wire \POWERLED.mult1_un75_sum_cry_5 ;
    wire \POWERLED.mult1_un68_sum_cry_6_s ;
    wire \POWERLED.mult1_un68_sum_i_0_8 ;
    wire \POWERLED.mult1_un75_sum_cry_6 ;
    wire \POWERLED.mult1_un75_sum_axb_8 ;
    wire \POWERLED.mult1_un75_sum_cry_7 ;
    wire \POWERLED.mult1_un75_sum_s_8_cascade_ ;
    wire bfn_6_16_0_;
    wire \POWERLED.mult1_un82_sum_cry_3_s ;
    wire \POWERLED.mult1_un82_sum_cry_2 ;
    wire \POWERLED.mult1_un75_sum_cry_3_s ;
    wire \POWERLED.mult1_un82_sum_cry_4_s ;
    wire \POWERLED.mult1_un82_sum_cry_3 ;
    wire \POWERLED.mult1_un75_sum_cry_4_s ;
    wire \POWERLED.mult1_un82_sum_cry_5_s ;
    wire \POWERLED.mult1_un82_sum_cry_4 ;
    wire \POWERLED.mult1_un75_sum_s_8 ;
    wire \POWERLED.mult1_un75_sum_cry_5_s ;
    wire \POWERLED.mult1_un82_sum_cry_6_s ;
    wire \POWERLED.mult1_un82_sum_cry_5 ;
    wire \POWERLED.mult1_un75_sum_cry_6_s ;
    wire \POWERLED.mult1_un75_sum_i_0_8 ;
    wire \POWERLED.mult1_un89_sum_axb_8 ;
    wire \POWERLED.mult1_un82_sum_cry_6 ;
    wire \POWERLED.mult1_un82_sum_axb_8 ;
    wire \POWERLED.mult1_un82_sum_cry_7 ;
    wire \POWERLED.mult1_un82_sum_s_8 ;
    wire \POWERLED.mult1_un75_sum_i ;
    wire \POWERLED.count_off_0_9 ;
    wire \POWERLED.count_offZ0Z_9_cascade_ ;
    wire \POWERLED.count_off_0_10 ;
    wire \POWERLED.count_off_0_11 ;
    wire bfn_7_3_0_;
    wire \POWERLED.un3_count_off_1_cry_1_cZ0 ;
    wire \POWERLED.un3_count_off_1_cry_2 ;
    wire \POWERLED.un3_count_off_1_cry_3 ;
    wire \POWERLED.un3_count_off_1_cry_4 ;
    wire \POWERLED.un3_count_off_1_cry_5 ;
    wire \POWERLED.un3_count_off_1_cry_6 ;
    wire \POWERLED.un3_count_off_1_cry_7 ;
    wire \POWERLED.un3_count_off_1_cry_8 ;
    wire \POWERLED.count_offZ0Z_9 ;
    wire \POWERLED.count_off_1_9 ;
    wire bfn_7_4_0_;
    wire \POWERLED.count_offZ0Z_10 ;
    wire \POWERLED.count_off_1_10 ;
    wire \POWERLED.un3_count_off_1_cry_9 ;
    wire \POWERLED.count_offZ0Z_11 ;
    wire \POWERLED.count_off_1_11 ;
    wire \POWERLED.un3_count_off_1_cry_10 ;
    wire \POWERLED.count_offZ0Z_12 ;
    wire \POWERLED.un3_count_off_1_cry_11 ;
    wire \POWERLED.un3_count_off_1_cry_12 ;
    wire \POWERLED.un3_count_off_1_cry_13 ;
    wire \POWERLED.un3_count_off_1_cry_14 ;
    wire \POWERLED.count_off_1_12 ;
    wire \POWERLED.count_off_0_12 ;
    wire \COUNTER.counterZ0Z_19 ;
    wire \COUNTER.counterZ0Z_17 ;
    wire \COUNTER.counterZ0Z_18 ;
    wire \COUNTER.counterZ0Z_16 ;
    wire \COUNTER.counterZ0Z_23 ;
    wire \COUNTER.counterZ0Z_20 ;
    wire \COUNTER.counterZ0Z_21 ;
    wire \COUNTER.counterZ0Z_22 ;
    wire N_555;
    wire G_14;
    wire N_662;
    wire RSMRST_PWRGD_curr_state_0;
    wire \RSMRST_PWRGD.curr_stateZ0Z_1 ;
    wire VCCST_EN_i_1_cascade_;
    wire \POWERLED.un1_func_state25_6_0_o_N_5_cascade_ ;
    wire \POWERLED.N_432 ;
    wire \POWERLED.un1_func_state25_6_0_o_N_7_2 ;
    wire \POWERLED.func_state_1_ss0_i_0_0_1_1_cascade_ ;
    wire \POWERLED.N_423 ;
    wire \POWERLED.N_671 ;
    wire \POWERLED.func_state_enZ0 ;
    wire \POWERLED.func_stateZ0Z_1 ;
    wire \POWERLED.N_512_cascade_ ;
    wire \POWERLED.un1_clk_100khz_39_and_i_1_cascade_ ;
    wire \POWERLED.N_514 ;
    wire \POWERLED.N_508 ;
    wire \POWERLED.un1_clk_100khz_33_and_i_1_cascade_ ;
    wire \POWERLED.count_off_1_7 ;
    wire \POWERLED.count_off_0_7 ;
    wire \POWERLED.count_off_1_8 ;
    wire \POWERLED.count_off_0_8 ;
    wire bfn_7_11_0_;
    wire \POWERLED.mult1_un54_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6 ;
    wire \POWERLED.mult1_un54_sum_cry_7 ;
    wire \POWERLED.mult1_un47_sum_l_fx_6 ;
    wire bfn_7_12_0_;
    wire \POWERLED.mult1_un54_sum_i ;
    wire \POWERLED.mult1_un61_sum_cry_3_s ;
    wire \POWERLED.mult1_un61_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3_s ;
    wire \POWERLED.mult1_un61_sum_cry_4_s ;
    wire \POWERLED.mult1_un61_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4_s ;
    wire \POWERLED.mult1_un61_sum_cry_5_s ;
    wire \POWERLED.mult1_un61_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_cry_5_s ;
    wire \POWERLED.mult1_un61_sum_cry_6_s ;
    wire \POWERLED.mult1_un61_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6_s ;
    wire \POWERLED.mult1_un68_sum_axb_8 ;
    wire \POWERLED.mult1_un61_sum_cry_6 ;
    wire \POWERLED.mult1_un61_sum_axb_8 ;
    wire \POWERLED.mult1_un61_sum_cry_7 ;
    wire \POWERLED.mult1_un61_sum_s_8 ;
    wire \POWERLED.un1_dutycycle_53_i_28 ;
    wire \POWERLED.un1_dutycycle_53_axb_0 ;
    wire bfn_7_13_0_;
    wire \POWERLED.mult1_un138_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_0 ;
    wire \POWERLED.mult1_un131_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_1 ;
    wire \POWERLED.mult1_un124_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_2 ;
    wire \POWERLED.mult1_un117_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_3 ;
    wire \POWERLED.mult1_un110_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_4 ;
    wire \POWERLED.mult1_un103_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_5 ;
    wire \POWERLED.mult1_un96_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_6 ;
    wire \POWERLED.un1_dutycycle_53_cry_7 ;
    wire \POWERLED.mult1_un89_sum ;
    wire bfn_7_14_0_;
    wire \POWERLED.un1_dutycycle_53_cry_8 ;
    wire \POWERLED.mult1_un75_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_9 ;
    wire \POWERLED.un1_dutycycle_53_cry_10 ;
    wire \POWERLED.un1_dutycycle_53_cry_11 ;
    wire \POWERLED.mult1_un54_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_12 ;
    wire \POWERLED.un1_dutycycle_53_cry_13 ;
    wire \POWERLED.un1_dutycycle_53_cry_14 ;
    wire \POWERLED.un1_dutycycle_53_cry_15 ;
    wire bfn_7_15_0_;
    wire \POWERLED.CO2 ;
    wire \POWERLED.CO2_THRU_CO ;
    wire \POWERLED.dutycycle_RNIZ0Z_14 ;
    wire \POWERLED.mult1_un68_sum ;
    wire \POWERLED.mult1_un68_sum_i ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_15 ;
    wire \POWERLED.mult1_un82_sum ;
    wire \POWERLED.mult1_un82_sum_i ;
    wire \POWERLED.mult1_un61_sum ;
    wire \POWERLED.mult1_un61_sum_i ;
    wire \POWERLED.N_598_cascade_ ;
    wire \POWERLED.N_450_cascade_ ;
    wire \POWERLED.N_599 ;
    wire \POWERLED.N_449_cascade_ ;
    wire \POWERLED.N_2376_i ;
    wire \POWERLED.N_2376_i_cascade_ ;
    wire \POWERLED.count_offZ0Z_0_cascade_ ;
    wire \POWERLED.count_off_0_5 ;
    wire \POWERLED.count_off_1_5 ;
    wire \POWERLED.count_offZ0Z_5 ;
    wire \POWERLED.count_offZ0Z_5_cascade_ ;
    wire \POWERLED.count_off_0_0 ;
    wire \POWERLED.count_off_1_0 ;
    wire \POWERLED.count_off_0_2 ;
    wire \POWERLED.count_off_1_2 ;
    wire \POWERLED.count_offZ0Z_2 ;
    wire \POWERLED.count_off_1_13 ;
    wire \POWERLED.count_off_0_13 ;
    wire \POWERLED.count_off_1_14 ;
    wire \POWERLED.count_off_0_14 ;
    wire \POWERLED.un3_count_off_1_cry_14_c_RNIPGZ0Z497 ;
    wire \POWERLED.count_off_0_15 ;
    wire \POWERLED.count_offZ0Z_15 ;
    wire \POWERLED.count_offZ0Z_13 ;
    wire \POWERLED.count_offZ0Z_14 ;
    wire \POWERLED.count_offZ0Z_15_cascade_ ;
    wire \POWERLED.count_offZ0Z_0 ;
    wire \POWERLED.count_off_0_6 ;
    wire \POWERLED.count_off_1_6 ;
    wire \POWERLED.count_offZ0Z_6 ;
    wire \COUNTER.un4_counter_0_and ;
    wire bfn_8_4_0_;
    wire \COUNTER.un4_counter_1_and ;
    wire \COUNTER.un4_counter_0 ;
    wire \COUNTER.un4_counter_2_and ;
    wire \COUNTER.un4_counter_1 ;
    wire \COUNTER.un4_counter_3_and ;
    wire \COUNTER.un4_counter_2 ;
    wire \COUNTER.un4_counter_4_and ;
    wire \COUNTER.un4_counter_3 ;
    wire \COUNTER.un4_counter_5_and ;
    wire \COUNTER.un4_counter_4 ;
    wire \COUNTER.un4_counter_6_and ;
    wire \COUNTER.un4_counter_5 ;
    wire \COUNTER.un4_counter_7_and ;
    wire \COUNTER.un4_counter_6 ;
    wire COUNTER_un4_counter_7;
    wire bfn_8_5_0_;
    wire \POWERLED.N_673_0_cascade_ ;
    wire \POWERLED.N_423_0 ;
    wire v5s_enn_cascade_;
    wire \POWERLED.func_state_en_0_0 ;
    wire \POWERLED.func_stateZ1Z_0 ;
    wire \POWERLED.func_state_en_0_0_cascade_ ;
    wire RSMRSTn_fast;
    wire \POWERLED.un1_func_state25_6_0_0_0_2 ;
    wire \POWERLED.func_state_RNI5SKJ1Z0Z_1 ;
    wire vddq_ok;
    wire func_state_RNI_2_0_cascade_;
    wire \POWERLED.func_state_1_m0_1_1 ;
    wire \POWERLED.N_540_1 ;
    wire \POWERLED.N_542 ;
    wire \POWERLED.N_673 ;
    wire \POWERLED.func_state_1_m2s2_i_0_1_cascade_ ;
    wire \POWERLED.N_6_1 ;
    wire \POWERLED.N_74_cascade_ ;
    wire \POWERLED.func_state_1_m2_ns_1_1 ;
    wire \POWERLED.func_state_1_m2_1 ;
    wire \POWERLED.func_state_RNIBVNSZ0Z_0 ;
    wire \POWERLED.N_6_2 ;
    wire \POWERLED.dutycycle_1_0_iv_i_0_a2_0_1_2 ;
    wire \POWERLED.dutycycle_1_0_iv_i_0_0_2_cascade_ ;
    wire \POWERLED.N_71_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_0_cascade_ ;
    wire \POWERLED.mult1_un152_sum_i ;
    wire \POWERLED.N_426_i_cascade_ ;
    wire \POWERLED.dutycycle_eena_1 ;
    wire \POWERLED.N_71 ;
    wire \POWERLED.dutycycle_eena_1_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_2 ;
    wire COUNTER_un4_counter_7_THRU_CO;
    wire \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1GZ0 ;
    wire \POWERLED.dutycycleZ1Z_7 ;
    wire \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1GZ0_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434 ;
    wire bfn_8_11_0_;
    wire \POWERLED.un1_dutycycle_53_i_29 ;
    wire \POWERLED.mult1_un47_sum_cry_2 ;
    wire \POWERLED.mult1_un47_sum_cry_4_s ;
    wire \POWERLED.mult1_un47_sum_cry_3 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_4 ;
    wire \POWERLED.mult1_un47_sum_cry_5_s ;
    wire \POWERLED.mult1_un47_sum_cry_4 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_5 ;
    wire \POWERLED.mult1_un47_sum_cry_6_s ;
    wire \POWERLED.mult1_un47_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_7_THRU_CO ;
    wire \POWERLED.mult1_un47_sum_cry_6 ;
    wire \POWERLED.mult1_un54_sum_s_8 ;
    wire \POWERLED.mult1_un54_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un54_sum_i_8 ;
    wire \POWERLED.mult1_un47_sum_cry_3_s ;
    wire \POWERLED.mult1_un47_sum_l_fx_3 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_0 ;
    wire \POWERLED.dutycycle_RNIZ0Z_3_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_8 ;
    wire \POWERLED.dutycycle_RNIZ0Z_2 ;
    wire \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ;
    wire \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ;
    wire \POWERLED.mult1_un47_sum_axb_4 ;
    wire \POWERLED.mult1_un159_sum_i ;
    wire \POWERLED.dutycycle_en_10 ;
    wire \POWERLED.dutycycleZ0Z_13 ;
    wire \POWERLED.un1_dutycycle_53_41_0 ;
    wire \POWERLED.un1_dutycycle_53_40_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_13 ;
    wire \POWERLED.dutycycleZ1Z_9 ;
    wire \POWERLED.dutycycleZ0Z_4_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_8_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_6_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_7 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_8 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_5 ;
    wire \POWERLED.un1_dutycycle_53_31_a4_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_31_a5_1 ;
    wire \POWERLED.un1_dutycycle_53_31_a0_2 ;
    wire \POWERLED.dutycycle_RNIZ0Z_12 ;
    wire \POWERLED.dutycycleZ1Z_14 ;
    wire \POWERLED.dutycycle_RNI_12Z0Z_8_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_15 ;
    wire \POWERLED.dutycycleZ0Z_15 ;
    wire \POWERLED.dutycycleZ0Z_14_cascade_ ;
    wire \POWERLED.N_2381_i_cascade_ ;
    wire \POWERLED.un2_count_clk_17_0_0_a2_0_5 ;
    wire \POWERLED.dutycycle_RNIZ0Z_13 ;
    wire \POWERLED.dutycycleZ1Z_11 ;
    wire \POWERLED.dutycycle_en_7 ;
    wire \POWERLED.dutycycleZ0Z_9_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_11_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_2_1 ;
    wire \POWERLED.un1_dutycycle_53_2_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_13 ;
    wire \VPP_VDDQ.un6_count_8_cascade_ ;
    wire \VPP_VDDQ.un6_count_10 ;
    wire \VPP_VDDQ.un6_count_11 ;
    wire \VPP_VDDQ.un6_count_9 ;
    wire \POWERLED.G_30Z0Z_0_cascade_ ;
    wire VPP_VDDQ_un6_count;
    wire G_30_cascade_;
    wire N_626;
    wire VPP_VDDQ_curr_state_1;
    wire VPP_VDDQ_curr_state_0;
    wire \POWERLED.count_off_0_3 ;
    wire \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ;
    wire \POWERLED.count_offZ0Z_3 ;
    wire \POWERLED.count_offZ0Z_7 ;
    wire \POWERLED.count_offZ0Z_3_cascade_ ;
    wire \POWERLED.count_offZ0Z_8 ;
    wire \POWERLED.un34_clk_100khz_10 ;
    wire \POWERLED.un34_clk_100khz_11 ;
    wire \POWERLED.un34_clk_100khz_8_cascade_ ;
    wire \POWERLED.un34_clk_100khz_9 ;
    wire \POWERLED.count_offZ0Z_4 ;
    wire \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ;
    wire \POWERLED.count_off_0_4 ;
    wire \POWERLED.count_off_RNIZ0Z_1 ;
    wire \POWERLED.count_off_0_1 ;
    wire \POWERLED.func_state_RNI7LSV8Z0Z_0 ;
    wire \POWERLED.count_offZ0Z_1 ;
    wire N_7_cascade_;
    wire N_8_0_cascade_;
    wire \POWERLED.g0_5Z0Z_1_cascade_ ;
    wire POWERLED_g2_1_0_0;
    wire \POWERLED.N_74 ;
    wire \POWERLED.N_4_0_cascade_ ;
    wire \POWERLED.func_state_1_m2_0_0_0 ;
    wire \POWERLED.g1_0_0 ;
    wire \POWERLED.func_state_1_m2_N_3_7_1 ;
    wire clk_100Khz_signalkeep_3_fast;
    wire \POWERLED.N_671_0 ;
    wire G_7_i_a4_1_0_cascade_;
    wire \RSMRST_PWRGD.G_7_i_0 ;
    wire \POWERLED.N_533_cascade_ ;
    wire \POWERLED.N_533 ;
    wire \POWERLED.un1_clk_100khz_51_and_i_3_0_sx ;
    wire \POWERLED.un1_dutycycle_164_0_a3_0_a2_0 ;
    wire \POWERLED.count_clkZ0Z_7_cascade_ ;
    wire \POWERLED.un1_func_state25_6_0_o_N_4 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_9_0 ;
    wire \POWERLED.count_clk_0_7 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_5_cascade_ ;
    wire \POWERLED.un1_dutycycle_172_m3 ;
    wire \POWERLED.un1_clk_100khz_52_and_i_0_m2_ns_1_cascade_ ;
    wire \POWERLED.N_448_cascade_ ;
    wire \POWERLED.N_656_0 ;
    wire \POWERLED.N_133_cascade_ ;
    wire \POWERLED.un1_dutycycle_172_m4 ;
    wire \POWERLED.dutycycle_eena_14_c ;
    wire \POWERLED.N_488_cascade_ ;
    wire \POWERLED.un1_dutycycle_172_m2 ;
    wire \POWERLED.un1_clk_100khz_30_and_i_0_0_sx_cascade_ ;
    wire \POWERLED.func_state_1_m2s2_i_0_a2_1_0 ;
    wire \POWERLED.un1_dutycycle_96_0_a3_0_a2_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_3 ;
    wire \POWERLED.N_251_cascade_ ;
    wire \POWERLED.N_506 ;
    wire bfn_9_10_0_;
    wire \POWERLED.un1_dutycycle_94_cry_0_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_1_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_2_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_3_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_4 ;
    wire \POWERLED.un1_dutycycle_94_cry_5_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ;
    wire \POWERLED.un1_dutycycle_94_cry_6_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_7_cZ0 ;
    wire bfn_9_11_0_;
    wire \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61 ;
    wire \POWERLED.un1_dutycycle_94_cry_8 ;
    wire \POWERLED.un1_dutycycle_94_cry_9 ;
    wire \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_10 ;
    wire \POWERLED.un1_dutycycle_94_cry_11_cZ0 ;
    wire \POWERLED.dutycycleZ0Z_11 ;
    wire \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_12 ;
    wire \POWERLED.N_435_i ;
    wire \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_13_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_14 ;
    wire \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ;
    wire vccst_en;
    wire \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ;
    wire \POWERLED.dutycycle_RNIP1UTZ0Z_4_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_5_cascade_ ;
    wire \POWERLED.dutycycle_RNIF86R3Z0Z_4 ;
    wire \POWERLED.dutycycle_RNIP1UTZ0Z_4 ;
    wire \POWERLED.dutycycle_RNIF86R3Z0Z_4_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_4 ;
    wire \POWERLED.un1_dutycycle_53_31_0_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_9_3 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_11 ;
    wire \POWERLED.dutycycleZ1Z_8 ;
    wire \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ;
    wire \POWERLED.dutycycle_RNIRT5H5Z0Z_8 ;
    wire \POWERLED.dutycycleZ0Z_3_cascade_ ;
    wire \POWERLED.dutycycle_RNI_10_8_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_9_4 ;
    wire \POWERLED.un1_dutycycle_53_9_4_0 ;
    wire \POWERLED.un1_dutycycle_53_9_4_1 ;
    wire \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0 ;
    wire \POWERLED.dutycycleZ0Z_12 ;
    wire \POWERLED.dutycycleZ0Z_7_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_9_a0_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_10_4 ;
    wire \POWERLED.un1_dutycycle_53_40_0 ;
    wire \POWERLED.un1_dutycycle_53_axb_11_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_axb_11_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_14 ;
    wire \POWERLED.un1_dutycycle_53_45_0 ;
    wire \POWERLED.dutycycle_RNIZ0Z_4 ;
    wire \POWERLED.un1_dutycycle_53_35_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_22 ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_6 ;
    wire \POWERLED.dutycycle_RNI_10_8 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_6 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_6_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_35_1 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_6 ;
    wire \POWERLED.un1_dutycycle_53_50_a0_0 ;
    wire \POWERLED.un1_dutycycle_53_50_a0_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_50_a0_0_0 ;
    wire \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ;
    wire \POWERLED.dutycycle_en_4 ;
    wire \POWERLED.dutycycleZ1Z_10 ;
    wire \POWERLED.dutycycleZ0Z_2_cascade_ ;
    wire \POWERLED.un2_count_clk_17_0_0_a2_0_0 ;
    wire \POWERLED.un1_dutycycle_53_50_0_0 ;
    wire \POWERLED.un1_dutycycle_53_4_0 ;
    wire \POWERLED.un1_dutycycle_53_10_2_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_10_3 ;
    wire \POWERLED.un1_dutycycle_53_9_a1_0 ;
    wire \POWERLED.dutycycleZ0Z_2 ;
    wire \POWERLED.dutycycleZ0Z_9 ;
    wire \POWERLED.dutycycleZ0Z_3 ;
    wire \POWERLED.un1_dutycycle_53_50_3_0 ;
    wire \VPP_VDDQ.N_64_i ;
    wire \VPP_VDDQ.countZ0Z_0 ;
    wire bfn_11_2_0_;
    wire \VPP_VDDQ.countZ0Z_1 ;
    wire \VPP_VDDQ.un1_count_1_cry_0 ;
    wire \VPP_VDDQ.countZ0Z_2 ;
    wire \VPP_VDDQ.un1_count_1_cry_1 ;
    wire \VPP_VDDQ.countZ0Z_3 ;
    wire \VPP_VDDQ.un1_count_1_cry_2 ;
    wire \VPP_VDDQ.countZ0Z_4 ;
    wire \VPP_VDDQ.un1_count_1_cry_3 ;
    wire \VPP_VDDQ.countZ0Z_5 ;
    wire \VPP_VDDQ.un1_count_1_cry_4 ;
    wire \VPP_VDDQ.countZ0Z_6 ;
    wire \VPP_VDDQ.un1_count_1_cry_5 ;
    wire \VPP_VDDQ.countZ0Z_7 ;
    wire \VPP_VDDQ.un1_count_1_cry_6 ;
    wire \VPP_VDDQ.un1_count_1_cry_7 ;
    wire \VPP_VDDQ.countZ0Z_8 ;
    wire bfn_11_3_0_;
    wire \VPP_VDDQ.countZ0Z_9 ;
    wire \VPP_VDDQ.un1_count_1_cry_8 ;
    wire \VPP_VDDQ.countZ0Z_10 ;
    wire \VPP_VDDQ.un1_count_1_cry_9 ;
    wire \VPP_VDDQ.countZ0Z_11 ;
    wire \VPP_VDDQ.un1_count_1_cry_10 ;
    wire \VPP_VDDQ.countZ0Z_12 ;
    wire \VPP_VDDQ.un1_count_1_cry_11 ;
    wire \VPP_VDDQ.countZ0Z_13 ;
    wire \VPP_VDDQ.un1_count_1_cry_12 ;
    wire N_92_g;
    wire \VPP_VDDQ.countZ0Z_14 ;
    wire \VPP_VDDQ.un1_count_1_cry_13 ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \VPP_VDDQ.un1_count_1_cry_14 ;
    wire \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_11_4_0_;
    wire \VPP_VDDQ.countZ0Z_15 ;
    wire \VPP_VDDQ.N_92_0 ;
    wire G_30;
    wire \POWERLED.count_clk_0_4 ;
    wire \POWERLED.count_clk_0_5 ;
    wire \POWERLED.count_clk_0_6 ;
    wire clk_100Khz_signalkeep_3;
    wire clk_100Khz_signalkeep_3_rep1;
    wire \POWERLED.count_clk_RNIZ0Z_0_cascade_ ;
    wire \POWERLED.count_clkZ0Z_1_cascade_ ;
    wire \POWERLED.count_clk_0_1 ;
    wire \POWERLED.count_clk_0_11 ;
    wire \POWERLED.count_off_RNI_0Z0Z_10 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_8_3_cascade_ ;
    wire \POWERLED.N_668_cascade_ ;
    wire \POWERLED.N_490 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_1_cascade_ ;
    wire \POWERLED.N_123 ;
    wire \POWERLED.N_443 ;
    wire \POWERLED.count_off_RNIH9TEZ0Z_10 ;
    wire \POWERLED.un1_func_state25_6_0_0_0_2_1 ;
    wire \POWERLED.N_668 ;
    wire \POWERLED.count_off_1_sqmuxa ;
    wire \POWERLED.un1_dutycycle_172_m0 ;
    wire \POWERLED.un1_dutycycle_172_m1_ns_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_172_m1 ;
    wire \POWERLED.func_state_RNI_3Z0Z_1 ;
    wire N_247;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_2 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_1_cascade_ ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_4 ;
    wire \POWERLED.func_state_RNI_0Z0Z_1 ;
    wire func_state_RNI_4_1;
    wire func_state_RNI_0_0;
    wire \POWERLED.dutycycle_RNI_4Z0Z_0 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_0_cascade_ ;
    wire \POWERLED.dutycycle_N_3_mux_0 ;
    wire \POWERLED.N_546_cascade_ ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_0 ;
    wire \POWERLED.N_482 ;
    wire \POWERLED.g0_i_m2_rn_1_0 ;
    wire \POWERLED.dutycycleZ0Z_1_cascade_ ;
    wire \POWERLED.dutycycle_eena_0_0 ;
    wire \POWERLED.g0_1 ;
    wire \POWERLED.dutycycle_eena_0_0_cascade_ ;
    wire \POWERLED.dutycycle_eena_cascade_ ;
    wire \POWERLED.dutycycle ;
    wire \POWERLED.g0_i_m2_sn ;
    wire \POWERLED.func_stateZ0Z_0 ;
    wire \POWERLED.g0_i_m2_rn_1 ;
    wire \POWERLED.dutycycleZ1Z_1 ;
    wire \POWERLED.dutycycle_1_0_0 ;
    wire \POWERLED.dutycycle_eena ;
    wire \POWERLED.dutycycleZ1Z_0 ;
    wire \POWERLED.N_510 ;
    wire \POWERLED.un1_clk_100khz_36_and_i_0_a2_c_cascade_ ;
    wire rsmrst_pwrgd_signal;
    wire \POWERLED.un1_clk_100khz_36_and_i_0_a2_d ;
    wire \POWERLED.un1_clk_100khz_36_and_i_0_a2_1_0_2 ;
    wire \POWERLED.un1_clk_100khz_36_and_i_0_a2_1_d_cascade_ ;
    wire \POWERLED.dutycycle_eena_5 ;
    wire gpio_fpga_soc_4;
    wire \POWERLED.N_249_cascade_ ;
    wire \POWERLED.un1_clk_100khz_40_and_i_0_a2_1_0_3_1 ;
    wire \POWERLED.N_203_cascade_ ;
    wire \POWERLED.N_521_cascade_ ;
    wire \POWERLED.un1_clk_100khz_43_and_i_1_cascade_ ;
    wire \POWERLED.N_523 ;
    wire \POWERLED.N_503_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_4 ;
    wire \POWERLED.un1_clk_100khz_30_and_i_0_a2_5_0_0_cascade_ ;
    wire \POWERLED.dutycycle_eena_2_0_0_tz_1 ;
    wire \POWERLED.dutycycle_eena_2_d_0_cascade_ ;
    wire \POWERLED.dutycycle_RNIRUFD6Z0Z_9 ;
    wire \POWERLED.func_state_RNI2MQDZ0Z_1 ;
    wire RSMRSTn_rep1;
    wire \POWERLED.dutycycleZ1Z_6 ;
    wire \POWERLED.N_520_cascade_ ;
    wire \POWERLED.dutycycle_RNIRUFD6Z0Z_12 ;
    wire \POWERLED.dutycycleZ0Z_7 ;
    wire \POWERLED.N_518_cascade_ ;
    wire \POWERLED.un1_clk_100khz_42_and_i_1 ;
    wire \POWERLED.un1_clk_100khz_40_and_i_0_a2_1_d ;
    wire \POWERLED.N_526_cascade_ ;
    wire \POWERLED.dutycycle_RNI36306Z0Z_14 ;
    wire \POWERLED.func_state_RNI_8Z0Z_1 ;
    wire \POWERLED.N_203 ;
    wire \POWERLED.dutycycleZ0Z_10 ;
    wire \POWERLED.N_524_cascade_ ;
    wire \POWERLED.un1_clk_100khz_47_and_i_1 ;
    wire rsmrstn;
    wire \POWERLED.dutycycleZ0Z_14 ;
    wire \POWERLED.N_2381_i ;
    wire \POWERLED.N_91_1_N ;
    wire \POWERLED.N_527_cascade_ ;
    wire \POWERLED.un1_clk_100khz_48_and_i_1_cascade_ ;
    wire \POWERLED.N_529 ;
    wire \POWERLED.dutycycle_en_12 ;
    wire \POWERLED.count_clk_0_8 ;
    wire \POWERLED.count_clk_0_9 ;
    wire \POWERLED.count_clk_0_2 ;
    wire \POWERLED.count_clkZ0Z_3_cascade_ ;
    wire \POWERLED.un1_dutycycle_168_0_0_o2_4_cascade_ ;
    wire \POWERLED.count_clk_0_3 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_10_0_cascade_ ;
    wire \POWERLED.N_625 ;
    wire \POWERLED.count_clk_RNIZ0Z_1 ;
    wire \POWERLED.N_625_cascade_ ;
    wire \POWERLED.count_clk_RNIPGQN2_5Z0Z_3 ;
    wire \POWERLED.count_clkZ0Z_1 ;
    wire bfn_12_5_0_;
    wire \POWERLED.count_clkZ0Z_2 ;
    wire \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_1 ;
    wire \POWERLED.count_clkZ0Z_3 ;
    wire \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_2 ;
    wire \POWERLED.count_clkZ0Z_4 ;
    wire \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_3 ;
    wire \POWERLED.count_clkZ0Z_5 ;
    wire \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_4 ;
    wire \POWERLED.count_clkZ0Z_6 ;
    wire \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_5 ;
    wire \POWERLED.count_clkZ0Z_7 ;
    wire \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_6 ;
    wire \POWERLED.count_clkZ0Z_8 ;
    wire \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_7 ;
    wire \POWERLED.un1_count_clk_2_cry_8_cZ0 ;
    wire \POWERLED.count_clkZ0Z_9 ;
    wire \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ;
    wire bfn_12_6_0_;
    wire \POWERLED.un1_count_clk_2_cry_9 ;
    wire \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_10 ;
    wire \POWERLED.un1_count_clk_2_cry_11_cZ0 ;
    wire \POWERLED.un1_count_clk_2_cry_12 ;
    wire \POWERLED.un1_count_clk_2_cry_13_cZ0 ;
    wire \POWERLED.func_state_RNI2VV9A_0_0 ;
    wire \POWERLED.un1_count_clk_2_cry_14 ;
    wire \POWERLED.count_clk_0_15 ;
    wire \POWERLED.count_clk_1_15 ;
    wire \POWERLED.count_clkZ0Z_15 ;
    wire \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ;
    wire \POWERLED.count_clkZ0Z_10 ;
    wire \POWERLED.un1_count_clk_2_axb_10 ;
    wire \POWERLED.un1_count_clk_2_axb_14 ;
    wire \POWERLED.count_clk_0_0 ;
    wire \POWERLED.count_clk_RNI_0Z0Z_0 ;
    wire \POWERLED.count_clkZ0Z_0 ;
    wire \POWERLED.count_clk_1_14 ;
    wire \POWERLED.count_clkZ0Z_0_cascade_ ;
    wire \POWERLED.count_clkZ0Z_14 ;
    wire \POWERLED.count_clkZ0Z_11 ;
    wire \POWERLED.un2_count_clk_17_0_o2_1_1_cascade_ ;
    wire \POWERLED.un2_count_clk_17_0_o2_1_2 ;
    wire \POWERLED.count_clk_RNISLCE7Z0Z_10 ;
    wire \POWERLED.count_clk_en_917_0 ;
    wire \POWERLED.func_state_RNIBVNS_2Z0Z_0 ;
    wire \POWERLED.count_clk_en_1_cascade_ ;
    wire \POWERLED.N_617 ;
    wire \POWERLED.count_clk_en_cascade_ ;
    wire \POWERLED.un1_count_clk_2_axb_12 ;
    wire \POWERLED.count_clk_1_13 ;
    wire \POWERLED.count_clk_0_13 ;
    wire \POWERLED.count_clkZ0Z_13 ;
    wire \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ;
    wire \POWERLED.count_clk_en ;
    wire \POWERLED.count_clkZ0Z_13_cascade_ ;
    wire \POWERLED.count_clkZ0Z_12 ;
    wire \POWERLED.un2_count_clk_17_0_o2_1_0 ;
    wire \POWERLED.N_676 ;
    wire \POWERLED.N_492 ;
    wire \POWERLED.dutycycle_0_5 ;
    wire \POWERLED.func_state_RNIS28SBZ0Z_1 ;
    wire \POWERLED.dutycycleZ1Z_5_cascade_ ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_5_cascade_ ;
    wire \POWERLED.dutycycle_0_sqmuxa_i_i_a3_0_a2_0_cascade_ ;
    wire func_state_RNI_2_0;
    wire \POWERLED.un1_count_off_1_sqmuxa_8_ns_1 ;
    wire \POWERLED.dutycycle_RNI_8Z0Z_5_cascade_ ;
    wire \POWERLED.N_251 ;
    wire \POWERLED.N_633 ;
    wire \POWERLED.func_state_RNIOGRSZ0Z_1_cascade_ ;
    wire v5s_enn;
    wire \POWERLED.N_413_N ;
    wire \POWERLED.dutycycle_0_6 ;
    wire \POWERLED.dutycycleZ0Z_6_cascade_ ;
    wire \POWERLED.N_612 ;
    wire \POWERLED.N_672 ;
    wire \POWERLED.N_672_cascade_ ;
    wire \POWERLED.un1_dutycycle_168_0 ;
    wire \POWERLED.count_clk_RNIZ0Z_6 ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_0 ;
    wire \POWERLED.N_412_i_cascade_ ;
    wire \POWERLED.N_604 ;
    wire \POWERLED.dutycycle_RNI_6Z0Z_3 ;
    wire \POWERLED.N_435 ;
    wire \POWERLED.N_412_i ;
    wire \POWERLED.func_state_RNI_5Z0Z_1 ;
    wire \POWERLED.func_state_RNI_5Z0Z_1_cascade_ ;
    wire \POWERLED.N_23_i ;
    wire \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ;
    wire \POWERLED.N_85 ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_5 ;
    wire \POWERLED.func_state_RNI12ASZ0Z_1_cascade_ ;
    wire \POWERLED.N_613 ;
    wire slp_s4n;
    wire \POWERLED.func_state_RNI8AQHZ0Z_0 ;
    wire \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ;
    wire \POWERLED.func_state_RNI12ASZ0Z_1 ;
    wire \POWERLED.N_83 ;
    wire slp_s3n;
    wire func_state_RNIMJ6IF_0_1;
    wire RSMRSTn_rep2;
    wire \POWERLED.N_531 ;
    wire \POWERLED.un1_clk_100khz_51_and_i_3_0 ;
    wire \POWERLED.N_532_cascade_ ;
    wire \POWERLED.N_530 ;
    wire \POWERLED.dutycycle_eena_13_c_1 ;
    wire \POWERLED.N_430 ;
    wire \POWERLED.un1_clk_100khz_51_and_i_3_cascade_ ;
    wire G_141;
    wire \POWERLED.dutycycle_RNI0DF58Z0Z_5 ;
    wire fpga_osc;
    wire \POWERLED.N_430_iZ0 ;
    wire \POWERLED.dutycycle_en_8 ;
    wire \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ;
    wire \POWERLED.dutycycleZ1Z_3 ;
    wire \POWERLED.N_421 ;
    wire \POWERLED.dutycycleZ0Z_8_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_axb_3_1_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_5 ;
    wire \POWERLED.dutycycleZ1Z_5 ;
    wire \POWERLED.un1_i3_mux_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_3 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_5 ;
    wire \POWERLED.dutycycleZ0Z_6 ;
    wire \POWERLED.dutycycleZ0Z_8 ;
    wire \POWERLED.dutycycleZ0Z_1 ;
    wire \POWERLED.d_i3_mux ;
    wire \VPP_VDDQ.delayed_vddq_pwrgdZ0 ;
    wire VCCST_EN_i_1;
    wire vpp_en;
    wire vccst_cpu_ok;
    wire v5s_ok;
    wire \VCCIN_PWRGD.un10_outputZ0Z_1 ;
    wire v33s_ok;
    wire vccin_en;
    wire \POWERLED.dutycycleZ0Z_0 ;
    wire \POWERLED.un1_dutycycle_53_axb_3 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_2 ;
    wire _gnd_net_;

    defparam ipInertedIOPad_VR_READY_VCCINAUX_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VR_READY_VCCINAUX_iopad (
            .OE(N__33702),
            .DIN(N__33701),
            .DOUT(N__33700),
            .PACKAGEPIN(VR_READY_VCCINAUX));
    defparam ipInertedIOPad_VR_READY_VCCINAUX_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCINAUX_preio (
            .PADOEN(N__33702),
            .PADOUT(N__33701),
            .PADIN(N__33700),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_ENn_iopad (
            .OE(N__33693),
            .DIN(N__33692),
            .DOUT(N__33691),
            .PACKAGEPIN(V33A_ENn));
    defparam ipInertedIOPad_V33A_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33A_ENn_preio (
            .PADOEN(N__33693),
            .PADOUT(N__33692),
            .PADIN(N__33691),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__15680),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V1P8A_EN_iopad (
            .OE(N__33684),
            .DIN(N__33683),
            .DOUT(N__33682),
            .PACKAGEPIN(V1P8A_EN));
    defparam ipInertedIOPad_V1P8A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V1P8A_EN_preio (
            .PADOEN(N__33684),
            .PADOUT(N__33683),
            .PADIN(N__33682),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16225),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDDQ_EN_iopad (
            .OE(N__33675),
            .DIN(N__33674),
            .DOUT(N__33673),
            .PACKAGEPIN(VDDQ_EN));
    defparam ipInertedIOPad_VDDQ_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDDQ_EN_preio (
            .PADOEN(N__33675),
            .PADOUT(N__33674),
            .PADIN(N__33673),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__14081),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad (
            .OE(N__33666),
            .DIN(N__33665),
            .DOUT(N__33664),
            .PACKAGEPIN(VCCST_OVERRIDE_3V3));
    defparam ipInertedIOPad_VCCST_OVERRIDE_3V3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_OVERRIDE_3V3_preio (
            .PADOEN(N__33666),
            .PADOUT(N__33665),
            .PADIN(N__33664),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_OK_iopad (
            .OE(N__33657),
            .DIN(N__33656),
            .DOUT(N__33655),
            .PACKAGEPIN(V5S_OK));
    defparam ipInertedIOPad_V5S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5S_OK_preio (
            .PADOEN(N__33657),
            .PADOUT(N__33656),
            .PADIN(N__33655),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S3n_iopad (
            .OE(N__33648),
            .DIN(N__33647),
            .DOUT(N__33646),
            .PACKAGEPIN(SLP_S3n));
    defparam ipInertedIOPad_SLP_S3n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S3n_preio (
            .PADOEN(N__33648),
            .PADOUT(N__33647),
            .PADIN(N__33646),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s3n),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S0n_iopad (
            .OE(N__33639),
            .DIN(N__33638),
            .DOUT(N__33637),
            .PACKAGEPIN(SLP_S0n));
    defparam ipInertedIOPad_SLP_S0n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S0n_preio (
            .PADOEN(N__33639),
            .PADOUT(N__33638),
            .PADIN(N__33637),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_ENn_iopad (
            .OE(N__33630),
            .DIN(N__33629),
            .DOUT(N__33628),
            .PACKAGEPIN(V5S_ENn));
    defparam ipInertedIOPad_V5S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5S_ENn_preio (
            .PADOEN(N__33630),
            .PADOUT(N__33629),
            .PADIN(N__33628),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29626),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V1P8A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V1P8A_OK_iopad (
            .OE(N__33621),
            .DIN(N__33620),
            .DOUT(N__33619),
            .PACKAGEPIN(V1P8A_OK));
    defparam ipInertedIOPad_V1P8A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V1P8A_OK_preio (
            .PADOEN(N__33621),
            .PADOUT(N__33620),
            .PADIN(N__33619),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v1p8a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTNn_iopad (
            .OE(N__33612),
            .DIN(N__33611),
            .DOUT(N__33610),
            .PACKAGEPIN(PWRBTNn));
    defparam ipInertedIOPad_PWRBTNn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PWRBTNn_preio (
            .PADOEN(N__33612),
            .PADOUT(N__33611),
            .PADIN(N__33610),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTN_LED_iopad (
            .OE(N__33603),
            .DIN(N__33602),
            .DOUT(N__33601),
            .PACKAGEPIN(PWRBTN_LED));
    defparam ipInertedIOPad_PWRBTN_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PWRBTN_LED_preio (
            .PADOEN(N__33603),
            .PADOUT(N__33602),
            .PADIN(N__33601),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__14102),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_2_iopad (
            .OE(N__33594),
            .DIN(N__33593),
            .DOUT(N__33592),
            .PACKAGEPIN(GPIO_FPGA_SoC_2));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_2_preio (
            .PADOEN(N__33594),
            .PADOUT(N__33593),
            .PADIN(N__33592),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad (
            .OE(N__33585),
            .DIN(N__33584),
            .DOUT(N__33583),
            .PACKAGEPIN(VCCIN_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__33585),
            .PADOUT(N__33584),
            .PADIN(N__33583),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_SLP_SUSn_iopad.PULLUP=1'b0;
    IO_PAD ipInertedIOPad_SLP_SUSn_iopad (
            .OE(N__33576),
            .DIN(N__33575),
            .DOUT(N__33574),
            .PACKAGEPIN(SLP_SUSn));
    defparam ipInertedIOPad_SLP_SUSn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_SUSn_preio (
            .PADOEN(N__33576),
            .PADOUT(N__33575),
            .PADIN(N__33574),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_susn),
            .DIN1());
    IO_PAD ipInertedIOPad_CPU_C10_GATE_N_iopad (
            .OE(N__33567),
            .DIN(N__33566),
            .DOUT(N__33565),
            .PACKAGEPIN(CPU_C10_GATE_N));
    defparam ipInertedIOPad_CPU_C10_GATE_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_CPU_C10_GATE_N_preio (
            .PADOEN(N__33567),
            .PADOUT(N__33566),
            .PADIN(N__33565),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_EN_iopad (
            .OE(N__33558),
            .DIN(N__33557),
            .DOUT(N__33556),
            .PACKAGEPIN(VCCST_EN));
    defparam ipInertedIOPad_VCCST_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_EN_preio (
            .PADOEN(N__33558),
            .PADOUT(N__33557),
            .PADIN(N__33556),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23918),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V33DSW_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V33DSW_OK_iopad (
            .OE(N__33549),
            .DIN(N__33548),
            .DOUT(N__33547),
            .PACKAGEPIN(V33DSW_OK));
    defparam ipInertedIOPad_V33DSW_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33DSW_OK_preio (
            .PADOEN(N__33549),
            .PADOUT(N__33548),
            .PADIN(N__33547),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_TPM_GPIO_iopad (
            .OE(N__33540),
            .DIN(N__33539),
            .DOUT(N__33538),
            .PACKAGEPIN(TPM_GPIO));
    defparam ipInertedIOPad_TPM_GPIO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_TPM_GPIO_preio (
            .PADOEN(N__33540),
            .PADOUT(N__33539),
            .PADIN(N__33538),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSWARN_N_iopad (
            .OE(N__33531),
            .DIN(N__33530),
            .DOUT(N__33529),
            .PACKAGEPIN(SUSWARN_N));
    defparam ipInertedIOPad_SUSWARN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSWARN_N_preio (
            .PADOEN(N__33531),
            .PADOUT(N__33530),
            .PADIN(N__33529),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PLTRSTn_iopad (
            .OE(N__33522),
            .DIN(N__33521),
            .DOUT(N__33520),
            .PACKAGEPIN(PLTRSTn));
    defparam ipInertedIOPad_PLTRSTn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PLTRSTn_preio (
            .PADOEN(N__33522),
            .PADOUT(N__33521),
            .PADIN(N__33520),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_4_iopad (
            .OE(N__33513),
            .DIN(N__33512),
            .DOUT(N__33511),
            .PACKAGEPIN(GPIO_FPGA_SoC_4));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_4_preio (
            .PADOEN(N__33513),
            .PADOUT(N__33512),
            .PADIN(N__33511),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_4),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_READY_VCCIN_iopad (
            .OE(N__33504),
            .DIN(N__33503),
            .DOUT(N__33502),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam ipInertedIOPad_VR_READY_VCCIN_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCIN_preio (
            .PADOEN(N__33504),
            .PADOUT(N__33503),
            .PADIN(N__33502),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccin),
            .DIN1());
    defparam ipInertedIOPad_V5A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V5A_OK_iopad (
            .OE(N__33495),
            .DIN(N__33494),
            .DOUT(N__33493),
            .PACKAGEPIN(V5A_OK));
    defparam ipInertedIOPad_V5A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5A_OK_preio (
            .PADOEN(N__33495),
            .PADOUT(N__33494),
            .PADIN(N__33493),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_RSMRSTn_iopad (
            .OE(N__33486),
            .DIN(N__33485),
            .DOUT(N__33484),
            .PACKAGEPIN(RSMRSTn));
    defparam ipInertedIOPad_RSMRSTn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RSMRSTn_preio (
            .PADOEN(N__33486),
            .PADOUT(N__33485),
            .PADIN(N__33484),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27692),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_OSC_iopad (
            .OE(N__33477),
            .DIN(N__33476),
            .DOUT(N__33475),
            .PACKAGEPIN(FPGA_OSC));
    defparam ipInertedIOPad_FPGA_OSC_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_OSC_preio (
            .PADOEN(N__33477),
            .PADOUT(N__33476),
            .PADIN(N__33475),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(fpga_osc),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_PWRGD_iopad (
            .OE(N__33468),
            .DIN(N__33467),
            .DOUT(N__33466),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam ipInertedIOPad_VCCST_PWRGD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_PWRGD_preio (
            .PADOEN(N__33468),
            .PADOUT(N__33467),
            .PADIN(N__33466),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__15461),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SYS_PWROK_iopad (
            .OE(N__33459),
            .DIN(N__33458),
            .DOUT(N__33457),
            .PACKAGEPIN(SYS_PWROK));
    defparam ipInertedIOPad_SYS_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SYS_PWROK_preio (
            .PADOEN(N__33459),
            .PADOUT(N__33458),
            .PADIN(N__33457),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__15439),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO2_iopad (
            .OE(N__33450),
            .DIN(N__33449),
            .DOUT(N__33448),
            .PACKAGEPIN(SPI_FP_IO2));
    defparam ipInertedIOPad_SPI_FP_IO2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO2_preio (
            .PADOEN(N__33450),
            .PADOUT(N__33449),
            .PADIN(N__33448),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE1_FPGA_iopad (
            .OE(N__33441),
            .DIN(N__33440),
            .DOUT(N__33439),
            .PACKAGEPIN(SATAXPCIE1_FPGA));
    defparam ipInertedIOPad_SATAXPCIE1_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE1_FPGA_preio (
            .PADOEN(N__33441),
            .PADOUT(N__33440),
            .PADIN(N__33439),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_1_iopad (
            .OE(N__33432),
            .DIN(N__33431),
            .DOUT(N__33430),
            .PACKAGEPIN(GPIO_FPGA_EXP_1));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_1_preio (
            .PADOEN(N__33432),
            .PADOUT(N__33431),
            .PADIN(N__33430),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad (
            .OE(N__33423),
            .DIN(N__33422),
            .DOUT(N__33421),
            .PACKAGEPIN(VCCINAUX_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__33423),
            .PADOUT(N__33422),
            .PADIN(N__33421),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PE_iopad (
            .OE(N__33414),
            .DIN(N__33413),
            .DOUT(N__33412),
            .PACKAGEPIN(VCCINAUX_VR_PE));
    defparam ipInertedIOPad_VCCINAUX_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PE_preio (
            .PADOEN(N__33414),
            .PADOUT(N__33413),
            .PADIN(N__33412),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_HDA_SDO_ATP_iopad (
            .OE(N__33405),
            .DIN(N__33404),
            .DOUT(N__33403),
            .PACKAGEPIN(HDA_SDO_ATP));
    defparam ipInertedIOPad_HDA_SDO_ATP_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_HDA_SDO_ATP_preio (
            .PADOEN(N__33405),
            .PADOUT(N__33404),
            .PADIN(N__33403),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__15884),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_2_iopad (
            .OE(N__33396),
            .DIN(N__33395),
            .DOUT(N__33394),
            .PACKAGEPIN(GPIO_FPGA_EXP_2));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_2_preio (
            .PADOEN(N__33396),
            .PADOUT(N__33395),
            .PADIN(N__33394),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VPP_EN_iopad (
            .OE(N__33387),
            .DIN(N__33386),
            .DOUT(N__33385),
            .PACKAGEPIN(VPP_EN));
    defparam ipInertedIOPad_VPP_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VPP_EN_preio (
            .PADOEN(N__33387),
            .PADOUT(N__33386),
            .PADIN(N__33385),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__33026),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VDDQ_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VDDQ_OK_iopad (
            .OE(N__33378),
            .DIN(N__33377),
            .DOUT(N__33376),
            .PACKAGEPIN(VDDQ_OK));
    defparam ipInertedIOPad_VDDQ_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDDQ_OK_preio (
            .PADOEN(N__33378),
            .PADOUT(N__33377),
            .PADIN(N__33376),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vddq_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSACK_N_iopad (
            .OE(N__33369),
            .DIN(N__33368),
            .DOUT(N__33367),
            .PACKAGEPIN(SUSACK_N));
    defparam ipInertedIOPad_SUSACK_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSACK_N_preio (
            .PADOEN(N__33369),
            .PADOUT(N__33368),
            .PADIN(N__33367),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S4n_iopad (
            .OE(N__33360),
            .DIN(N__33359),
            .DOUT(N__33358),
            .PACKAGEPIN(SLP_S4n));
    defparam ipInertedIOPad_SLP_S4n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S4n_preio (
            .PADOEN(N__33360),
            .PADOUT(N__33359),
            .PADIN(N__33358),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s4n),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_CPU_OK_iopad (
            .OE(N__33351),
            .DIN(N__33350),
            .DOUT(N__33349),
            .PACKAGEPIN(VCCST_CPU_OK));
    defparam ipInertedIOPad_VCCST_CPU_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_CPU_OK_preio (
            .PADOEN(N__33351),
            .PADOUT(N__33350),
            .PADIN(N__33349),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vccst_cpu_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_EN_iopad (
            .OE(N__33342),
            .DIN(N__33341),
            .DOUT(N__33340),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam ipInertedIOPad_VCCINAUX_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_EN_preio (
            .PADOEN(N__33342),
            .PADOUT(N__33341),
            .PADIN(N__33340),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16181),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_OK_iopad (
            .OE(N__33333),
            .DIN(N__33332),
            .DOUT(N__33331),
            .PACKAGEPIN(V33S_OK));
    defparam ipInertedIOPad_V33S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33S_OK_preio (
            .PADOEN(N__33333),
            .PADOUT(N__33332),
            .PADIN(N__33331),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_ENn_iopad (
            .OE(N__33324),
            .DIN(N__33323),
            .DOUT(N__33322),
            .PACKAGEPIN(V33S_ENn));
    defparam ipInertedIOPad_V33S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33S_ENn_preio (
            .PADOEN(N__33324),
            .PADOUT(N__33323),
            .PADIN(N__33322),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29630),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_1_iopad (
            .OE(N__33315),
            .DIN(N__33314),
            .DOUT(N__33313),
            .PACKAGEPIN(GPIO_FPGA_SoC_1));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_1_preio (
            .PADOEN(N__33315),
            .PADOUT(N__33314),
            .PADIN(N__33313),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_1),
            .DIN1());
    defparam ipInertedIOPad_DSW_PWROK_iopad.PULLUP=1'b0;
    IO_PAD ipInertedIOPad_DSW_PWROK_iopad (
            .OE(N__33306),
            .DIN(N__33305),
            .DOUT(N__33304),
            .PACKAGEPIN(DSW_PWROK));
    defparam ipInertedIOPad_DSW_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DSW_PWROK_preio (
            .PADOEN(N__33306),
            .PADOUT(N__33305),
            .PADIN(N__33304),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25181),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5A_EN_iopad (
            .OE(N__33297),
            .DIN(N__33296),
            .DOUT(N__33295),
            .PACKAGEPIN(V5A_EN));
    defparam ipInertedIOPad_V5A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5A_EN_preio (
            .PADOEN(N__33297),
            .PADOUT(N__33296),
            .PADIN(N__33295),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16226),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_3_iopad (
            .OE(N__33288),
            .DIN(N__33287),
            .DOUT(N__33286),
            .PACKAGEPIN(GPIO_FPGA_SoC_3));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_3_preio (
            .PADOEN(N__33288),
            .PADOUT(N__33287),
            .PADIN(N__33286),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad (
            .OE(N__33279),
            .DIN(N__33278),
            .DOUT(N__33277),
            .PACKAGEPIN(VR_PROCHOT_FPGA_OUT_N));
    defparam ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio (
            .PADOEN(N__33279),
            .PADOUT(N__33278),
            .PADIN(N__33277),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VPP_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VPP_OK_iopad (
            .OE(N__33270),
            .DIN(N__33269),
            .DOUT(N__33268),
            .PACKAGEPIN(VPP_OK));
    defparam ipInertedIOPad_VPP_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VPP_OK_preio (
            .PADOEN(N__33270),
            .PADOUT(N__33269),
            .PADIN(N__33268),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vpp_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PE_iopad (
            .OE(N__33261),
            .DIN(N__33260),
            .DOUT(N__33259),
            .PACKAGEPIN(VCCIN_VR_PE));
    defparam ipInertedIOPad_VCCIN_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PE_preio (
            .PADOEN(N__33261),
            .PADOUT(N__33260),
            .PADIN(N__33259),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25202),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_EN_iopad (
            .OE(N__33252),
            .DIN(N__33251),
            .DOUT(N__33250),
            .PACKAGEPIN(VCCIN_EN));
    defparam ipInertedIOPad_VCCIN_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_EN_preio (
            .PADOEN(N__33252),
            .PADOUT(N__33251),
            .PADIN(N__33250),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__32969),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SOC_SPKR_iopad (
            .OE(N__33243),
            .DIN(N__33242),
            .DOUT(N__33241),
            .PACKAGEPIN(SOC_SPKR));
    defparam ipInertedIOPad_SOC_SPKR_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SOC_SPKR_preio (
            .PADOEN(N__33243),
            .PADOUT(N__33242),
            .PADIN(N__33241),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S5n_iopad (
            .OE(N__33234),
            .DIN(N__33233),
            .DOUT(N__33232),
            .PACKAGEPIN(SLP_S5n));
    defparam ipInertedIOPad_SLP_S5n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S5n_preio (
            .PADOEN(N__33234),
            .PADOUT(N__33233),
            .PADIN(N__33232),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V12_MAIN_MON_iopad (
            .OE(N__33225),
            .DIN(N__33224),
            .DOUT(N__33223),
            .PACKAGEPIN(V12_MAIN_MON));
    defparam ipInertedIOPad_V12_MAIN_MON_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V12_MAIN_MON_preio (
            .PADOEN(N__33225),
            .PADOUT(N__33224),
            .PADIN(N__33223),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO3_iopad (
            .OE(N__33216),
            .DIN(N__33215),
            .DOUT(N__33214),
            .PACKAGEPIN(SPI_FP_IO3));
    defparam ipInertedIOPad_SPI_FP_IO3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO3_preio (
            .PADOEN(N__33216),
            .PADOUT(N__33215),
            .PADIN(N__33214),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE0_FPGA_iopad (
            .OE(N__33207),
            .DIN(N__33206),
            .DOUT(N__33205),
            .PACKAGEPIN(SATAXPCIE0_FPGA));
    defparam ipInertedIOPad_SATAXPCIE0_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE0_FPGA_preio (
            .PADOEN(N__33207),
            .PADOUT(N__33206),
            .PADIN(N__33205),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_OK_iopad (
            .OE(N__33198),
            .DIN(N__33197),
            .DOUT(N__33196),
            .PACKAGEPIN(V33A_OK));
    defparam ipInertedIOPad_V33A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33A_OK_preio (
            .PADOEN(N__33198),
            .PADOUT(N__33197),
            .PADIN(N__33196),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PCH_PWROK_iopad (
            .OE(N__33189),
            .DIN(N__33188),
            .DOUT(N__33187),
            .PACKAGEPIN(PCH_PWROK));
    defparam ipInertedIOPad_PCH_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PCH_PWROK_preio (
            .PADOEN(N__33189),
            .PADOUT(N__33188),
            .PADIN(N__33187),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__15440),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_SLP_WLAN_N_iopad (
            .OE(N__33180),
            .DIN(N__33179),
            .DOUT(N__33178),
            .PACKAGEPIN(FPGA_SLP_WLAN_N));
    defparam ipInertedIOPad_FPGA_SLP_WLAN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_SLP_WLAN_N_preio (
            .PADOEN(N__33180),
            .PADOUT(N__33179),
            .PADIN(N__33178),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    InMux I__7709 (
            .O(N__33161),
            .I(N__33158));
    LocalMux I__7708 (
            .O(N__33158),
            .I(N__33155));
    Span4Mux_v I__7707 (
            .O(N__33155),
            .I(N__33152));
    Span4Mux_h I__7706 (
            .O(N__33152),
            .I(N__33149));
    Span4Mux_v I__7705 (
            .O(N__33149),
            .I(N__33146));
    Span4Mux_v I__7704 (
            .O(N__33146),
            .I(N__33141));
    InMux I__7703 (
            .O(N__33145),
            .I(N__33136));
    InMux I__7702 (
            .O(N__33144),
            .I(N__33136));
    Odrv4 I__7701 (
            .O(N__33141),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    LocalMux I__7700 (
            .O(N__33136),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    InMux I__7699 (
            .O(N__33131),
            .I(N__33124));
    InMux I__7698 (
            .O(N__33130),
            .I(N__33120));
    InMux I__7697 (
            .O(N__33129),
            .I(N__33117));
    InMux I__7696 (
            .O(N__33128),
            .I(N__33112));
    InMux I__7695 (
            .O(N__33127),
            .I(N__33112));
    LocalMux I__7694 (
            .O(N__33124),
            .I(N__33109));
    InMux I__7693 (
            .O(N__33123),
            .I(N__33106));
    LocalMux I__7692 (
            .O(N__33120),
            .I(N__33101));
    LocalMux I__7691 (
            .O(N__33117),
            .I(N__33101));
    LocalMux I__7690 (
            .O(N__33112),
            .I(N__33098));
    Span4Mux_v I__7689 (
            .O(N__33109),
            .I(N__33095));
    LocalMux I__7688 (
            .O(N__33106),
            .I(N__33092));
    Span4Mux_v I__7687 (
            .O(N__33101),
            .I(N__33087));
    Span4Mux_s2_v I__7686 (
            .O(N__33098),
            .I(N__33087));
    Span4Mux_h I__7685 (
            .O(N__33095),
            .I(N__33081));
    Span4Mux_v I__7684 (
            .O(N__33092),
            .I(N__33078));
    Span4Mux_h I__7683 (
            .O(N__33087),
            .I(N__33074));
    InMux I__7682 (
            .O(N__33086),
            .I(N__33069));
    InMux I__7681 (
            .O(N__33085),
            .I(N__33069));
    CascadeMux I__7680 (
            .O(N__33084),
            .I(N__33064));
    Span4Mux_v I__7679 (
            .O(N__33081),
            .I(N__33060));
    Span4Mux_h I__7678 (
            .O(N__33078),
            .I(N__33057));
    InMux I__7677 (
            .O(N__33077),
            .I(N__33054));
    Span4Mux_v I__7676 (
            .O(N__33074),
            .I(N__33049));
    LocalMux I__7675 (
            .O(N__33069),
            .I(N__33049));
    InMux I__7674 (
            .O(N__33068),
            .I(N__33044));
    InMux I__7673 (
            .O(N__33067),
            .I(N__33044));
    InMux I__7672 (
            .O(N__33064),
            .I(N__33039));
    InMux I__7671 (
            .O(N__33063),
            .I(N__33039));
    Odrv4 I__7670 (
            .O(N__33060),
            .I(VCCST_EN_i_1));
    Odrv4 I__7669 (
            .O(N__33057),
            .I(VCCST_EN_i_1));
    LocalMux I__7668 (
            .O(N__33054),
            .I(VCCST_EN_i_1));
    Odrv4 I__7667 (
            .O(N__33049),
            .I(VCCST_EN_i_1));
    LocalMux I__7666 (
            .O(N__33044),
            .I(VCCST_EN_i_1));
    LocalMux I__7665 (
            .O(N__33039),
            .I(VCCST_EN_i_1));
    IoInMux I__7664 (
            .O(N__33026),
            .I(N__33023));
    LocalMux I__7663 (
            .O(N__33023),
            .I(vpp_en));
    InMux I__7662 (
            .O(N__33020),
            .I(N__33017));
    LocalMux I__7661 (
            .O(N__33017),
            .I(N__33014));
    Span4Mux_s2_h I__7660 (
            .O(N__33014),
            .I(N__33011));
    Sp12to4 I__7659 (
            .O(N__33011),
            .I(N__33008));
    Span12Mux_v I__7658 (
            .O(N__33008),
            .I(N__33005));
    Odrv12 I__7657 (
            .O(N__33005),
            .I(vccst_cpu_ok));
    InMux I__7656 (
            .O(N__33002),
            .I(N__32999));
    LocalMux I__7655 (
            .O(N__32999),
            .I(N__32996));
    IoSpan4Mux I__7654 (
            .O(N__32996),
            .I(N__32993));
    IoSpan4Mux I__7653 (
            .O(N__32993),
            .I(N__32990));
    Odrv4 I__7652 (
            .O(N__32990),
            .I(v5s_ok));
    CascadeMux I__7651 (
            .O(N__32987),
            .I(N__32984));
    InMux I__7650 (
            .O(N__32984),
            .I(N__32981));
    LocalMux I__7649 (
            .O(N__32981),
            .I(N__32978));
    Odrv4 I__7648 (
            .O(N__32978),
            .I(\VCCIN_PWRGD.un10_outputZ0Z_1 ));
    InMux I__7647 (
            .O(N__32975),
            .I(N__32972));
    LocalMux I__7646 (
            .O(N__32972),
            .I(v33s_ok));
    IoInMux I__7645 (
            .O(N__32969),
            .I(N__32966));
    LocalMux I__7644 (
            .O(N__32966),
            .I(N__32963));
    Span4Mux_s3_v I__7643 (
            .O(N__32963),
            .I(N__32960));
    Odrv4 I__7642 (
            .O(N__32960),
            .I(vccin_en));
    CascadeMux I__7641 (
            .O(N__32957),
            .I(N__32950));
    CascadeMux I__7640 (
            .O(N__32956),
            .I(N__32945));
    InMux I__7639 (
            .O(N__32955),
            .I(N__32941));
    InMux I__7638 (
            .O(N__32954),
            .I(N__32937));
    InMux I__7637 (
            .O(N__32953),
            .I(N__32934));
    InMux I__7636 (
            .O(N__32950),
            .I(N__32929));
    InMux I__7635 (
            .O(N__32949),
            .I(N__32929));
    InMux I__7634 (
            .O(N__32948),
            .I(N__32926));
    InMux I__7633 (
            .O(N__32945),
            .I(N__32923));
    InMux I__7632 (
            .O(N__32944),
            .I(N__32920));
    LocalMux I__7631 (
            .O(N__32941),
            .I(N__32917));
    CascadeMux I__7630 (
            .O(N__32940),
            .I(N__32914));
    LocalMux I__7629 (
            .O(N__32937),
            .I(N__32910));
    LocalMux I__7628 (
            .O(N__32934),
            .I(N__32905));
    LocalMux I__7627 (
            .O(N__32929),
            .I(N__32905));
    LocalMux I__7626 (
            .O(N__32926),
            .I(N__32902));
    LocalMux I__7625 (
            .O(N__32923),
            .I(N__32899));
    LocalMux I__7624 (
            .O(N__32920),
            .I(N__32896));
    Span12Mux_s7_h I__7623 (
            .O(N__32917),
            .I(N__32893));
    InMux I__7622 (
            .O(N__32914),
            .I(N__32890));
    InMux I__7621 (
            .O(N__32913),
            .I(N__32887));
    Span4Mux_v I__7620 (
            .O(N__32910),
            .I(N__32880));
    Span4Mux_v I__7619 (
            .O(N__32905),
            .I(N__32880));
    Span4Mux_v I__7618 (
            .O(N__32902),
            .I(N__32880));
    Span4Mux_s3_h I__7617 (
            .O(N__32899),
            .I(N__32875));
    Span4Mux_s3_h I__7616 (
            .O(N__32896),
            .I(N__32875));
    Odrv12 I__7615 (
            .O(N__32893),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__7614 (
            .O(N__32890),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__7613 (
            .O(N__32887),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__7612 (
            .O(N__32880),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__7611 (
            .O(N__32875),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    InMux I__7610 (
            .O(N__32864),
            .I(N__32861));
    LocalMux I__7609 (
            .O(N__32861),
            .I(\POWERLED.un1_dutycycle_53_axb_3 ));
    InMux I__7608 (
            .O(N__32858),
            .I(N__32855));
    LocalMux I__7607 (
            .O(N__32855),
            .I(N__32852));
    Odrv12 I__7606 (
            .O(N__32852),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_2 ));
    InMux I__7605 (
            .O(N__32849),
            .I(N__32846));
    LocalMux I__7604 (
            .O(N__32846),
            .I(\POWERLED.dutycycle_eena_13_c_1 ));
    InMux I__7603 (
            .O(N__32843),
            .I(N__32837));
    InMux I__7602 (
            .O(N__32842),
            .I(N__32837));
    LocalMux I__7601 (
            .O(N__32837),
            .I(N__32828));
    CascadeMux I__7600 (
            .O(N__32836),
            .I(N__32822));
    InMux I__7599 (
            .O(N__32835),
            .I(N__32816));
    InMux I__7598 (
            .O(N__32834),
            .I(N__32816));
    InMux I__7597 (
            .O(N__32833),
            .I(N__32806));
    InMux I__7596 (
            .O(N__32832),
            .I(N__32806));
    InMux I__7595 (
            .O(N__32831),
            .I(N__32803));
    Span4Mux_s1_v I__7594 (
            .O(N__32828),
            .I(N__32800));
    InMux I__7593 (
            .O(N__32827),
            .I(N__32797));
    InMux I__7592 (
            .O(N__32826),
            .I(N__32794));
    InMux I__7591 (
            .O(N__32825),
            .I(N__32789));
    InMux I__7590 (
            .O(N__32822),
            .I(N__32784));
    InMux I__7589 (
            .O(N__32821),
            .I(N__32784));
    LocalMux I__7588 (
            .O(N__32816),
            .I(N__32780));
    InMux I__7587 (
            .O(N__32815),
            .I(N__32775));
    InMux I__7586 (
            .O(N__32814),
            .I(N__32775));
    InMux I__7585 (
            .O(N__32813),
            .I(N__32772));
    InMux I__7584 (
            .O(N__32812),
            .I(N__32769));
    InMux I__7583 (
            .O(N__32811),
            .I(N__32765));
    LocalMux I__7582 (
            .O(N__32806),
            .I(N__32754));
    LocalMux I__7581 (
            .O(N__32803),
            .I(N__32754));
    Span4Mux_h I__7580 (
            .O(N__32800),
            .I(N__32754));
    LocalMux I__7579 (
            .O(N__32797),
            .I(N__32754));
    LocalMux I__7578 (
            .O(N__32794),
            .I(N__32754));
    InMux I__7577 (
            .O(N__32793),
            .I(N__32749));
    InMux I__7576 (
            .O(N__32792),
            .I(N__32749));
    LocalMux I__7575 (
            .O(N__32789),
            .I(N__32746));
    LocalMux I__7574 (
            .O(N__32784),
            .I(N__32741));
    InMux I__7573 (
            .O(N__32783),
            .I(N__32737));
    Span4Mux_v I__7572 (
            .O(N__32780),
            .I(N__32732));
    LocalMux I__7571 (
            .O(N__32775),
            .I(N__32732));
    LocalMux I__7570 (
            .O(N__32772),
            .I(N__32727));
    LocalMux I__7569 (
            .O(N__32769),
            .I(N__32727));
    InMux I__7568 (
            .O(N__32768),
            .I(N__32724));
    LocalMux I__7567 (
            .O(N__32765),
            .I(N__32715));
    Span4Mux_v I__7566 (
            .O(N__32754),
            .I(N__32715));
    LocalMux I__7565 (
            .O(N__32749),
            .I(N__32715));
    Span4Mux_s1_h I__7564 (
            .O(N__32746),
            .I(N__32715));
    InMux I__7563 (
            .O(N__32745),
            .I(N__32712));
    InMux I__7562 (
            .O(N__32744),
            .I(N__32709));
    Span4Mux_s3_h I__7561 (
            .O(N__32741),
            .I(N__32706));
    InMux I__7560 (
            .O(N__32740),
            .I(N__32703));
    LocalMux I__7559 (
            .O(N__32737),
            .I(N__32698));
    Span4Mux_s3_h I__7558 (
            .O(N__32732),
            .I(N__32698));
    Span4Mux_v I__7557 (
            .O(N__32727),
            .I(N__32691));
    LocalMux I__7556 (
            .O(N__32724),
            .I(N__32691));
    Span4Mux_v I__7555 (
            .O(N__32715),
            .I(N__32691));
    LocalMux I__7554 (
            .O(N__32712),
            .I(\POWERLED.N_430 ));
    LocalMux I__7553 (
            .O(N__32709),
            .I(\POWERLED.N_430 ));
    Odrv4 I__7552 (
            .O(N__32706),
            .I(\POWERLED.N_430 ));
    LocalMux I__7551 (
            .O(N__32703),
            .I(\POWERLED.N_430 ));
    Odrv4 I__7550 (
            .O(N__32698),
            .I(\POWERLED.N_430 ));
    Odrv4 I__7549 (
            .O(N__32691),
            .I(\POWERLED.N_430 ));
    CascadeMux I__7548 (
            .O(N__32678),
            .I(\POWERLED.un1_clk_100khz_51_and_i_3_cascade_ ));
    InMux I__7547 (
            .O(N__32675),
            .I(N__32664));
    IoInMux I__7546 (
            .O(N__32674),
            .I(N__32661));
    InMux I__7545 (
            .O(N__32673),
            .I(N__32656));
    InMux I__7544 (
            .O(N__32672),
            .I(N__32656));
    InMux I__7543 (
            .O(N__32671),
            .I(N__32653));
    InMux I__7542 (
            .O(N__32670),
            .I(N__32650));
    InMux I__7541 (
            .O(N__32669),
            .I(N__32647));
    CascadeMux I__7540 (
            .O(N__32668),
            .I(N__32641));
    CascadeMux I__7539 (
            .O(N__32667),
            .I(N__32634));
    LocalMux I__7538 (
            .O(N__32664),
            .I(N__32631));
    LocalMux I__7537 (
            .O(N__32661),
            .I(N__32621));
    LocalMux I__7536 (
            .O(N__32656),
            .I(N__32621));
    LocalMux I__7535 (
            .O(N__32653),
            .I(N__32614));
    LocalMux I__7534 (
            .O(N__32650),
            .I(N__32614));
    LocalMux I__7533 (
            .O(N__32647),
            .I(N__32614));
    InMux I__7532 (
            .O(N__32646),
            .I(N__32611));
    InMux I__7531 (
            .O(N__32645),
            .I(N__32608));
    InMux I__7530 (
            .O(N__32644),
            .I(N__32604));
    InMux I__7529 (
            .O(N__32641),
            .I(N__32601));
    InMux I__7528 (
            .O(N__32640),
            .I(N__32594));
    InMux I__7527 (
            .O(N__32639),
            .I(N__32594));
    InMux I__7526 (
            .O(N__32638),
            .I(N__32594));
    InMux I__7525 (
            .O(N__32637),
            .I(N__32590));
    InMux I__7524 (
            .O(N__32634),
            .I(N__32587));
    Span4Mux_v I__7523 (
            .O(N__32631),
            .I(N__32584));
    InMux I__7522 (
            .O(N__32630),
            .I(N__32579));
    InMux I__7521 (
            .O(N__32629),
            .I(N__32579));
    CascadeMux I__7520 (
            .O(N__32628),
            .I(N__32576));
    InMux I__7519 (
            .O(N__32627),
            .I(N__32570));
    InMux I__7518 (
            .O(N__32626),
            .I(N__32570));
    Span4Mux_s3_v I__7517 (
            .O(N__32621),
            .I(N__32567));
    Span4Mux_s3_v I__7516 (
            .O(N__32614),
            .I(N__32562));
    LocalMux I__7515 (
            .O(N__32611),
            .I(N__32562));
    LocalMux I__7514 (
            .O(N__32608),
            .I(N__32559));
    InMux I__7513 (
            .O(N__32607),
            .I(N__32556));
    LocalMux I__7512 (
            .O(N__32604),
            .I(N__32553));
    LocalMux I__7511 (
            .O(N__32601),
            .I(N__32548));
    LocalMux I__7510 (
            .O(N__32594),
            .I(N__32548));
    InMux I__7509 (
            .O(N__32593),
            .I(N__32545));
    LocalMux I__7508 (
            .O(N__32590),
            .I(N__32542));
    LocalMux I__7507 (
            .O(N__32587),
            .I(N__32539));
    Span4Mux_h I__7506 (
            .O(N__32584),
            .I(N__32534));
    LocalMux I__7505 (
            .O(N__32579),
            .I(N__32534));
    InMux I__7504 (
            .O(N__32576),
            .I(N__32529));
    InMux I__7503 (
            .O(N__32575),
            .I(N__32529));
    LocalMux I__7502 (
            .O(N__32570),
            .I(N__32522));
    Span4Mux_v I__7501 (
            .O(N__32567),
            .I(N__32522));
    Span4Mux_v I__7500 (
            .O(N__32562),
            .I(N__32522));
    Span4Mux_s3_h I__7499 (
            .O(N__32559),
            .I(N__32515));
    LocalMux I__7498 (
            .O(N__32556),
            .I(N__32515));
    Span4Mux_s3_h I__7497 (
            .O(N__32553),
            .I(N__32515));
    Span4Mux_s3_h I__7496 (
            .O(N__32548),
            .I(N__32510));
    LocalMux I__7495 (
            .O(N__32545),
            .I(N__32510));
    Span4Mux_s3_h I__7494 (
            .O(N__32542),
            .I(N__32507));
    Odrv4 I__7493 (
            .O(N__32539),
            .I(G_141));
    Odrv4 I__7492 (
            .O(N__32534),
            .I(G_141));
    LocalMux I__7491 (
            .O(N__32529),
            .I(G_141));
    Odrv4 I__7490 (
            .O(N__32522),
            .I(G_141));
    Odrv4 I__7489 (
            .O(N__32515),
            .I(G_141));
    Odrv4 I__7488 (
            .O(N__32510),
            .I(G_141));
    Odrv4 I__7487 (
            .O(N__32507),
            .I(G_141));
    CascadeMux I__7486 (
            .O(N__32492),
            .I(N__32489));
    InMux I__7485 (
            .O(N__32489),
            .I(N__32483));
    InMux I__7484 (
            .O(N__32488),
            .I(N__32483));
    LocalMux I__7483 (
            .O(N__32483),
            .I(\POWERLED.dutycycle_RNI0DF58Z0Z_5 ));
    ClkMux I__7482 (
            .O(N__32480),
            .I(N__32476));
    ClkMux I__7481 (
            .O(N__32479),
            .I(N__32473));
    LocalMux I__7480 (
            .O(N__32476),
            .I(N__32454));
    LocalMux I__7479 (
            .O(N__32473),
            .I(N__32454));
    ClkMux I__7478 (
            .O(N__32472),
            .I(N__32451));
    ClkMux I__7477 (
            .O(N__32471),
            .I(N__32446));
    ClkMux I__7476 (
            .O(N__32470),
            .I(N__32443));
    ClkMux I__7475 (
            .O(N__32469),
            .I(N__32440));
    ClkMux I__7474 (
            .O(N__32468),
            .I(N__32437));
    ClkMux I__7473 (
            .O(N__32467),
            .I(N__32432));
    ClkMux I__7472 (
            .O(N__32466),
            .I(N__32427));
    ClkMux I__7471 (
            .O(N__32465),
            .I(N__32424));
    ClkMux I__7470 (
            .O(N__32464),
            .I(N__32420));
    ClkMux I__7469 (
            .O(N__32463),
            .I(N__32416));
    ClkMux I__7468 (
            .O(N__32462),
            .I(N__32413));
    ClkMux I__7467 (
            .O(N__32461),
            .I(N__32408));
    ClkMux I__7466 (
            .O(N__32460),
            .I(N__32403));
    ClkMux I__7465 (
            .O(N__32459),
            .I(N__32398));
    Span4Mux_s1_v I__7464 (
            .O(N__32454),
            .I(N__32392));
    LocalMux I__7463 (
            .O(N__32451),
            .I(N__32392));
    ClkMux I__7462 (
            .O(N__32450),
            .I(N__32389));
    ClkMux I__7461 (
            .O(N__32449),
            .I(N__32386));
    LocalMux I__7460 (
            .O(N__32446),
            .I(N__32381));
    LocalMux I__7459 (
            .O(N__32443),
            .I(N__32377));
    LocalMux I__7458 (
            .O(N__32440),
            .I(N__32372));
    LocalMux I__7457 (
            .O(N__32437),
            .I(N__32372));
    ClkMux I__7456 (
            .O(N__32436),
            .I(N__32369));
    ClkMux I__7455 (
            .O(N__32435),
            .I(N__32366));
    LocalMux I__7454 (
            .O(N__32432),
            .I(N__32363));
    ClkMux I__7453 (
            .O(N__32431),
            .I(N__32360));
    ClkMux I__7452 (
            .O(N__32430),
            .I(N__32357));
    LocalMux I__7451 (
            .O(N__32427),
            .I(N__32351));
    LocalMux I__7450 (
            .O(N__32424),
            .I(N__32346));
    ClkMux I__7449 (
            .O(N__32423),
            .I(N__32343));
    LocalMux I__7448 (
            .O(N__32420),
            .I(N__32339));
    ClkMux I__7447 (
            .O(N__32419),
            .I(N__32336));
    LocalMux I__7446 (
            .O(N__32416),
            .I(N__32329));
    LocalMux I__7445 (
            .O(N__32413),
            .I(N__32326));
    ClkMux I__7444 (
            .O(N__32412),
            .I(N__32323));
    ClkMux I__7443 (
            .O(N__32411),
            .I(N__32319));
    LocalMux I__7442 (
            .O(N__32408),
            .I(N__32313));
    ClkMux I__7441 (
            .O(N__32407),
            .I(N__32310));
    ClkMux I__7440 (
            .O(N__32406),
            .I(N__32306));
    LocalMux I__7439 (
            .O(N__32403),
            .I(N__32303));
    ClkMux I__7438 (
            .O(N__32402),
            .I(N__32300));
    ClkMux I__7437 (
            .O(N__32401),
            .I(N__32296));
    LocalMux I__7436 (
            .O(N__32398),
            .I(N__32293));
    ClkMux I__7435 (
            .O(N__32397),
            .I(N__32290));
    Span4Mux_v I__7434 (
            .O(N__32392),
            .I(N__32285));
    LocalMux I__7433 (
            .O(N__32389),
            .I(N__32285));
    LocalMux I__7432 (
            .O(N__32386),
            .I(N__32276));
    ClkMux I__7431 (
            .O(N__32385),
            .I(N__32273));
    ClkMux I__7430 (
            .O(N__32384),
            .I(N__32270));
    Span4Mux_v I__7429 (
            .O(N__32381),
            .I(N__32266));
    ClkMux I__7428 (
            .O(N__32380),
            .I(N__32262));
    Span4Mux_v I__7427 (
            .O(N__32377),
            .I(N__32252));
    Span4Mux_v I__7426 (
            .O(N__32372),
            .I(N__32252));
    LocalMux I__7425 (
            .O(N__32369),
            .I(N__32252));
    LocalMux I__7424 (
            .O(N__32366),
            .I(N__32252));
    Span4Mux_v I__7423 (
            .O(N__32363),
            .I(N__32245));
    LocalMux I__7422 (
            .O(N__32360),
            .I(N__32245));
    LocalMux I__7421 (
            .O(N__32357),
            .I(N__32245));
    ClkMux I__7420 (
            .O(N__32356),
            .I(N__32242));
    ClkMux I__7419 (
            .O(N__32355),
            .I(N__32239));
    ClkMux I__7418 (
            .O(N__32354),
            .I(N__32236));
    Span4Mux_h I__7417 (
            .O(N__32351),
            .I(N__32232));
    ClkMux I__7416 (
            .O(N__32350),
            .I(N__32229));
    ClkMux I__7415 (
            .O(N__32349),
            .I(N__32221));
    Span4Mux_s1_h I__7414 (
            .O(N__32346),
            .I(N__32215));
    LocalMux I__7413 (
            .O(N__32343),
            .I(N__32215));
    ClkMux I__7412 (
            .O(N__32342),
            .I(N__32212));
    Span4Mux_s1_h I__7411 (
            .O(N__32339),
            .I(N__32207));
    LocalMux I__7410 (
            .O(N__32336),
            .I(N__32207));
    ClkMux I__7409 (
            .O(N__32335),
            .I(N__32202));
    ClkMux I__7408 (
            .O(N__32334),
            .I(N__32198));
    ClkMux I__7407 (
            .O(N__32333),
            .I(N__32195));
    ClkMux I__7406 (
            .O(N__32332),
            .I(N__32192));
    Span4Mux_h I__7405 (
            .O(N__32329),
            .I(N__32189));
    Span4Mux_s1_h I__7404 (
            .O(N__32326),
            .I(N__32184));
    LocalMux I__7403 (
            .O(N__32323),
            .I(N__32184));
    ClkMux I__7402 (
            .O(N__32322),
            .I(N__32181));
    LocalMux I__7401 (
            .O(N__32319),
            .I(N__32176));
    ClkMux I__7400 (
            .O(N__32318),
            .I(N__32173));
    ClkMux I__7399 (
            .O(N__32317),
            .I(N__32170));
    ClkMux I__7398 (
            .O(N__32316),
            .I(N__32167));
    Span4Mux_v I__7397 (
            .O(N__32313),
            .I(N__32161));
    LocalMux I__7396 (
            .O(N__32310),
            .I(N__32161));
    ClkMux I__7395 (
            .O(N__32309),
            .I(N__32158));
    LocalMux I__7394 (
            .O(N__32306),
            .I(N__32155));
    Span4Mux_v I__7393 (
            .O(N__32303),
            .I(N__32150));
    LocalMux I__7392 (
            .O(N__32300),
            .I(N__32150));
    ClkMux I__7391 (
            .O(N__32299),
            .I(N__32147));
    LocalMux I__7390 (
            .O(N__32296),
            .I(N__32144));
    Span4Mux_h I__7389 (
            .O(N__32293),
            .I(N__32139));
    LocalMux I__7388 (
            .O(N__32290),
            .I(N__32139));
    Span4Mux_v I__7387 (
            .O(N__32285),
            .I(N__32136));
    ClkMux I__7386 (
            .O(N__32284),
            .I(N__32133));
    ClkMux I__7385 (
            .O(N__32283),
            .I(N__32130));
    ClkMux I__7384 (
            .O(N__32282),
            .I(N__32127));
    ClkMux I__7383 (
            .O(N__32281),
            .I(N__32123));
    ClkMux I__7382 (
            .O(N__32280),
            .I(N__32120));
    ClkMux I__7381 (
            .O(N__32279),
            .I(N__32117));
    Span4Mux_v I__7380 (
            .O(N__32276),
            .I(N__32112));
    LocalMux I__7379 (
            .O(N__32273),
            .I(N__32112));
    LocalMux I__7378 (
            .O(N__32270),
            .I(N__32109));
    ClkMux I__7377 (
            .O(N__32269),
            .I(N__32106));
    Span4Mux_s0_v I__7376 (
            .O(N__32266),
            .I(N__32103));
    ClkMux I__7375 (
            .O(N__32265),
            .I(N__32100));
    LocalMux I__7374 (
            .O(N__32262),
            .I(N__32097));
    ClkMux I__7373 (
            .O(N__32261),
            .I(N__32094));
    Span4Mux_v I__7372 (
            .O(N__32252),
            .I(N__32083));
    Span4Mux_v I__7371 (
            .O(N__32245),
            .I(N__32083));
    LocalMux I__7370 (
            .O(N__32242),
            .I(N__32083));
    LocalMux I__7369 (
            .O(N__32239),
            .I(N__32083));
    LocalMux I__7368 (
            .O(N__32236),
            .I(N__32083));
    ClkMux I__7367 (
            .O(N__32235),
            .I(N__32080));
    Span4Mux_v I__7366 (
            .O(N__32232),
            .I(N__32075));
    LocalMux I__7365 (
            .O(N__32229),
            .I(N__32075));
    ClkMux I__7364 (
            .O(N__32228),
            .I(N__32072));
    ClkMux I__7363 (
            .O(N__32227),
            .I(N__32069));
    ClkMux I__7362 (
            .O(N__32226),
            .I(N__32066));
    ClkMux I__7361 (
            .O(N__32225),
            .I(N__32063));
    ClkMux I__7360 (
            .O(N__32224),
            .I(N__32060));
    LocalMux I__7359 (
            .O(N__32221),
            .I(N__32057));
    ClkMux I__7358 (
            .O(N__32220),
            .I(N__32054));
    Span4Mux_v I__7357 (
            .O(N__32215),
            .I(N__32047));
    LocalMux I__7356 (
            .O(N__32212),
            .I(N__32047));
    Span4Mux_h I__7355 (
            .O(N__32207),
            .I(N__32042));
    ClkMux I__7354 (
            .O(N__32206),
            .I(N__32039));
    ClkMux I__7353 (
            .O(N__32205),
            .I(N__32036));
    LocalMux I__7352 (
            .O(N__32202),
            .I(N__32033));
    ClkMux I__7351 (
            .O(N__32201),
            .I(N__32030));
    LocalMux I__7350 (
            .O(N__32198),
            .I(N__32025));
    LocalMux I__7349 (
            .O(N__32195),
            .I(N__32025));
    LocalMux I__7348 (
            .O(N__32192),
            .I(N__32022));
    Span4Mux_v I__7347 (
            .O(N__32189),
            .I(N__32017));
    Span4Mux_h I__7346 (
            .O(N__32184),
            .I(N__32017));
    LocalMux I__7345 (
            .O(N__32181),
            .I(N__32014));
    ClkMux I__7344 (
            .O(N__32180),
            .I(N__32011));
    ClkMux I__7343 (
            .O(N__32179),
            .I(N__32008));
    Span4Mux_s2_h I__7342 (
            .O(N__32176),
            .I(N__32003));
    LocalMux I__7341 (
            .O(N__32173),
            .I(N__32003));
    LocalMux I__7340 (
            .O(N__32170),
            .I(N__32000));
    LocalMux I__7339 (
            .O(N__32167),
            .I(N__31997));
    ClkMux I__7338 (
            .O(N__32166),
            .I(N__31994));
    Span4Mux_v I__7337 (
            .O(N__32161),
            .I(N__31991));
    LocalMux I__7336 (
            .O(N__32158),
            .I(N__31988));
    Span4Mux_v I__7335 (
            .O(N__32155),
            .I(N__31981));
    Span4Mux_h I__7334 (
            .O(N__32150),
            .I(N__31981));
    LocalMux I__7333 (
            .O(N__32147),
            .I(N__31981));
    Span4Mux_h I__7332 (
            .O(N__32144),
            .I(N__31968));
    Span4Mux_v I__7331 (
            .O(N__32139),
            .I(N__31968));
    Span4Mux_h I__7330 (
            .O(N__32136),
            .I(N__31968));
    LocalMux I__7329 (
            .O(N__32133),
            .I(N__31968));
    LocalMux I__7328 (
            .O(N__32130),
            .I(N__31968));
    LocalMux I__7327 (
            .O(N__32127),
            .I(N__31968));
    ClkMux I__7326 (
            .O(N__32126),
            .I(N__31965));
    LocalMux I__7325 (
            .O(N__32123),
            .I(N__31958));
    LocalMux I__7324 (
            .O(N__32120),
            .I(N__31958));
    LocalMux I__7323 (
            .O(N__32117),
            .I(N__31958));
    Span4Mux_v I__7322 (
            .O(N__32112),
            .I(N__31947));
    Span4Mux_v I__7321 (
            .O(N__32109),
            .I(N__31947));
    LocalMux I__7320 (
            .O(N__32106),
            .I(N__31947));
    Span4Mux_h I__7319 (
            .O(N__32103),
            .I(N__31947));
    LocalMux I__7318 (
            .O(N__32100),
            .I(N__31947));
    IoSpan4Mux I__7317 (
            .O(N__32097),
            .I(N__31944));
    LocalMux I__7316 (
            .O(N__32094),
            .I(N__31941));
    Span4Mux_v I__7315 (
            .O(N__32083),
            .I(N__31936));
    LocalMux I__7314 (
            .O(N__32080),
            .I(N__31936));
    Span4Mux_v I__7313 (
            .O(N__32075),
            .I(N__31925));
    LocalMux I__7312 (
            .O(N__32072),
            .I(N__31925));
    LocalMux I__7311 (
            .O(N__32069),
            .I(N__31925));
    LocalMux I__7310 (
            .O(N__32066),
            .I(N__31925));
    LocalMux I__7309 (
            .O(N__32063),
            .I(N__31925));
    LocalMux I__7308 (
            .O(N__32060),
            .I(N__31918));
    Span4Mux_h I__7307 (
            .O(N__32057),
            .I(N__31918));
    LocalMux I__7306 (
            .O(N__32054),
            .I(N__31918));
    ClkMux I__7305 (
            .O(N__32053),
            .I(N__31915));
    ClkMux I__7304 (
            .O(N__32052),
            .I(N__31912));
    Span4Mux_v I__7303 (
            .O(N__32047),
            .I(N__31909));
    ClkMux I__7302 (
            .O(N__32046),
            .I(N__31906));
    ClkMux I__7301 (
            .O(N__32045),
            .I(N__31903));
    Span4Mux_v I__7300 (
            .O(N__32042),
            .I(N__31896));
    LocalMux I__7299 (
            .O(N__32039),
            .I(N__31896));
    LocalMux I__7298 (
            .O(N__32036),
            .I(N__31896));
    Span4Mux_s2_h I__7297 (
            .O(N__32033),
            .I(N__31891));
    LocalMux I__7296 (
            .O(N__32030),
            .I(N__31891));
    Span4Mux_v I__7295 (
            .O(N__32025),
            .I(N__31886));
    Span4Mux_s1_h I__7294 (
            .O(N__32022),
            .I(N__31886));
    Span4Mux_v I__7293 (
            .O(N__32017),
            .I(N__31877));
    Span4Mux_v I__7292 (
            .O(N__32014),
            .I(N__31877));
    LocalMux I__7291 (
            .O(N__32011),
            .I(N__31877));
    LocalMux I__7290 (
            .O(N__32008),
            .I(N__31877));
    Span4Mux_v I__7289 (
            .O(N__32003),
            .I(N__31868));
    Span4Mux_s2_h I__7288 (
            .O(N__32000),
            .I(N__31868));
    Span4Mux_s2_h I__7287 (
            .O(N__31997),
            .I(N__31868));
    LocalMux I__7286 (
            .O(N__31994),
            .I(N__31868));
    IoSpan4Mux I__7285 (
            .O(N__31991),
            .I(N__31863));
    IoSpan4Mux I__7284 (
            .O(N__31988),
            .I(N__31863));
    Span4Mux_v I__7283 (
            .O(N__31981),
            .I(N__31856));
    Span4Mux_v I__7282 (
            .O(N__31968),
            .I(N__31856));
    LocalMux I__7281 (
            .O(N__31965),
            .I(N__31856));
    Span4Mux_v I__7280 (
            .O(N__31958),
            .I(N__31851));
    Span4Mux_v I__7279 (
            .O(N__31947),
            .I(N__31851));
    IoSpan4Mux I__7278 (
            .O(N__31944),
            .I(N__31846));
    IoSpan4Mux I__7277 (
            .O(N__31941),
            .I(N__31846));
    Span4Mux_h I__7276 (
            .O(N__31936),
            .I(N__31837));
    Span4Mux_v I__7275 (
            .O(N__31925),
            .I(N__31837));
    Span4Mux_v I__7274 (
            .O(N__31918),
            .I(N__31837));
    LocalMux I__7273 (
            .O(N__31915),
            .I(N__31837));
    LocalMux I__7272 (
            .O(N__31912),
            .I(N__31833));
    Span4Mux_h I__7271 (
            .O(N__31909),
            .I(N__31826));
    LocalMux I__7270 (
            .O(N__31906),
            .I(N__31826));
    LocalMux I__7269 (
            .O(N__31903),
            .I(N__31826));
    Span4Mux_v I__7268 (
            .O(N__31896),
            .I(N__31821));
    Span4Mux_h I__7267 (
            .O(N__31891),
            .I(N__31821));
    Span4Mux_h I__7266 (
            .O(N__31886),
            .I(N__31814));
    Span4Mux_v I__7265 (
            .O(N__31877),
            .I(N__31814));
    Span4Mux_h I__7264 (
            .O(N__31868),
            .I(N__31814));
    IoSpan4Mux I__7263 (
            .O(N__31863),
            .I(N__31807));
    IoSpan4Mux I__7262 (
            .O(N__31856),
            .I(N__31807));
    IoSpan4Mux I__7261 (
            .O(N__31851),
            .I(N__31807));
    IoSpan4Mux I__7260 (
            .O(N__31846),
            .I(N__31802));
    IoSpan4Mux I__7259 (
            .O(N__31837),
            .I(N__31802));
    ClkMux I__7258 (
            .O(N__31836),
            .I(N__31799));
    Sp12to4 I__7257 (
            .O(N__31833),
            .I(N__31794));
    Sp12to4 I__7256 (
            .O(N__31826),
            .I(N__31794));
    Odrv4 I__7255 (
            .O(N__31821),
            .I(fpga_osc));
    Odrv4 I__7254 (
            .O(N__31814),
            .I(fpga_osc));
    Odrv4 I__7253 (
            .O(N__31807),
            .I(fpga_osc));
    Odrv4 I__7252 (
            .O(N__31802),
            .I(fpga_osc));
    LocalMux I__7251 (
            .O(N__31799),
            .I(fpga_osc));
    Odrv12 I__7250 (
            .O(N__31794),
            .I(fpga_osc));
    SRMux I__7249 (
            .O(N__31781),
            .I(N__31777));
    SRMux I__7248 (
            .O(N__31780),
            .I(N__31774));
    LocalMux I__7247 (
            .O(N__31777),
            .I(N__31768));
    LocalMux I__7246 (
            .O(N__31774),
            .I(N__31764));
    SRMux I__7245 (
            .O(N__31773),
            .I(N__31761));
    SRMux I__7244 (
            .O(N__31772),
            .I(N__31758));
    SRMux I__7243 (
            .O(N__31771),
            .I(N__31751));
    Span4Mux_h I__7242 (
            .O(N__31768),
            .I(N__31747));
    SRMux I__7241 (
            .O(N__31767),
            .I(N__31744));
    Span4Mux_h I__7240 (
            .O(N__31764),
            .I(N__31741));
    LocalMux I__7239 (
            .O(N__31761),
            .I(N__31738));
    LocalMux I__7238 (
            .O(N__31758),
            .I(N__31735));
    SRMux I__7237 (
            .O(N__31757),
            .I(N__31732));
    SRMux I__7236 (
            .O(N__31756),
            .I(N__31728));
    SRMux I__7235 (
            .O(N__31755),
            .I(N__31725));
    SRMux I__7234 (
            .O(N__31754),
            .I(N__31722));
    LocalMux I__7233 (
            .O(N__31751),
            .I(N__31718));
    SRMux I__7232 (
            .O(N__31750),
            .I(N__31715));
    Span4Mux_s1_v I__7231 (
            .O(N__31747),
            .I(N__31710));
    LocalMux I__7230 (
            .O(N__31744),
            .I(N__31710));
    Span4Mux_s0_v I__7229 (
            .O(N__31741),
            .I(N__31707));
    Span4Mux_s1_h I__7228 (
            .O(N__31738),
            .I(N__31700));
    Span4Mux_v I__7227 (
            .O(N__31735),
            .I(N__31700));
    LocalMux I__7226 (
            .O(N__31732),
            .I(N__31700));
    SRMux I__7225 (
            .O(N__31731),
            .I(N__31697));
    LocalMux I__7224 (
            .O(N__31728),
            .I(N__31694));
    LocalMux I__7223 (
            .O(N__31725),
            .I(N__31691));
    LocalMux I__7222 (
            .O(N__31722),
            .I(N__31688));
    SRMux I__7221 (
            .O(N__31721),
            .I(N__31685));
    Span4Mux_h I__7220 (
            .O(N__31718),
            .I(N__31680));
    LocalMux I__7219 (
            .O(N__31715),
            .I(N__31680));
    Span4Mux_v I__7218 (
            .O(N__31710),
            .I(N__31677));
    Span4Mux_v I__7217 (
            .O(N__31707),
            .I(N__31672));
    Span4Mux_h I__7216 (
            .O(N__31700),
            .I(N__31672));
    LocalMux I__7215 (
            .O(N__31697),
            .I(N__31669));
    Span4Mux_s0_h I__7214 (
            .O(N__31694),
            .I(N__31664));
    Span4Mux_v I__7213 (
            .O(N__31691),
            .I(N__31664));
    Span4Mux_v I__7212 (
            .O(N__31688),
            .I(N__31657));
    LocalMux I__7211 (
            .O(N__31685),
            .I(N__31657));
    Span4Mux_s3_v I__7210 (
            .O(N__31680),
            .I(N__31657));
    Span4Mux_v I__7209 (
            .O(N__31677),
            .I(N__31654));
    Span4Mux_v I__7208 (
            .O(N__31672),
            .I(N__31651));
    Span4Mux_v I__7207 (
            .O(N__31669),
            .I(N__31644));
    Span4Mux_h I__7206 (
            .O(N__31664),
            .I(N__31644));
    Span4Mux_v I__7205 (
            .O(N__31657),
            .I(N__31644));
    Odrv4 I__7204 (
            .O(N__31654),
            .I(\POWERLED.N_430_iZ0 ));
    Odrv4 I__7203 (
            .O(N__31651),
            .I(\POWERLED.N_430_iZ0 ));
    Odrv4 I__7202 (
            .O(N__31644),
            .I(\POWERLED.N_430_iZ0 ));
    CascadeMux I__7201 (
            .O(N__31637),
            .I(N__31634));
    InMux I__7200 (
            .O(N__31634),
            .I(N__31630));
    InMux I__7199 (
            .O(N__31633),
            .I(N__31627));
    LocalMux I__7198 (
            .O(N__31630),
            .I(\POWERLED.dutycycle_en_8 ));
    LocalMux I__7197 (
            .O(N__31627),
            .I(\POWERLED.dutycycle_en_8 ));
    InMux I__7196 (
            .O(N__31622),
            .I(N__31618));
    InMux I__7195 (
            .O(N__31621),
            .I(N__31615));
    LocalMux I__7194 (
            .O(N__31618),
            .I(N__31610));
    LocalMux I__7193 (
            .O(N__31615),
            .I(N__31610));
    Span4Mux_v I__7192 (
            .O(N__31610),
            .I(N__31607));
    Odrv4 I__7191 (
            .O(N__31607),
            .I(\POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ));
    CascadeMux I__7190 (
            .O(N__31604),
            .I(N__31600));
    InMux I__7189 (
            .O(N__31603),
            .I(N__31595));
    InMux I__7188 (
            .O(N__31600),
            .I(N__31595));
    LocalMux I__7187 (
            .O(N__31595),
            .I(\POWERLED.dutycycleZ1Z_3 ));
    CascadeMux I__7186 (
            .O(N__31592),
            .I(N__31576));
    InMux I__7185 (
            .O(N__31591),
            .I(N__31572));
    InMux I__7184 (
            .O(N__31590),
            .I(N__31569));
    InMux I__7183 (
            .O(N__31589),
            .I(N__31560));
    InMux I__7182 (
            .O(N__31588),
            .I(N__31557));
    InMux I__7181 (
            .O(N__31587),
            .I(N__31554));
    InMux I__7180 (
            .O(N__31586),
            .I(N__31545));
    InMux I__7179 (
            .O(N__31585),
            .I(N__31545));
    InMux I__7178 (
            .O(N__31584),
            .I(N__31545));
    InMux I__7177 (
            .O(N__31583),
            .I(N__31545));
    InMux I__7176 (
            .O(N__31582),
            .I(N__31540));
    InMux I__7175 (
            .O(N__31581),
            .I(N__31540));
    InMux I__7174 (
            .O(N__31580),
            .I(N__31535));
    InMux I__7173 (
            .O(N__31579),
            .I(N__31535));
    InMux I__7172 (
            .O(N__31576),
            .I(N__31530));
    InMux I__7171 (
            .O(N__31575),
            .I(N__31530));
    LocalMux I__7170 (
            .O(N__31572),
            .I(N__31527));
    LocalMux I__7169 (
            .O(N__31569),
            .I(N__31524));
    InMux I__7168 (
            .O(N__31568),
            .I(N__31515));
    InMux I__7167 (
            .O(N__31567),
            .I(N__31515));
    InMux I__7166 (
            .O(N__31566),
            .I(N__31515));
    InMux I__7165 (
            .O(N__31565),
            .I(N__31515));
    InMux I__7164 (
            .O(N__31564),
            .I(N__31512));
    CascadeMux I__7163 (
            .O(N__31563),
            .I(N__31509));
    LocalMux I__7162 (
            .O(N__31560),
            .I(N__31505));
    LocalMux I__7161 (
            .O(N__31557),
            .I(N__31502));
    LocalMux I__7160 (
            .O(N__31554),
            .I(N__31499));
    LocalMux I__7159 (
            .O(N__31545),
            .I(N__31488));
    LocalMux I__7158 (
            .O(N__31540),
            .I(N__31488));
    LocalMux I__7157 (
            .O(N__31535),
            .I(N__31488));
    LocalMux I__7156 (
            .O(N__31530),
            .I(N__31488));
    Span4Mux_s3_h I__7155 (
            .O(N__31527),
            .I(N__31479));
    Span4Mux_v I__7154 (
            .O(N__31524),
            .I(N__31479));
    LocalMux I__7153 (
            .O(N__31515),
            .I(N__31479));
    LocalMux I__7152 (
            .O(N__31512),
            .I(N__31479));
    InMux I__7151 (
            .O(N__31509),
            .I(N__31474));
    InMux I__7150 (
            .O(N__31508),
            .I(N__31474));
    Span12Mux_s10_h I__7149 (
            .O(N__31505),
            .I(N__31471));
    Span4Mux_v I__7148 (
            .O(N__31502),
            .I(N__31468));
    Span4Mux_v I__7147 (
            .O(N__31499),
            .I(N__31465));
    InMux I__7146 (
            .O(N__31498),
            .I(N__31460));
    InMux I__7145 (
            .O(N__31497),
            .I(N__31460));
    Span4Mux_s3_v I__7144 (
            .O(N__31488),
            .I(N__31453));
    Span4Mux_v I__7143 (
            .O(N__31479),
            .I(N__31453));
    LocalMux I__7142 (
            .O(N__31474),
            .I(N__31453));
    Odrv12 I__7141 (
            .O(N__31471),
            .I(\POWERLED.N_421 ));
    Odrv4 I__7140 (
            .O(N__31468),
            .I(\POWERLED.N_421 ));
    Odrv4 I__7139 (
            .O(N__31465),
            .I(\POWERLED.N_421 ));
    LocalMux I__7138 (
            .O(N__31460),
            .I(\POWERLED.N_421 ));
    Odrv4 I__7137 (
            .O(N__31453),
            .I(\POWERLED.N_421 ));
    CascadeMux I__7136 (
            .O(N__31442),
            .I(\POWERLED.dutycycleZ0Z_8_cascade_ ));
    CascadeMux I__7135 (
            .O(N__31439),
            .I(\POWERLED.un1_dutycycle_53_axb_3_1_cascade_ ));
    CascadeMux I__7134 (
            .O(N__31436),
            .I(N__31427));
    InMux I__7133 (
            .O(N__31435),
            .I(N__31418));
    InMux I__7132 (
            .O(N__31434),
            .I(N__31413));
    InMux I__7131 (
            .O(N__31433),
            .I(N__31413));
    InMux I__7130 (
            .O(N__31432),
            .I(N__31410));
    InMux I__7129 (
            .O(N__31431),
            .I(N__31407));
    CascadeMux I__7128 (
            .O(N__31430),
            .I(N__31402));
    InMux I__7127 (
            .O(N__31427),
            .I(N__31395));
    InMux I__7126 (
            .O(N__31426),
            .I(N__31392));
    InMux I__7125 (
            .O(N__31425),
            .I(N__31385));
    InMux I__7124 (
            .O(N__31424),
            .I(N__31385));
    InMux I__7123 (
            .O(N__31423),
            .I(N__31385));
    InMux I__7122 (
            .O(N__31422),
            .I(N__31380));
    InMux I__7121 (
            .O(N__31421),
            .I(N__31380));
    LocalMux I__7120 (
            .O(N__31418),
            .I(N__31377));
    LocalMux I__7119 (
            .O(N__31413),
            .I(N__31374));
    LocalMux I__7118 (
            .O(N__31410),
            .I(N__31369));
    LocalMux I__7117 (
            .O(N__31407),
            .I(N__31369));
    InMux I__7116 (
            .O(N__31406),
            .I(N__31358));
    InMux I__7115 (
            .O(N__31405),
            .I(N__31358));
    InMux I__7114 (
            .O(N__31402),
            .I(N__31358));
    InMux I__7113 (
            .O(N__31401),
            .I(N__31358));
    InMux I__7112 (
            .O(N__31400),
            .I(N__31358));
    InMux I__7111 (
            .O(N__31399),
            .I(N__31353));
    InMux I__7110 (
            .O(N__31398),
            .I(N__31353));
    LocalMux I__7109 (
            .O(N__31395),
            .I(N__31348));
    LocalMux I__7108 (
            .O(N__31392),
            .I(N__31348));
    LocalMux I__7107 (
            .O(N__31385),
            .I(N__31345));
    LocalMux I__7106 (
            .O(N__31380),
            .I(N__31340));
    Span4Mux_s2_h I__7105 (
            .O(N__31377),
            .I(N__31340));
    Span4Mux_s2_h I__7104 (
            .O(N__31374),
            .I(N__31337));
    Odrv4 I__7103 (
            .O(N__31369),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__7102 (
            .O(N__31358),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__7101 (
            .O(N__31353),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__7100 (
            .O(N__31348),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__7099 (
            .O(N__31345),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__7098 (
            .O(N__31340),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__7097 (
            .O(N__31337),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    CascadeMux I__7096 (
            .O(N__31322),
            .I(N__31318));
    InMux I__7095 (
            .O(N__31321),
            .I(N__31315));
    InMux I__7094 (
            .O(N__31318),
            .I(N__31311));
    LocalMux I__7093 (
            .O(N__31315),
            .I(N__31302));
    InMux I__7092 (
            .O(N__31314),
            .I(N__31299));
    LocalMux I__7091 (
            .O(N__31311),
            .I(N__31294));
    InMux I__7090 (
            .O(N__31310),
            .I(N__31291));
    InMux I__7089 (
            .O(N__31309),
            .I(N__31288));
    InMux I__7088 (
            .O(N__31308),
            .I(N__31285));
    CascadeMux I__7087 (
            .O(N__31307),
            .I(N__31282));
    InMux I__7086 (
            .O(N__31306),
            .I(N__31277));
    InMux I__7085 (
            .O(N__31305),
            .I(N__31277));
    Span4Mux_v I__7084 (
            .O(N__31302),
            .I(N__31273));
    LocalMux I__7083 (
            .O(N__31299),
            .I(N__31270));
    InMux I__7082 (
            .O(N__31298),
            .I(N__31265));
    InMux I__7081 (
            .O(N__31297),
            .I(N__31265));
    Span4Mux_h I__7080 (
            .O(N__31294),
            .I(N__31260));
    LocalMux I__7079 (
            .O(N__31291),
            .I(N__31257));
    LocalMux I__7078 (
            .O(N__31288),
            .I(N__31252));
    LocalMux I__7077 (
            .O(N__31285),
            .I(N__31252));
    InMux I__7076 (
            .O(N__31282),
            .I(N__31249));
    LocalMux I__7075 (
            .O(N__31277),
            .I(N__31244));
    InMux I__7074 (
            .O(N__31276),
            .I(N__31241));
    Span4Mux_h I__7073 (
            .O(N__31273),
            .I(N__31238));
    Span4Mux_v I__7072 (
            .O(N__31270),
            .I(N__31233));
    LocalMux I__7071 (
            .O(N__31265),
            .I(N__31233));
    InMux I__7070 (
            .O(N__31264),
            .I(N__31230));
    InMux I__7069 (
            .O(N__31263),
            .I(N__31227));
    Span4Mux_v I__7068 (
            .O(N__31260),
            .I(N__31222));
    Span4Mux_h I__7067 (
            .O(N__31257),
            .I(N__31222));
    Span4Mux_v I__7066 (
            .O(N__31252),
            .I(N__31217));
    LocalMux I__7065 (
            .O(N__31249),
            .I(N__31217));
    InMux I__7064 (
            .O(N__31248),
            .I(N__31212));
    InMux I__7063 (
            .O(N__31247),
            .I(N__31212));
    Span4Mux_h I__7062 (
            .O(N__31244),
            .I(N__31199));
    LocalMux I__7061 (
            .O(N__31241),
            .I(N__31199));
    Span4Mux_s0_h I__7060 (
            .O(N__31238),
            .I(N__31199));
    Span4Mux_h I__7059 (
            .O(N__31233),
            .I(N__31199));
    LocalMux I__7058 (
            .O(N__31230),
            .I(N__31199));
    LocalMux I__7057 (
            .O(N__31227),
            .I(N__31199));
    Odrv4 I__7056 (
            .O(N__31222),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    Odrv4 I__7055 (
            .O(N__31217),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__7054 (
            .O(N__31212),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    Odrv4 I__7053 (
            .O(N__31199),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    CascadeMux I__7052 (
            .O(N__31190),
            .I(\POWERLED.un1_i3_mux_cascade_ ));
    InMux I__7051 (
            .O(N__31187),
            .I(N__31183));
    CascadeMux I__7050 (
            .O(N__31186),
            .I(N__31180));
    LocalMux I__7049 (
            .O(N__31183),
            .I(N__31177));
    InMux I__7048 (
            .O(N__31180),
            .I(N__31174));
    Odrv12 I__7047 (
            .O(N__31177),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_3 ));
    LocalMux I__7046 (
            .O(N__31174),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_3 ));
    InMux I__7045 (
            .O(N__31169),
            .I(N__31166));
    LocalMux I__7044 (
            .O(N__31166),
            .I(N__31163));
    Span4Mux_h I__7043 (
            .O(N__31163),
            .I(N__31160));
    Span4Mux_h I__7042 (
            .O(N__31160),
            .I(N__31157));
    Odrv4 I__7041 (
            .O(N__31157),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_5 ));
    CascadeMux I__7040 (
            .O(N__31154),
            .I(N__31141));
    InMux I__7039 (
            .O(N__31153),
            .I(N__31133));
    InMux I__7038 (
            .O(N__31152),
            .I(N__31133));
    InMux I__7037 (
            .O(N__31151),
            .I(N__31133));
    InMux I__7036 (
            .O(N__31150),
            .I(N__31128));
    InMux I__7035 (
            .O(N__31149),
            .I(N__31128));
    InMux I__7034 (
            .O(N__31148),
            .I(N__31123));
    InMux I__7033 (
            .O(N__31147),
            .I(N__31123));
    CascadeMux I__7032 (
            .O(N__31146),
            .I(N__31119));
    InMux I__7031 (
            .O(N__31145),
            .I(N__31116));
    InMux I__7030 (
            .O(N__31144),
            .I(N__31109));
    InMux I__7029 (
            .O(N__31141),
            .I(N__31109));
    InMux I__7028 (
            .O(N__31140),
            .I(N__31109));
    LocalMux I__7027 (
            .O(N__31133),
            .I(N__31106));
    LocalMux I__7026 (
            .O(N__31128),
            .I(N__31097));
    LocalMux I__7025 (
            .O(N__31123),
            .I(N__31097));
    InMux I__7024 (
            .O(N__31122),
            .I(N__31094));
    InMux I__7023 (
            .O(N__31119),
            .I(N__31091));
    LocalMux I__7022 (
            .O(N__31116),
            .I(N__31084));
    LocalMux I__7021 (
            .O(N__31109),
            .I(N__31079));
    Span4Mux_s2_v I__7020 (
            .O(N__31106),
            .I(N__31079));
    InMux I__7019 (
            .O(N__31105),
            .I(N__31076));
    InMux I__7018 (
            .O(N__31104),
            .I(N__31069));
    InMux I__7017 (
            .O(N__31103),
            .I(N__31069));
    InMux I__7016 (
            .O(N__31102),
            .I(N__31069));
    Span4Mux_v I__7015 (
            .O(N__31097),
            .I(N__31064));
    LocalMux I__7014 (
            .O(N__31094),
            .I(N__31064));
    LocalMux I__7013 (
            .O(N__31091),
            .I(N__31061));
    InMux I__7012 (
            .O(N__31090),
            .I(N__31056));
    InMux I__7011 (
            .O(N__31089),
            .I(N__31056));
    InMux I__7010 (
            .O(N__31088),
            .I(N__31051));
    InMux I__7009 (
            .O(N__31087),
            .I(N__31051));
    Span4Mux_v I__7008 (
            .O(N__31084),
            .I(N__31046));
    Span4Mux_v I__7007 (
            .O(N__31079),
            .I(N__31046));
    LocalMux I__7006 (
            .O(N__31076),
            .I(N__31039));
    LocalMux I__7005 (
            .O(N__31069),
            .I(N__31039));
    Span4Mux_h I__7004 (
            .O(N__31064),
            .I(N__31039));
    Odrv12 I__7003 (
            .O(N__31061),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__7002 (
            .O(N__31056),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__7001 (
            .O(N__31051),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__7000 (
            .O(N__31046),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__6999 (
            .O(N__31039),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    CascadeMux I__6998 (
            .O(N__31028),
            .I(N__31025));
    InMux I__6997 (
            .O(N__31025),
            .I(N__31015));
    InMux I__6996 (
            .O(N__31024),
            .I(N__31010));
    InMux I__6995 (
            .O(N__31023),
            .I(N__31007));
    CascadeMux I__6994 (
            .O(N__31022),
            .I(N__31004));
    InMux I__6993 (
            .O(N__31021),
            .I(N__30999));
    InMux I__6992 (
            .O(N__31020),
            .I(N__30994));
    InMux I__6991 (
            .O(N__31019),
            .I(N__30994));
    InMux I__6990 (
            .O(N__31018),
            .I(N__30991));
    LocalMux I__6989 (
            .O(N__31015),
            .I(N__30988));
    InMux I__6988 (
            .O(N__31014),
            .I(N__30983));
    InMux I__6987 (
            .O(N__31013),
            .I(N__30983));
    LocalMux I__6986 (
            .O(N__31010),
            .I(N__30978));
    LocalMux I__6985 (
            .O(N__31007),
            .I(N__30975));
    InMux I__6984 (
            .O(N__31004),
            .I(N__30968));
    InMux I__6983 (
            .O(N__31003),
            .I(N__30968));
    InMux I__6982 (
            .O(N__31002),
            .I(N__30968));
    LocalMux I__6981 (
            .O(N__30999),
            .I(N__30963));
    LocalMux I__6980 (
            .O(N__30994),
            .I(N__30963));
    LocalMux I__6979 (
            .O(N__30991),
            .I(N__30960));
    Span12Mux_s4_v I__6978 (
            .O(N__30988),
            .I(N__30955));
    LocalMux I__6977 (
            .O(N__30983),
            .I(N__30955));
    InMux I__6976 (
            .O(N__30982),
            .I(N__30950));
    InMux I__6975 (
            .O(N__30981),
            .I(N__30950));
    Span4Mux_h I__6974 (
            .O(N__30978),
            .I(N__30945));
    Span4Mux_h I__6973 (
            .O(N__30975),
            .I(N__30945));
    LocalMux I__6972 (
            .O(N__30968),
            .I(N__30938));
    Span4Mux_h I__6971 (
            .O(N__30963),
            .I(N__30938));
    Span4Mux_h I__6970 (
            .O(N__30960),
            .I(N__30938));
    Odrv12 I__6969 (
            .O(N__30955),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__6968 (
            .O(N__30950),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__6967 (
            .O(N__30945),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__6966 (
            .O(N__30938),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    InMux I__6965 (
            .O(N__30929),
            .I(N__30921));
    InMux I__6964 (
            .O(N__30928),
            .I(N__30913));
    InMux I__6963 (
            .O(N__30927),
            .I(N__30906));
    InMux I__6962 (
            .O(N__30926),
            .I(N__30906));
    InMux I__6961 (
            .O(N__30925),
            .I(N__30906));
    CascadeMux I__6960 (
            .O(N__30924),
            .I(N__30902));
    LocalMux I__6959 (
            .O(N__30921),
            .I(N__30899));
    CascadeMux I__6958 (
            .O(N__30920),
            .I(N__30896));
    CascadeMux I__6957 (
            .O(N__30919),
            .I(N__30893));
    InMux I__6956 (
            .O(N__30918),
            .I(N__30886));
    InMux I__6955 (
            .O(N__30917),
            .I(N__30886));
    InMux I__6954 (
            .O(N__30916),
            .I(N__30886));
    LocalMux I__6953 (
            .O(N__30913),
            .I(N__30883));
    LocalMux I__6952 (
            .O(N__30906),
            .I(N__30880));
    InMux I__6951 (
            .O(N__30905),
            .I(N__30875));
    InMux I__6950 (
            .O(N__30902),
            .I(N__30875));
    Span12Mux_s6_v I__6949 (
            .O(N__30899),
            .I(N__30872));
    InMux I__6948 (
            .O(N__30896),
            .I(N__30867));
    InMux I__6947 (
            .O(N__30893),
            .I(N__30867));
    LocalMux I__6946 (
            .O(N__30886),
            .I(N__30864));
    Span4Mux_v I__6945 (
            .O(N__30883),
            .I(N__30857));
    Span4Mux_v I__6944 (
            .O(N__30880),
            .I(N__30857));
    LocalMux I__6943 (
            .O(N__30875),
            .I(N__30857));
    Odrv12 I__6942 (
            .O(N__30872),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__6941 (
            .O(N__30867),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__6940 (
            .O(N__30864),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__6939 (
            .O(N__30857),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    InMux I__6938 (
            .O(N__30848),
            .I(N__30845));
    LocalMux I__6937 (
            .O(N__30845),
            .I(\POWERLED.d_i3_mux ));
    CascadeMux I__6936 (
            .O(N__30842),
            .I(\POWERLED.func_state_RNI_5Z0Z_1_cascade_ ));
    InMux I__6935 (
            .O(N__30839),
            .I(N__30836));
    LocalMux I__6934 (
            .O(N__30836),
            .I(N__30832));
    InMux I__6933 (
            .O(N__30835),
            .I(N__30829));
    Odrv4 I__6932 (
            .O(N__30832),
            .I(\POWERLED.N_23_i ));
    LocalMux I__6931 (
            .O(N__30829),
            .I(\POWERLED.N_23_i ));
    InMux I__6930 (
            .O(N__30824),
            .I(N__30821));
    LocalMux I__6929 (
            .O(N__30821),
            .I(N__30818));
    Span4Mux_s2_h I__6928 (
            .O(N__30818),
            .I(N__30815));
    Odrv4 I__6927 (
            .O(N__30815),
            .I(\POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ));
    InMux I__6926 (
            .O(N__30812),
            .I(N__30806));
    InMux I__6925 (
            .O(N__30811),
            .I(N__30806));
    LocalMux I__6924 (
            .O(N__30806),
            .I(\POWERLED.N_85 ));
    InMux I__6923 (
            .O(N__30803),
            .I(N__30800));
    LocalMux I__6922 (
            .O(N__30800),
            .I(N__30796));
    InMux I__6921 (
            .O(N__30799),
            .I(N__30793));
    Odrv4 I__6920 (
            .O(N__30796),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_5 ));
    LocalMux I__6919 (
            .O(N__30793),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_5 ));
    CascadeMux I__6918 (
            .O(N__30788),
            .I(\POWERLED.func_state_RNI12ASZ0Z_1_cascade_ ));
    InMux I__6917 (
            .O(N__30785),
            .I(N__30778));
    InMux I__6916 (
            .O(N__30784),
            .I(N__30775));
    InMux I__6915 (
            .O(N__30783),
            .I(N__30770));
    InMux I__6914 (
            .O(N__30782),
            .I(N__30770));
    InMux I__6913 (
            .O(N__30781),
            .I(N__30766));
    LocalMux I__6912 (
            .O(N__30778),
            .I(N__30759));
    LocalMux I__6911 (
            .O(N__30775),
            .I(N__30759));
    LocalMux I__6910 (
            .O(N__30770),
            .I(N__30759));
    InMux I__6909 (
            .O(N__30769),
            .I(N__30756));
    LocalMux I__6908 (
            .O(N__30766),
            .I(N__30751));
    Span4Mux_s1_h I__6907 (
            .O(N__30759),
            .I(N__30751));
    LocalMux I__6906 (
            .O(N__30756),
            .I(N__30748));
    Span4Mux_h I__6905 (
            .O(N__30751),
            .I(N__30745));
    Odrv12 I__6904 (
            .O(N__30748),
            .I(\POWERLED.N_613 ));
    Odrv4 I__6903 (
            .O(N__30745),
            .I(\POWERLED.N_613 ));
    InMux I__6902 (
            .O(N__30740),
            .I(N__30729));
    CascadeMux I__6901 (
            .O(N__30739),
            .I(N__30724));
    InMux I__6900 (
            .O(N__30738),
            .I(N__30713));
    InMux I__6899 (
            .O(N__30737),
            .I(N__30713));
    InMux I__6898 (
            .O(N__30736),
            .I(N__30713));
    InMux I__6897 (
            .O(N__30735),
            .I(N__30710));
    InMux I__6896 (
            .O(N__30734),
            .I(N__30700));
    InMux I__6895 (
            .O(N__30733),
            .I(N__30700));
    InMux I__6894 (
            .O(N__30732),
            .I(N__30697));
    LocalMux I__6893 (
            .O(N__30729),
            .I(N__30691));
    InMux I__6892 (
            .O(N__30728),
            .I(N__30688));
    InMux I__6891 (
            .O(N__30727),
            .I(N__30684));
    InMux I__6890 (
            .O(N__30724),
            .I(N__30681));
    InMux I__6889 (
            .O(N__30723),
            .I(N__30676));
    InMux I__6888 (
            .O(N__30722),
            .I(N__30676));
    CascadeMux I__6887 (
            .O(N__30721),
            .I(N__30673));
    InMux I__6886 (
            .O(N__30720),
            .I(N__30667));
    LocalMux I__6885 (
            .O(N__30713),
            .I(N__30659));
    LocalMux I__6884 (
            .O(N__30710),
            .I(N__30659));
    InMux I__6883 (
            .O(N__30709),
            .I(N__30656));
    InMux I__6882 (
            .O(N__30708),
            .I(N__30647));
    InMux I__6881 (
            .O(N__30707),
            .I(N__30647));
    InMux I__6880 (
            .O(N__30706),
            .I(N__30647));
    InMux I__6879 (
            .O(N__30705),
            .I(N__30647));
    LocalMux I__6878 (
            .O(N__30700),
            .I(N__30642));
    LocalMux I__6877 (
            .O(N__30697),
            .I(N__30642));
    InMux I__6876 (
            .O(N__30696),
            .I(N__30639));
    InMux I__6875 (
            .O(N__30695),
            .I(N__30634));
    InMux I__6874 (
            .O(N__30694),
            .I(N__30634));
    Span4Mux_s0_h I__6873 (
            .O(N__30691),
            .I(N__30629));
    LocalMux I__6872 (
            .O(N__30688),
            .I(N__30629));
    InMux I__6871 (
            .O(N__30687),
            .I(N__30626));
    LocalMux I__6870 (
            .O(N__30684),
            .I(N__30619));
    LocalMux I__6869 (
            .O(N__30681),
            .I(N__30619));
    LocalMux I__6868 (
            .O(N__30676),
            .I(N__30619));
    InMux I__6867 (
            .O(N__30673),
            .I(N__30612));
    InMux I__6866 (
            .O(N__30672),
            .I(N__30612));
    InMux I__6865 (
            .O(N__30671),
            .I(N__30612));
    InMux I__6864 (
            .O(N__30670),
            .I(N__30609));
    LocalMux I__6863 (
            .O(N__30667),
            .I(N__30606));
    InMux I__6862 (
            .O(N__30666),
            .I(N__30603));
    CascadeMux I__6861 (
            .O(N__30665),
            .I(N__30599));
    CascadeMux I__6860 (
            .O(N__30664),
            .I(N__30595));
    Span4Mux_v I__6859 (
            .O(N__30659),
            .I(N__30588));
    LocalMux I__6858 (
            .O(N__30656),
            .I(N__30588));
    LocalMux I__6857 (
            .O(N__30647),
            .I(N__30588));
    Span4Mux_v I__6856 (
            .O(N__30642),
            .I(N__30581));
    LocalMux I__6855 (
            .O(N__30639),
            .I(N__30581));
    LocalMux I__6854 (
            .O(N__30634),
            .I(N__30581));
    Span4Mux_v I__6853 (
            .O(N__30629),
            .I(N__30572));
    LocalMux I__6852 (
            .O(N__30626),
            .I(N__30569));
    Span4Mux_v I__6851 (
            .O(N__30619),
            .I(N__30564));
    LocalMux I__6850 (
            .O(N__30612),
            .I(N__30564));
    LocalMux I__6849 (
            .O(N__30609),
            .I(N__30557));
    Span4Mux_v I__6848 (
            .O(N__30606),
            .I(N__30557));
    LocalMux I__6847 (
            .O(N__30603),
            .I(N__30557));
    InMux I__6846 (
            .O(N__30602),
            .I(N__30554));
    InMux I__6845 (
            .O(N__30599),
            .I(N__30551));
    InMux I__6844 (
            .O(N__30598),
            .I(N__30545));
    InMux I__6843 (
            .O(N__30595),
            .I(N__30545));
    Span4Mux_v I__6842 (
            .O(N__30588),
            .I(N__30540));
    Span4Mux_v I__6841 (
            .O(N__30581),
            .I(N__30540));
    InMux I__6840 (
            .O(N__30580),
            .I(N__30533));
    InMux I__6839 (
            .O(N__30579),
            .I(N__30533));
    InMux I__6838 (
            .O(N__30578),
            .I(N__30533));
    InMux I__6837 (
            .O(N__30577),
            .I(N__30526));
    InMux I__6836 (
            .O(N__30576),
            .I(N__30526));
    InMux I__6835 (
            .O(N__30575),
            .I(N__30526));
    Span4Mux_v I__6834 (
            .O(N__30572),
            .I(N__30521));
    Span4Mux_v I__6833 (
            .O(N__30569),
            .I(N__30521));
    Span4Mux_v I__6832 (
            .O(N__30564),
            .I(N__30514));
    Span4Mux_h I__6831 (
            .O(N__30557),
            .I(N__30514));
    LocalMux I__6830 (
            .O(N__30554),
            .I(N__30514));
    LocalMux I__6829 (
            .O(N__30551),
            .I(N__30511));
    InMux I__6828 (
            .O(N__30550),
            .I(N__30508));
    LocalMux I__6827 (
            .O(N__30545),
            .I(N__30501));
    Sp12to4 I__6826 (
            .O(N__30540),
            .I(N__30501));
    LocalMux I__6825 (
            .O(N__30533),
            .I(N__30501));
    LocalMux I__6824 (
            .O(N__30526),
            .I(N__30498));
    Span4Mux_h I__6823 (
            .O(N__30521),
            .I(N__30493));
    Span4Mux_v I__6822 (
            .O(N__30514),
            .I(N__30493));
    Span4Mux_h I__6821 (
            .O(N__30511),
            .I(N__30488));
    LocalMux I__6820 (
            .O(N__30508),
            .I(N__30488));
    Span12Mux_s8_h I__6819 (
            .O(N__30501),
            .I(N__30485));
    Span12Mux_s8_h I__6818 (
            .O(N__30498),
            .I(N__30482));
    IoSpan4Mux I__6817 (
            .O(N__30493),
            .I(N__30477));
    IoSpan4Mux I__6816 (
            .O(N__30488),
            .I(N__30477));
    Odrv12 I__6815 (
            .O(N__30485),
            .I(slp_s4n));
    Odrv12 I__6814 (
            .O(N__30482),
            .I(slp_s4n));
    Odrv4 I__6813 (
            .O(N__30477),
            .I(slp_s4n));
    InMux I__6812 (
            .O(N__30470),
            .I(N__30464));
    InMux I__6811 (
            .O(N__30469),
            .I(N__30464));
    LocalMux I__6810 (
            .O(N__30464),
            .I(N__30461));
    Span4Mux_v I__6809 (
            .O(N__30461),
            .I(N__30458));
    Odrv4 I__6808 (
            .O(N__30458),
            .I(\POWERLED.func_state_RNI8AQHZ0Z_0 ));
    InMux I__6807 (
            .O(N__30455),
            .I(N__30452));
    LocalMux I__6806 (
            .O(N__30452),
            .I(N__30449));
    Span12Mux_s6_v I__6805 (
            .O(N__30449),
            .I(N__30446));
    Odrv12 I__6804 (
            .O(N__30446),
            .I(\POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ));
    InMux I__6803 (
            .O(N__30443),
            .I(N__30437));
    InMux I__6802 (
            .O(N__30442),
            .I(N__30437));
    LocalMux I__6801 (
            .O(N__30437),
            .I(\POWERLED.func_state_RNI12ASZ0Z_1 ));
    InMux I__6800 (
            .O(N__30434),
            .I(N__30428));
    InMux I__6799 (
            .O(N__30433),
            .I(N__30428));
    LocalMux I__6798 (
            .O(N__30428),
            .I(N__30425));
    Odrv4 I__6797 (
            .O(N__30425),
            .I(\POWERLED.N_83 ));
    CascadeMux I__6796 (
            .O(N__30422),
            .I(N__30417));
    InMux I__6795 (
            .O(N__30421),
            .I(N__30402));
    InMux I__6794 (
            .O(N__30420),
            .I(N__30402));
    InMux I__6793 (
            .O(N__30417),
            .I(N__30402));
    InMux I__6792 (
            .O(N__30416),
            .I(N__30395));
    InMux I__6791 (
            .O(N__30415),
            .I(N__30395));
    InMux I__6790 (
            .O(N__30414),
            .I(N__30395));
    InMux I__6789 (
            .O(N__30413),
            .I(N__30390));
    InMux I__6788 (
            .O(N__30412),
            .I(N__30390));
    CascadeMux I__6787 (
            .O(N__30411),
            .I(N__30384));
    CascadeMux I__6786 (
            .O(N__30410),
            .I(N__30381));
    CascadeMux I__6785 (
            .O(N__30409),
            .I(N__30378));
    LocalMux I__6784 (
            .O(N__30402),
            .I(N__30374));
    LocalMux I__6783 (
            .O(N__30395),
            .I(N__30369));
    LocalMux I__6782 (
            .O(N__30390),
            .I(N__30369));
    InMux I__6781 (
            .O(N__30389),
            .I(N__30364));
    InMux I__6780 (
            .O(N__30388),
            .I(N__30364));
    InMux I__6779 (
            .O(N__30387),
            .I(N__30355));
    InMux I__6778 (
            .O(N__30384),
            .I(N__30355));
    InMux I__6777 (
            .O(N__30381),
            .I(N__30355));
    InMux I__6776 (
            .O(N__30378),
            .I(N__30355));
    CascadeMux I__6775 (
            .O(N__30377),
            .I(N__30349));
    Span4Mux_h I__6774 (
            .O(N__30374),
            .I(N__30337));
    Span4Mux_v I__6773 (
            .O(N__30369),
            .I(N__30337));
    LocalMux I__6772 (
            .O(N__30364),
            .I(N__30337));
    LocalMux I__6771 (
            .O(N__30355),
            .I(N__30337));
    InMux I__6770 (
            .O(N__30354),
            .I(N__30332));
    InMux I__6769 (
            .O(N__30353),
            .I(N__30332));
    InMux I__6768 (
            .O(N__30352),
            .I(N__30325));
    InMux I__6767 (
            .O(N__30349),
            .I(N__30325));
    InMux I__6766 (
            .O(N__30348),
            .I(N__30325));
    CascadeMux I__6765 (
            .O(N__30347),
            .I(N__30322));
    CascadeMux I__6764 (
            .O(N__30346),
            .I(N__30319));
    Span4Mux_v I__6763 (
            .O(N__30337),
            .I(N__30311));
    LocalMux I__6762 (
            .O(N__30332),
            .I(N__30306));
    LocalMux I__6761 (
            .O(N__30325),
            .I(N__30306));
    InMux I__6760 (
            .O(N__30322),
            .I(N__30299));
    InMux I__6759 (
            .O(N__30319),
            .I(N__30299));
    InMux I__6758 (
            .O(N__30318),
            .I(N__30299));
    InMux I__6757 (
            .O(N__30317),
            .I(N__30296));
    CascadeMux I__6756 (
            .O(N__30316),
            .I(N__30293));
    CascadeMux I__6755 (
            .O(N__30315),
            .I(N__30290));
    CascadeMux I__6754 (
            .O(N__30314),
            .I(N__30285));
    Span4Mux_h I__6753 (
            .O(N__30311),
            .I(N__30281));
    Span4Mux_v I__6752 (
            .O(N__30306),
            .I(N__30274));
    LocalMux I__6751 (
            .O(N__30299),
            .I(N__30274));
    LocalMux I__6750 (
            .O(N__30296),
            .I(N__30274));
    InMux I__6749 (
            .O(N__30293),
            .I(N__30267));
    InMux I__6748 (
            .O(N__30290),
            .I(N__30267));
    InMux I__6747 (
            .O(N__30289),
            .I(N__30267));
    InMux I__6746 (
            .O(N__30288),
            .I(N__30259));
    InMux I__6745 (
            .O(N__30285),
            .I(N__30259));
    CascadeMux I__6744 (
            .O(N__30284),
            .I(N__30255));
    IoSpan4Mux I__6743 (
            .O(N__30281),
            .I(N__30248));
    Span4Mux_v I__6742 (
            .O(N__30274),
            .I(N__30248));
    LocalMux I__6741 (
            .O(N__30267),
            .I(N__30248));
    InMux I__6740 (
            .O(N__30266),
            .I(N__30245));
    CascadeMux I__6739 (
            .O(N__30265),
            .I(N__30240));
    CascadeMux I__6738 (
            .O(N__30264),
            .I(N__30236));
    LocalMux I__6737 (
            .O(N__30259),
            .I(N__30232));
    InMux I__6736 (
            .O(N__30258),
            .I(N__30229));
    InMux I__6735 (
            .O(N__30255),
            .I(N__30224));
    IoSpan4Mux I__6734 (
            .O(N__30248),
            .I(N__30221));
    LocalMux I__6733 (
            .O(N__30245),
            .I(N__30218));
    InMux I__6732 (
            .O(N__30244),
            .I(N__30213));
    InMux I__6731 (
            .O(N__30243),
            .I(N__30213));
    InMux I__6730 (
            .O(N__30240),
            .I(N__30208));
    InMux I__6729 (
            .O(N__30239),
            .I(N__30208));
    InMux I__6728 (
            .O(N__30236),
            .I(N__30205));
    InMux I__6727 (
            .O(N__30235),
            .I(N__30202));
    Span4Mux_h I__6726 (
            .O(N__30232),
            .I(N__30197));
    LocalMux I__6725 (
            .O(N__30229),
            .I(N__30197));
    InMux I__6724 (
            .O(N__30228),
            .I(N__30192));
    InMux I__6723 (
            .O(N__30227),
            .I(N__30192));
    LocalMux I__6722 (
            .O(N__30224),
            .I(N__30189));
    IoSpan4Mux I__6721 (
            .O(N__30221),
            .I(N__30186));
    Span12Mux_s10_h I__6720 (
            .O(N__30218),
            .I(N__30177));
    LocalMux I__6719 (
            .O(N__30213),
            .I(N__30177));
    LocalMux I__6718 (
            .O(N__30208),
            .I(N__30177));
    LocalMux I__6717 (
            .O(N__30205),
            .I(N__30177));
    LocalMux I__6716 (
            .O(N__30202),
            .I(N__30174));
    Span4Mux_v I__6715 (
            .O(N__30197),
            .I(N__30169));
    LocalMux I__6714 (
            .O(N__30192),
            .I(N__30169));
    Odrv12 I__6713 (
            .O(N__30189),
            .I(slp_s3n));
    Odrv4 I__6712 (
            .O(N__30186),
            .I(slp_s3n));
    Odrv12 I__6711 (
            .O(N__30177),
            .I(slp_s3n));
    Odrv4 I__6710 (
            .O(N__30174),
            .I(slp_s3n));
    Odrv4 I__6709 (
            .O(N__30169),
            .I(slp_s3n));
    CascadeMux I__6708 (
            .O(N__30158),
            .I(N__30154));
    InMux I__6707 (
            .O(N__30157),
            .I(N__30134));
    InMux I__6706 (
            .O(N__30154),
            .I(N__30134));
    InMux I__6705 (
            .O(N__30153),
            .I(N__30134));
    InMux I__6704 (
            .O(N__30152),
            .I(N__30134));
    InMux I__6703 (
            .O(N__30151),
            .I(N__30129));
    InMux I__6702 (
            .O(N__30150),
            .I(N__30129));
    InMux I__6701 (
            .O(N__30149),
            .I(N__30126));
    CascadeMux I__6700 (
            .O(N__30148),
            .I(N__30119));
    InMux I__6699 (
            .O(N__30147),
            .I(N__30112));
    InMux I__6698 (
            .O(N__30146),
            .I(N__30109));
    CascadeMux I__6697 (
            .O(N__30145),
            .I(N__30106));
    InMux I__6696 (
            .O(N__30144),
            .I(N__30102));
    InMux I__6695 (
            .O(N__30143),
            .I(N__30099));
    LocalMux I__6694 (
            .O(N__30134),
            .I(N__30096));
    LocalMux I__6693 (
            .O(N__30129),
            .I(N__30091));
    LocalMux I__6692 (
            .O(N__30126),
            .I(N__30091));
    InMux I__6691 (
            .O(N__30125),
            .I(N__30086));
    InMux I__6690 (
            .O(N__30124),
            .I(N__30086));
    InMux I__6689 (
            .O(N__30123),
            .I(N__30083));
    InMux I__6688 (
            .O(N__30122),
            .I(N__30080));
    InMux I__6687 (
            .O(N__30119),
            .I(N__30076));
    InMux I__6686 (
            .O(N__30118),
            .I(N__30070));
    InMux I__6685 (
            .O(N__30117),
            .I(N__30065));
    InMux I__6684 (
            .O(N__30116),
            .I(N__30065));
    InMux I__6683 (
            .O(N__30115),
            .I(N__30062));
    LocalMux I__6682 (
            .O(N__30112),
            .I(N__30058));
    LocalMux I__6681 (
            .O(N__30109),
            .I(N__30055));
    InMux I__6680 (
            .O(N__30106),
            .I(N__30050));
    InMux I__6679 (
            .O(N__30105),
            .I(N__30050));
    LocalMux I__6678 (
            .O(N__30102),
            .I(N__30046));
    LocalMux I__6677 (
            .O(N__30099),
            .I(N__30037));
    Span4Mux_v I__6676 (
            .O(N__30096),
            .I(N__30037));
    Span4Mux_s3_v I__6675 (
            .O(N__30091),
            .I(N__30037));
    LocalMux I__6674 (
            .O(N__30086),
            .I(N__30037));
    LocalMux I__6673 (
            .O(N__30083),
            .I(N__30032));
    LocalMux I__6672 (
            .O(N__30080),
            .I(N__30032));
    InMux I__6671 (
            .O(N__30079),
            .I(N__30029));
    LocalMux I__6670 (
            .O(N__30076),
            .I(N__30026));
    InMux I__6669 (
            .O(N__30075),
            .I(N__30023));
    CascadeMux I__6668 (
            .O(N__30074),
            .I(N__30019));
    InMux I__6667 (
            .O(N__30073),
            .I(N__30015));
    LocalMux I__6666 (
            .O(N__30070),
            .I(N__30005));
    LocalMux I__6665 (
            .O(N__30065),
            .I(N__30005));
    LocalMux I__6664 (
            .O(N__30062),
            .I(N__30005));
    InMux I__6663 (
            .O(N__30061),
            .I(N__30002));
    Span4Mux_s2_h I__6662 (
            .O(N__30058),
            .I(N__29997));
    Span4Mux_s2_h I__6661 (
            .O(N__30055),
            .I(N__29997));
    LocalMux I__6660 (
            .O(N__30050),
            .I(N__29994));
    InMux I__6659 (
            .O(N__30049),
            .I(N__29991));
    Span4Mux_v I__6658 (
            .O(N__30046),
            .I(N__29982));
    Span4Mux_v I__6657 (
            .O(N__30037),
            .I(N__29982));
    Span4Mux_v I__6656 (
            .O(N__30032),
            .I(N__29982));
    LocalMux I__6655 (
            .O(N__30029),
            .I(N__29982));
    Span12Mux_s5_h I__6654 (
            .O(N__30026),
            .I(N__29977));
    LocalMux I__6653 (
            .O(N__30023),
            .I(N__29974));
    InMux I__6652 (
            .O(N__30022),
            .I(N__29969));
    InMux I__6651 (
            .O(N__30019),
            .I(N__29969));
    InMux I__6650 (
            .O(N__30018),
            .I(N__29966));
    LocalMux I__6649 (
            .O(N__30015),
            .I(N__29963));
    InMux I__6648 (
            .O(N__30014),
            .I(N__29960));
    InMux I__6647 (
            .O(N__30013),
            .I(N__29955));
    InMux I__6646 (
            .O(N__30012),
            .I(N__29955));
    Span4Mux_v I__6645 (
            .O(N__30005),
            .I(N__29946));
    LocalMux I__6644 (
            .O(N__30002),
            .I(N__29946));
    Span4Mux_v I__6643 (
            .O(N__29997),
            .I(N__29946));
    Span4Mux_s2_h I__6642 (
            .O(N__29994),
            .I(N__29946));
    LocalMux I__6641 (
            .O(N__29991),
            .I(N__29941));
    Span4Mux_h I__6640 (
            .O(N__29982),
            .I(N__29941));
    InMux I__6639 (
            .O(N__29981),
            .I(N__29936));
    InMux I__6638 (
            .O(N__29980),
            .I(N__29936));
    Odrv12 I__6637 (
            .O(N__29977),
            .I(func_state_RNIMJ6IF_0_1));
    Odrv4 I__6636 (
            .O(N__29974),
            .I(func_state_RNIMJ6IF_0_1));
    LocalMux I__6635 (
            .O(N__29969),
            .I(func_state_RNIMJ6IF_0_1));
    LocalMux I__6634 (
            .O(N__29966),
            .I(func_state_RNIMJ6IF_0_1));
    Odrv4 I__6633 (
            .O(N__29963),
            .I(func_state_RNIMJ6IF_0_1));
    LocalMux I__6632 (
            .O(N__29960),
            .I(func_state_RNIMJ6IF_0_1));
    LocalMux I__6631 (
            .O(N__29955),
            .I(func_state_RNIMJ6IF_0_1));
    Odrv4 I__6630 (
            .O(N__29946),
            .I(func_state_RNIMJ6IF_0_1));
    Odrv4 I__6629 (
            .O(N__29941),
            .I(func_state_RNIMJ6IF_0_1));
    LocalMux I__6628 (
            .O(N__29936),
            .I(func_state_RNIMJ6IF_0_1));
    InMux I__6627 (
            .O(N__29915),
            .I(N__29909));
    InMux I__6626 (
            .O(N__29914),
            .I(N__29904));
    InMux I__6625 (
            .O(N__29913),
            .I(N__29904));
    CascadeMux I__6624 (
            .O(N__29912),
            .I(N__29901));
    LocalMux I__6623 (
            .O(N__29909),
            .I(N__29889));
    LocalMux I__6622 (
            .O(N__29904),
            .I(N__29886));
    InMux I__6621 (
            .O(N__29901),
            .I(N__29881));
    InMux I__6620 (
            .O(N__29900),
            .I(N__29881));
    InMux I__6619 (
            .O(N__29899),
            .I(N__29876));
    InMux I__6618 (
            .O(N__29898),
            .I(N__29876));
    InMux I__6617 (
            .O(N__29897),
            .I(N__29869));
    InMux I__6616 (
            .O(N__29896),
            .I(N__29869));
    InMux I__6615 (
            .O(N__29895),
            .I(N__29869));
    InMux I__6614 (
            .O(N__29894),
            .I(N__29866));
    InMux I__6613 (
            .O(N__29893),
            .I(N__29863));
    InMux I__6612 (
            .O(N__29892),
            .I(N__29859));
    Span4Mux_s3_v I__6611 (
            .O(N__29889),
            .I(N__29848));
    Span4Mux_h I__6610 (
            .O(N__29886),
            .I(N__29848));
    LocalMux I__6609 (
            .O(N__29881),
            .I(N__29848));
    LocalMux I__6608 (
            .O(N__29876),
            .I(N__29848));
    LocalMux I__6607 (
            .O(N__29869),
            .I(N__29848));
    LocalMux I__6606 (
            .O(N__29866),
            .I(N__29845));
    LocalMux I__6605 (
            .O(N__29863),
            .I(N__29841));
    InMux I__6604 (
            .O(N__29862),
            .I(N__29838));
    LocalMux I__6603 (
            .O(N__29859),
            .I(N__29833));
    Span4Mux_v I__6602 (
            .O(N__29848),
            .I(N__29833));
    Span12Mux_s4_v I__6601 (
            .O(N__29845),
            .I(N__29830));
    InMux I__6600 (
            .O(N__29844),
            .I(N__29827));
    Span4Mux_h I__6599 (
            .O(N__29841),
            .I(N__29820));
    LocalMux I__6598 (
            .O(N__29838),
            .I(N__29820));
    Span4Mux_h I__6597 (
            .O(N__29833),
            .I(N__29820));
    Odrv12 I__6596 (
            .O(N__29830),
            .I(RSMRSTn_rep2));
    LocalMux I__6595 (
            .O(N__29827),
            .I(RSMRSTn_rep2));
    Odrv4 I__6594 (
            .O(N__29820),
            .I(RSMRSTn_rep2));
    InMux I__6593 (
            .O(N__29813),
            .I(N__29809));
    InMux I__6592 (
            .O(N__29812),
            .I(N__29806));
    LocalMux I__6591 (
            .O(N__29809),
            .I(N__29802));
    LocalMux I__6590 (
            .O(N__29806),
            .I(N__29799));
    InMux I__6589 (
            .O(N__29805),
            .I(N__29796));
    Odrv4 I__6588 (
            .O(N__29802),
            .I(\POWERLED.N_531 ));
    Odrv4 I__6587 (
            .O(N__29799),
            .I(\POWERLED.N_531 ));
    LocalMux I__6586 (
            .O(N__29796),
            .I(\POWERLED.N_531 ));
    InMux I__6585 (
            .O(N__29789),
            .I(N__29786));
    LocalMux I__6584 (
            .O(N__29786),
            .I(N__29783));
    Span4Mux_v I__6583 (
            .O(N__29783),
            .I(N__29780));
    Sp12to4 I__6582 (
            .O(N__29780),
            .I(N__29777));
    Span12Mux_s3_h I__6581 (
            .O(N__29777),
            .I(N__29774));
    Odrv12 I__6580 (
            .O(N__29774),
            .I(\POWERLED.un1_clk_100khz_51_and_i_3_0 ));
    CascadeMux I__6579 (
            .O(N__29771),
            .I(\POWERLED.N_532_cascade_ ));
    InMux I__6578 (
            .O(N__29768),
            .I(N__29765));
    LocalMux I__6577 (
            .O(N__29765),
            .I(\POWERLED.N_530 ));
    CascadeMux I__6576 (
            .O(N__29762),
            .I(\POWERLED.dutycycle_RNI_8Z0Z_5_cascade_ ));
    CascadeMux I__6575 (
            .O(N__29759),
            .I(N__29754));
    InMux I__6574 (
            .O(N__29758),
            .I(N__29749));
    InMux I__6573 (
            .O(N__29757),
            .I(N__29749));
    InMux I__6572 (
            .O(N__29754),
            .I(N__29745));
    LocalMux I__6571 (
            .O(N__29749),
            .I(N__29739));
    InMux I__6570 (
            .O(N__29748),
            .I(N__29736));
    LocalMux I__6569 (
            .O(N__29745),
            .I(N__29733));
    InMux I__6568 (
            .O(N__29744),
            .I(N__29730));
    CascadeMux I__6567 (
            .O(N__29743),
            .I(N__29727));
    CascadeMux I__6566 (
            .O(N__29742),
            .I(N__29722));
    Span4Mux_s3_v I__6565 (
            .O(N__29739),
            .I(N__29717));
    LocalMux I__6564 (
            .O(N__29736),
            .I(N__29717));
    Span4Mux_s3_v I__6563 (
            .O(N__29733),
            .I(N__29712));
    LocalMux I__6562 (
            .O(N__29730),
            .I(N__29712));
    InMux I__6561 (
            .O(N__29727),
            .I(N__29709));
    InMux I__6560 (
            .O(N__29726),
            .I(N__29706));
    InMux I__6559 (
            .O(N__29725),
            .I(N__29703));
    InMux I__6558 (
            .O(N__29722),
            .I(N__29700));
    Span4Mux_v I__6557 (
            .O(N__29717),
            .I(N__29694));
    Span4Mux_v I__6556 (
            .O(N__29712),
            .I(N__29694));
    LocalMux I__6555 (
            .O(N__29709),
            .I(N__29691));
    LocalMux I__6554 (
            .O(N__29706),
            .I(N__29688));
    LocalMux I__6553 (
            .O(N__29703),
            .I(N__29683));
    LocalMux I__6552 (
            .O(N__29700),
            .I(N__29683));
    InMux I__6551 (
            .O(N__29699),
            .I(N__29680));
    Odrv4 I__6550 (
            .O(N__29694),
            .I(\POWERLED.N_251 ));
    Odrv4 I__6549 (
            .O(N__29691),
            .I(\POWERLED.N_251 ));
    Odrv12 I__6548 (
            .O(N__29688),
            .I(\POWERLED.N_251 ));
    Odrv12 I__6547 (
            .O(N__29683),
            .I(\POWERLED.N_251 ));
    LocalMux I__6546 (
            .O(N__29680),
            .I(\POWERLED.N_251 ));
    InMux I__6545 (
            .O(N__29669),
            .I(N__29665));
    CascadeMux I__6544 (
            .O(N__29668),
            .I(N__29662));
    LocalMux I__6543 (
            .O(N__29665),
            .I(N__29659));
    InMux I__6542 (
            .O(N__29662),
            .I(N__29656));
    Span4Mux_v I__6541 (
            .O(N__29659),
            .I(N__29651));
    LocalMux I__6540 (
            .O(N__29656),
            .I(N__29648));
    InMux I__6539 (
            .O(N__29655),
            .I(N__29645));
    InMux I__6538 (
            .O(N__29654),
            .I(N__29642));
    Odrv4 I__6537 (
            .O(N__29651),
            .I(\POWERLED.N_633 ));
    Odrv4 I__6536 (
            .O(N__29648),
            .I(\POWERLED.N_633 ));
    LocalMux I__6535 (
            .O(N__29645),
            .I(\POWERLED.N_633 ));
    LocalMux I__6534 (
            .O(N__29642),
            .I(\POWERLED.N_633 ));
    CascadeMux I__6533 (
            .O(N__29633),
            .I(\POWERLED.func_state_RNIOGRSZ0Z_1_cascade_ ));
    IoInMux I__6532 (
            .O(N__29630),
            .I(N__29627));
    LocalMux I__6531 (
            .O(N__29627),
            .I(N__29623));
    IoInMux I__6530 (
            .O(N__29626),
            .I(N__29620));
    IoSpan4Mux I__6529 (
            .O(N__29623),
            .I(N__29614));
    LocalMux I__6528 (
            .O(N__29620),
            .I(N__29611));
    InMux I__6527 (
            .O(N__29619),
            .I(N__29605));
    CascadeMux I__6526 (
            .O(N__29618),
            .I(N__29601));
    InMux I__6525 (
            .O(N__29617),
            .I(N__29597));
    Span4Mux_s0_h I__6524 (
            .O(N__29614),
            .I(N__29594));
    Span4Mux_s0_h I__6523 (
            .O(N__29611),
            .I(N__29591));
    InMux I__6522 (
            .O(N__29610),
            .I(N__29586));
    InMux I__6521 (
            .O(N__29609),
            .I(N__29586));
    InMux I__6520 (
            .O(N__29608),
            .I(N__29583));
    LocalMux I__6519 (
            .O(N__29605),
            .I(N__29580));
    InMux I__6518 (
            .O(N__29604),
            .I(N__29577));
    InMux I__6517 (
            .O(N__29601),
            .I(N__29574));
    InMux I__6516 (
            .O(N__29600),
            .I(N__29569));
    LocalMux I__6515 (
            .O(N__29597),
            .I(N__29566));
    Sp12to4 I__6514 (
            .O(N__29594),
            .I(N__29559));
    Sp12to4 I__6513 (
            .O(N__29591),
            .I(N__29559));
    LocalMux I__6512 (
            .O(N__29586),
            .I(N__29559));
    LocalMux I__6511 (
            .O(N__29583),
            .I(N__29554));
    Span4Mux_v I__6510 (
            .O(N__29580),
            .I(N__29547));
    LocalMux I__6509 (
            .O(N__29577),
            .I(N__29547));
    LocalMux I__6508 (
            .O(N__29574),
            .I(N__29547));
    InMux I__6507 (
            .O(N__29573),
            .I(N__29544));
    InMux I__6506 (
            .O(N__29572),
            .I(N__29541));
    LocalMux I__6505 (
            .O(N__29569),
            .I(N__29538));
    Span4Mux_h I__6504 (
            .O(N__29566),
            .I(N__29533));
    Span12Mux_s10_v I__6503 (
            .O(N__29559),
            .I(N__29530));
    InMux I__6502 (
            .O(N__29558),
            .I(N__29527));
    InMux I__6501 (
            .O(N__29557),
            .I(N__29524));
    Span4Mux_v I__6500 (
            .O(N__29554),
            .I(N__29521));
    Span4Mux_v I__6499 (
            .O(N__29547),
            .I(N__29518));
    LocalMux I__6498 (
            .O(N__29544),
            .I(N__29511));
    LocalMux I__6497 (
            .O(N__29541),
            .I(N__29511));
    Span4Mux_s3_h I__6496 (
            .O(N__29538),
            .I(N__29511));
    InMux I__6495 (
            .O(N__29537),
            .I(N__29506));
    InMux I__6494 (
            .O(N__29536),
            .I(N__29506));
    Odrv4 I__6493 (
            .O(N__29533),
            .I(v5s_enn));
    Odrv12 I__6492 (
            .O(N__29530),
            .I(v5s_enn));
    LocalMux I__6491 (
            .O(N__29527),
            .I(v5s_enn));
    LocalMux I__6490 (
            .O(N__29524),
            .I(v5s_enn));
    Odrv4 I__6489 (
            .O(N__29521),
            .I(v5s_enn));
    Odrv4 I__6488 (
            .O(N__29518),
            .I(v5s_enn));
    Odrv4 I__6487 (
            .O(N__29511),
            .I(v5s_enn));
    LocalMux I__6486 (
            .O(N__29506),
            .I(v5s_enn));
    InMux I__6485 (
            .O(N__29489),
            .I(N__29486));
    LocalMux I__6484 (
            .O(N__29486),
            .I(N__29481));
    InMux I__6483 (
            .O(N__29485),
            .I(N__29476));
    InMux I__6482 (
            .O(N__29484),
            .I(N__29476));
    Odrv12 I__6481 (
            .O(N__29481),
            .I(\POWERLED.N_413_N ));
    LocalMux I__6480 (
            .O(N__29476),
            .I(\POWERLED.N_413_N ));
    CascadeMux I__6479 (
            .O(N__29471),
            .I(N__29467));
    InMux I__6478 (
            .O(N__29470),
            .I(N__29462));
    InMux I__6477 (
            .O(N__29467),
            .I(N__29462));
    LocalMux I__6476 (
            .O(N__29462),
            .I(\POWERLED.dutycycle_0_6 ));
    CascadeMux I__6475 (
            .O(N__29459),
            .I(\POWERLED.dutycycleZ0Z_6_cascade_ ));
    InMux I__6474 (
            .O(N__29456),
            .I(N__29452));
    InMux I__6473 (
            .O(N__29455),
            .I(N__29449));
    LocalMux I__6472 (
            .O(N__29452),
            .I(N__29446));
    LocalMux I__6471 (
            .O(N__29449),
            .I(N__29443));
    Span4Mux_v I__6470 (
            .O(N__29446),
            .I(N__29437));
    Span4Mux_s1_h I__6469 (
            .O(N__29443),
            .I(N__29437));
    InMux I__6468 (
            .O(N__29442),
            .I(N__29434));
    Span4Mux_h I__6467 (
            .O(N__29437),
            .I(N__29429));
    LocalMux I__6466 (
            .O(N__29434),
            .I(N__29429));
    Span4Mux_v I__6465 (
            .O(N__29429),
            .I(N__29426));
    Odrv4 I__6464 (
            .O(N__29426),
            .I(\POWERLED.N_612 ));
    InMux I__6463 (
            .O(N__29423),
            .I(N__29420));
    LocalMux I__6462 (
            .O(N__29420),
            .I(N__29417));
    Span4Mux_h I__6461 (
            .O(N__29417),
            .I(N__29414));
    Odrv4 I__6460 (
            .O(N__29414),
            .I(\POWERLED.N_672 ));
    CascadeMux I__6459 (
            .O(N__29411),
            .I(\POWERLED.N_672_cascade_ ));
    InMux I__6458 (
            .O(N__29408),
            .I(N__29405));
    LocalMux I__6457 (
            .O(N__29405),
            .I(N__29402));
    Span4Mux_h I__6456 (
            .O(N__29402),
            .I(N__29399));
    Odrv4 I__6455 (
            .O(N__29399),
            .I(\POWERLED.un1_dutycycle_168_0 ));
    InMux I__6454 (
            .O(N__29396),
            .I(N__29390));
    InMux I__6453 (
            .O(N__29395),
            .I(N__29390));
    LocalMux I__6452 (
            .O(N__29390),
            .I(N__29385));
    InMux I__6451 (
            .O(N__29389),
            .I(N__29380));
    InMux I__6450 (
            .O(N__29388),
            .I(N__29380));
    Span4Mux_v I__6449 (
            .O(N__29385),
            .I(N__29377));
    LocalMux I__6448 (
            .O(N__29380),
            .I(N__29374));
    Odrv4 I__6447 (
            .O(N__29377),
            .I(\POWERLED.count_clk_RNIZ0Z_6 ));
    Odrv12 I__6446 (
            .O(N__29374),
            .I(\POWERLED.count_clk_RNIZ0Z_6 ));
    InMux I__6445 (
            .O(N__29369),
            .I(N__29366));
    LocalMux I__6444 (
            .O(N__29366),
            .I(N__29361));
    InMux I__6443 (
            .O(N__29365),
            .I(N__29356));
    InMux I__6442 (
            .O(N__29364),
            .I(N__29356));
    Span4Mux_v I__6441 (
            .O(N__29361),
            .I(N__29352));
    LocalMux I__6440 (
            .O(N__29356),
            .I(N__29349));
    InMux I__6439 (
            .O(N__29355),
            .I(N__29346));
    Odrv4 I__6438 (
            .O(N__29352),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_0 ));
    Odrv4 I__6437 (
            .O(N__29349),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_0 ));
    LocalMux I__6436 (
            .O(N__29346),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_0 ));
    CascadeMux I__6435 (
            .O(N__29339),
            .I(\POWERLED.N_412_i_cascade_ ));
    InMux I__6434 (
            .O(N__29336),
            .I(N__29332));
    InMux I__6433 (
            .O(N__29335),
            .I(N__29329));
    LocalMux I__6432 (
            .O(N__29332),
            .I(N__29326));
    LocalMux I__6431 (
            .O(N__29329),
            .I(N__29323));
    Span4Mux_v I__6430 (
            .O(N__29326),
            .I(N__29320));
    Span4Mux_s2_v I__6429 (
            .O(N__29323),
            .I(N__29317));
    Odrv4 I__6428 (
            .O(N__29320),
            .I(\POWERLED.N_604 ));
    Odrv4 I__6427 (
            .O(N__29317),
            .I(\POWERLED.N_604 ));
    CascadeMux I__6426 (
            .O(N__29312),
            .I(N__29309));
    InMux I__6425 (
            .O(N__29309),
            .I(N__29303));
    InMux I__6424 (
            .O(N__29308),
            .I(N__29303));
    LocalMux I__6423 (
            .O(N__29303),
            .I(N__29300));
    Span12Mux_s9_v I__6422 (
            .O(N__29300),
            .I(N__29297));
    Odrv12 I__6421 (
            .O(N__29297),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_3 ));
    CascadeMux I__6420 (
            .O(N__29294),
            .I(N__29288));
    InMux I__6419 (
            .O(N__29293),
            .I(N__29285));
    InMux I__6418 (
            .O(N__29292),
            .I(N__29282));
    InMux I__6417 (
            .O(N__29291),
            .I(N__29279));
    InMux I__6416 (
            .O(N__29288),
            .I(N__29276));
    LocalMux I__6415 (
            .O(N__29285),
            .I(N__29271));
    LocalMux I__6414 (
            .O(N__29282),
            .I(N__29268));
    LocalMux I__6413 (
            .O(N__29279),
            .I(N__29264));
    LocalMux I__6412 (
            .O(N__29276),
            .I(N__29261));
    InMux I__6411 (
            .O(N__29275),
            .I(N__29256));
    InMux I__6410 (
            .O(N__29274),
            .I(N__29256));
    Span4Mux_s3_h I__6409 (
            .O(N__29271),
            .I(N__29253));
    Span4Mux_v I__6408 (
            .O(N__29268),
            .I(N__29250));
    InMux I__6407 (
            .O(N__29267),
            .I(N__29247));
    Span4Mux_s3_h I__6406 (
            .O(N__29264),
            .I(N__29240));
    Span4Mux_v I__6405 (
            .O(N__29261),
            .I(N__29240));
    LocalMux I__6404 (
            .O(N__29256),
            .I(N__29240));
    Odrv4 I__6403 (
            .O(N__29253),
            .I(\POWERLED.N_435 ));
    Odrv4 I__6402 (
            .O(N__29250),
            .I(\POWERLED.N_435 ));
    LocalMux I__6401 (
            .O(N__29247),
            .I(\POWERLED.N_435 ));
    Odrv4 I__6400 (
            .O(N__29240),
            .I(\POWERLED.N_435 ));
    InMux I__6399 (
            .O(N__29231),
            .I(N__29227));
    CascadeMux I__6398 (
            .O(N__29230),
            .I(N__29224));
    LocalMux I__6397 (
            .O(N__29227),
            .I(N__29219));
    InMux I__6396 (
            .O(N__29224),
            .I(N__29216));
    CascadeMux I__6395 (
            .O(N__29223),
            .I(N__29213));
    InMux I__6394 (
            .O(N__29222),
            .I(N__29210));
    Span4Mux_v I__6393 (
            .O(N__29219),
            .I(N__29206));
    LocalMux I__6392 (
            .O(N__29216),
            .I(N__29203));
    InMux I__6391 (
            .O(N__29213),
            .I(N__29200));
    LocalMux I__6390 (
            .O(N__29210),
            .I(N__29197));
    InMux I__6389 (
            .O(N__29209),
            .I(N__29194));
    Span4Mux_h I__6388 (
            .O(N__29206),
            .I(N__29187));
    Span4Mux_h I__6387 (
            .O(N__29203),
            .I(N__29187));
    LocalMux I__6386 (
            .O(N__29200),
            .I(N__29187));
    Odrv4 I__6385 (
            .O(N__29197),
            .I(\POWERLED.N_412_i ));
    LocalMux I__6384 (
            .O(N__29194),
            .I(\POWERLED.N_412_i ));
    Odrv4 I__6383 (
            .O(N__29187),
            .I(\POWERLED.N_412_i ));
    InMux I__6382 (
            .O(N__29180),
            .I(N__29177));
    LocalMux I__6381 (
            .O(N__29177),
            .I(N__29174));
    Span4Mux_h I__6380 (
            .O(N__29174),
            .I(N__29170));
    InMux I__6379 (
            .O(N__29173),
            .I(N__29167));
    Odrv4 I__6378 (
            .O(N__29170),
            .I(\POWERLED.func_state_RNI_5Z0Z_1 ));
    LocalMux I__6377 (
            .O(N__29167),
            .I(\POWERLED.func_state_RNI_5Z0Z_1 ));
    InMux I__6376 (
            .O(N__29162),
            .I(N__29156));
    InMux I__6375 (
            .O(N__29161),
            .I(N__29156));
    LocalMux I__6374 (
            .O(N__29156),
            .I(N__29153));
    Odrv4 I__6373 (
            .O(N__29153),
            .I(\POWERLED.count_clk_1_13 ));
    InMux I__6372 (
            .O(N__29150),
            .I(N__29147));
    LocalMux I__6371 (
            .O(N__29147),
            .I(\POWERLED.count_clk_0_13 ));
    InMux I__6370 (
            .O(N__29144),
            .I(N__29141));
    LocalMux I__6369 (
            .O(N__29141),
            .I(N__29138));
    Odrv12 I__6368 (
            .O(N__29138),
            .I(\POWERLED.count_clkZ0Z_13 ));
    InMux I__6367 (
            .O(N__29135),
            .I(N__29126));
    InMux I__6366 (
            .O(N__29134),
            .I(N__29126));
    InMux I__6365 (
            .O(N__29133),
            .I(N__29126));
    LocalMux I__6364 (
            .O(N__29126),
            .I(N__29123));
    Odrv4 I__6363 (
            .O(N__29123),
            .I(\POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ));
    CascadeMux I__6362 (
            .O(N__29120),
            .I(N__29114));
    CascadeMux I__6361 (
            .O(N__29119),
            .I(N__29111));
    CEMux I__6360 (
            .O(N__29118),
            .I(N__29107));
    CEMux I__6359 (
            .O(N__29117),
            .I(N__29100));
    InMux I__6358 (
            .O(N__29114),
            .I(N__29092));
    InMux I__6357 (
            .O(N__29111),
            .I(N__29092));
    CEMux I__6356 (
            .O(N__29110),
            .I(N__29092));
    LocalMux I__6355 (
            .O(N__29107),
            .I(N__29089));
    CEMux I__6354 (
            .O(N__29106),
            .I(N__29086));
    CascadeMux I__6353 (
            .O(N__29105),
            .I(N__29083));
    CascadeMux I__6352 (
            .O(N__29104),
            .I(N__29077));
    CEMux I__6351 (
            .O(N__29103),
            .I(N__29071));
    LocalMux I__6350 (
            .O(N__29100),
            .I(N__29066));
    InMux I__6349 (
            .O(N__29099),
            .I(N__29063));
    LocalMux I__6348 (
            .O(N__29092),
            .I(N__29057));
    Span4Mux_v I__6347 (
            .O(N__29089),
            .I(N__29052));
    LocalMux I__6346 (
            .O(N__29086),
            .I(N__29052));
    InMux I__6345 (
            .O(N__29083),
            .I(N__29047));
    InMux I__6344 (
            .O(N__29082),
            .I(N__29047));
    InMux I__6343 (
            .O(N__29081),
            .I(N__29040));
    InMux I__6342 (
            .O(N__29080),
            .I(N__29040));
    InMux I__6341 (
            .O(N__29077),
            .I(N__29040));
    CEMux I__6340 (
            .O(N__29076),
            .I(N__29034));
    InMux I__6339 (
            .O(N__29075),
            .I(N__29031));
    InMux I__6338 (
            .O(N__29074),
            .I(N__29028));
    LocalMux I__6337 (
            .O(N__29071),
            .I(N__29025));
    InMux I__6336 (
            .O(N__29070),
            .I(N__29020));
    CEMux I__6335 (
            .O(N__29069),
            .I(N__29020));
    Span4Mux_v I__6334 (
            .O(N__29066),
            .I(N__29017));
    LocalMux I__6333 (
            .O(N__29063),
            .I(N__29014));
    InMux I__6332 (
            .O(N__29062),
            .I(N__29007));
    InMux I__6331 (
            .O(N__29061),
            .I(N__29007));
    InMux I__6330 (
            .O(N__29060),
            .I(N__29007));
    Span4Mux_v I__6329 (
            .O(N__29057),
            .I(N__29000));
    Span4Mux_s3_v I__6328 (
            .O(N__29052),
            .I(N__29000));
    LocalMux I__6327 (
            .O(N__29047),
            .I(N__29000));
    LocalMux I__6326 (
            .O(N__29040),
            .I(N__28997));
    InMux I__6325 (
            .O(N__29039),
            .I(N__28992));
    InMux I__6324 (
            .O(N__29038),
            .I(N__28992));
    InMux I__6323 (
            .O(N__29037),
            .I(N__28987));
    LocalMux I__6322 (
            .O(N__29034),
            .I(N__28984));
    LocalMux I__6321 (
            .O(N__29031),
            .I(N__28977));
    LocalMux I__6320 (
            .O(N__29028),
            .I(N__28977));
    Span4Mux_h I__6319 (
            .O(N__29025),
            .I(N__28977));
    LocalMux I__6318 (
            .O(N__29020),
            .I(N__28970));
    Span4Mux_h I__6317 (
            .O(N__29017),
            .I(N__28970));
    Span4Mux_v I__6316 (
            .O(N__29014),
            .I(N__28970));
    LocalMux I__6315 (
            .O(N__29007),
            .I(N__28961));
    Span4Mux_s0_h I__6314 (
            .O(N__29000),
            .I(N__28961));
    Span4Mux_s3_v I__6313 (
            .O(N__28997),
            .I(N__28961));
    LocalMux I__6312 (
            .O(N__28992),
            .I(N__28961));
    InMux I__6311 (
            .O(N__28991),
            .I(N__28956));
    InMux I__6310 (
            .O(N__28990),
            .I(N__28956));
    LocalMux I__6309 (
            .O(N__28987),
            .I(\POWERLED.count_clk_en ));
    Odrv12 I__6308 (
            .O(N__28984),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__6307 (
            .O(N__28977),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__6306 (
            .O(N__28970),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__6305 (
            .O(N__28961),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__6304 (
            .O(N__28956),
            .I(\POWERLED.count_clk_en ));
    CascadeMux I__6303 (
            .O(N__28943),
            .I(\POWERLED.count_clkZ0Z_13_cascade_ ));
    InMux I__6302 (
            .O(N__28940),
            .I(N__28934));
    InMux I__6301 (
            .O(N__28939),
            .I(N__28934));
    LocalMux I__6300 (
            .O(N__28934),
            .I(\POWERLED.count_clkZ0Z_12 ));
    InMux I__6299 (
            .O(N__28931),
            .I(N__28928));
    LocalMux I__6298 (
            .O(N__28928),
            .I(\POWERLED.un2_count_clk_17_0_o2_1_0 ));
    InMux I__6297 (
            .O(N__28925),
            .I(N__28920));
    InMux I__6296 (
            .O(N__28924),
            .I(N__28915));
    InMux I__6295 (
            .O(N__28923),
            .I(N__28915));
    LocalMux I__6294 (
            .O(N__28920),
            .I(N__28912));
    LocalMux I__6293 (
            .O(N__28915),
            .I(N__28909));
    Span4Mux_h I__6292 (
            .O(N__28912),
            .I(N__28905));
    Span4Mux_v I__6291 (
            .O(N__28909),
            .I(N__28902));
    InMux I__6290 (
            .O(N__28908),
            .I(N__28899));
    Odrv4 I__6289 (
            .O(N__28905),
            .I(\POWERLED.N_676 ));
    Odrv4 I__6288 (
            .O(N__28902),
            .I(\POWERLED.N_676 ));
    LocalMux I__6287 (
            .O(N__28899),
            .I(\POWERLED.N_676 ));
    InMux I__6286 (
            .O(N__28892),
            .I(N__28889));
    LocalMux I__6285 (
            .O(N__28889),
            .I(\POWERLED.N_492 ));
    CascadeMux I__6284 (
            .O(N__28886),
            .I(N__28882));
    InMux I__6283 (
            .O(N__28885),
            .I(N__28877));
    InMux I__6282 (
            .O(N__28882),
            .I(N__28877));
    LocalMux I__6281 (
            .O(N__28877),
            .I(\POWERLED.dutycycle_0_5 ));
    InMux I__6280 (
            .O(N__28874),
            .I(N__28868));
    InMux I__6279 (
            .O(N__28873),
            .I(N__28868));
    LocalMux I__6278 (
            .O(N__28868),
            .I(N__28865));
    Span4Mux_s2_h I__6277 (
            .O(N__28865),
            .I(N__28862));
    Odrv4 I__6276 (
            .O(N__28862),
            .I(\POWERLED.func_state_RNIS28SBZ0Z_1 ));
    CascadeMux I__6275 (
            .O(N__28859),
            .I(\POWERLED.dutycycleZ1Z_5_cascade_ ));
    CascadeMux I__6274 (
            .O(N__28856),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_5_cascade_ ));
    CascadeMux I__6273 (
            .O(N__28853),
            .I(\POWERLED.dutycycle_0_sqmuxa_i_i_a3_0_a2_0_cascade_ ));
    InMux I__6272 (
            .O(N__28850),
            .I(N__28836));
    InMux I__6271 (
            .O(N__28849),
            .I(N__28836));
    InMux I__6270 (
            .O(N__28848),
            .I(N__28833));
    InMux I__6269 (
            .O(N__28847),
            .I(N__28829));
    InMux I__6268 (
            .O(N__28846),
            .I(N__28824));
    InMux I__6267 (
            .O(N__28845),
            .I(N__28824));
    InMux I__6266 (
            .O(N__28844),
            .I(N__28817));
    InMux I__6265 (
            .O(N__28843),
            .I(N__28817));
    InMux I__6264 (
            .O(N__28842),
            .I(N__28817));
    InMux I__6263 (
            .O(N__28841),
            .I(N__28810));
    LocalMux I__6262 (
            .O(N__28836),
            .I(N__28805));
    LocalMux I__6261 (
            .O(N__28833),
            .I(N__28805));
    InMux I__6260 (
            .O(N__28832),
            .I(N__28802));
    LocalMux I__6259 (
            .O(N__28829),
            .I(N__28797));
    LocalMux I__6258 (
            .O(N__28824),
            .I(N__28792));
    LocalMux I__6257 (
            .O(N__28817),
            .I(N__28792));
    InMux I__6256 (
            .O(N__28816),
            .I(N__28787));
    InMux I__6255 (
            .O(N__28815),
            .I(N__28782));
    InMux I__6254 (
            .O(N__28814),
            .I(N__28782));
    InMux I__6253 (
            .O(N__28813),
            .I(N__28779));
    LocalMux I__6252 (
            .O(N__28810),
            .I(N__28772));
    Span4Mux_s3_h I__6251 (
            .O(N__28805),
            .I(N__28772));
    LocalMux I__6250 (
            .O(N__28802),
            .I(N__28772));
    InMux I__6249 (
            .O(N__28801),
            .I(N__28767));
    InMux I__6248 (
            .O(N__28800),
            .I(N__28767));
    Span4Mux_v I__6247 (
            .O(N__28797),
            .I(N__28762));
    Span4Mux_v I__6246 (
            .O(N__28792),
            .I(N__28762));
    InMux I__6245 (
            .O(N__28791),
            .I(N__28757));
    InMux I__6244 (
            .O(N__28790),
            .I(N__28757));
    LocalMux I__6243 (
            .O(N__28787),
            .I(N__28754));
    LocalMux I__6242 (
            .O(N__28782),
            .I(func_state_RNI_2_0));
    LocalMux I__6241 (
            .O(N__28779),
            .I(func_state_RNI_2_0));
    Odrv4 I__6240 (
            .O(N__28772),
            .I(func_state_RNI_2_0));
    LocalMux I__6239 (
            .O(N__28767),
            .I(func_state_RNI_2_0));
    Odrv4 I__6238 (
            .O(N__28762),
            .I(func_state_RNI_2_0));
    LocalMux I__6237 (
            .O(N__28757),
            .I(func_state_RNI_2_0));
    Odrv4 I__6236 (
            .O(N__28754),
            .I(func_state_RNI_2_0));
    InMux I__6235 (
            .O(N__28739),
            .I(N__28736));
    LocalMux I__6234 (
            .O(N__28736),
            .I(\POWERLED.un1_count_off_1_sqmuxa_8_ns_1 ));
    InMux I__6233 (
            .O(N__28733),
            .I(N__28730));
    LocalMux I__6232 (
            .O(N__28730),
            .I(\POWERLED.count_clk_0_0 ));
    InMux I__6231 (
            .O(N__28727),
            .I(N__28724));
    LocalMux I__6230 (
            .O(N__28724),
            .I(\POWERLED.count_clk_RNI_0Z0Z_0 ));
    InMux I__6229 (
            .O(N__28721),
            .I(N__28718));
    LocalMux I__6228 (
            .O(N__28718),
            .I(N__28711));
    InMux I__6227 (
            .O(N__28717),
            .I(N__28702));
    InMux I__6226 (
            .O(N__28716),
            .I(N__28702));
    InMux I__6225 (
            .O(N__28715),
            .I(N__28702));
    InMux I__6224 (
            .O(N__28714),
            .I(N__28702));
    Odrv4 I__6223 (
            .O(N__28711),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__6222 (
            .O(N__28702),
            .I(\POWERLED.count_clkZ0Z_0 ));
    InMux I__6221 (
            .O(N__28697),
            .I(N__28688));
    InMux I__6220 (
            .O(N__28696),
            .I(N__28688));
    InMux I__6219 (
            .O(N__28695),
            .I(N__28688));
    LocalMux I__6218 (
            .O(N__28688),
            .I(\POWERLED.count_clk_1_14 ));
    CascadeMux I__6217 (
            .O(N__28685),
            .I(\POWERLED.count_clkZ0Z_0_cascade_ ));
    InMux I__6216 (
            .O(N__28682),
            .I(N__28676));
    InMux I__6215 (
            .O(N__28681),
            .I(N__28676));
    LocalMux I__6214 (
            .O(N__28676),
            .I(\POWERLED.count_clkZ0Z_14 ));
    InMux I__6213 (
            .O(N__28673),
            .I(N__28669));
    InMux I__6212 (
            .O(N__28672),
            .I(N__28666));
    LocalMux I__6211 (
            .O(N__28669),
            .I(\POWERLED.count_clkZ0Z_11 ));
    LocalMux I__6210 (
            .O(N__28666),
            .I(\POWERLED.count_clkZ0Z_11 ));
    CascadeMux I__6209 (
            .O(N__28661),
            .I(\POWERLED.un2_count_clk_17_0_o2_1_1_cascade_ ));
    InMux I__6208 (
            .O(N__28658),
            .I(N__28655));
    LocalMux I__6207 (
            .O(N__28655),
            .I(\POWERLED.un2_count_clk_17_0_o2_1_2 ));
    CascadeMux I__6206 (
            .O(N__28652),
            .I(N__28649));
    InMux I__6205 (
            .O(N__28649),
            .I(N__28645));
    InMux I__6204 (
            .O(N__28648),
            .I(N__28642));
    LocalMux I__6203 (
            .O(N__28645),
            .I(\POWERLED.count_clk_RNISLCE7Z0Z_10 ));
    LocalMux I__6202 (
            .O(N__28642),
            .I(\POWERLED.count_clk_RNISLCE7Z0Z_10 ));
    CascadeMux I__6201 (
            .O(N__28637),
            .I(N__28634));
    InMux I__6200 (
            .O(N__28634),
            .I(N__28631));
    LocalMux I__6199 (
            .O(N__28631),
            .I(\POWERLED.count_clk_en_917_0 ));
    CascadeMux I__6198 (
            .O(N__28628),
            .I(N__28625));
    InMux I__6197 (
            .O(N__28625),
            .I(N__28618));
    InMux I__6196 (
            .O(N__28624),
            .I(N__28618));
    InMux I__6195 (
            .O(N__28623),
            .I(N__28615));
    LocalMux I__6194 (
            .O(N__28618),
            .I(N__28612));
    LocalMux I__6193 (
            .O(N__28615),
            .I(N__28609));
    Span4Mux_v I__6192 (
            .O(N__28612),
            .I(N__28604));
    Span4Mux_s3_h I__6191 (
            .O(N__28609),
            .I(N__28604));
    Odrv4 I__6190 (
            .O(N__28604),
            .I(\POWERLED.func_state_RNIBVNS_2Z0Z_0 ));
    CascadeMux I__6189 (
            .O(N__28601),
            .I(\POWERLED.count_clk_en_1_cascade_ ));
    InMux I__6188 (
            .O(N__28598),
            .I(N__28594));
    InMux I__6187 (
            .O(N__28597),
            .I(N__28591));
    LocalMux I__6186 (
            .O(N__28594),
            .I(N__28585));
    LocalMux I__6185 (
            .O(N__28591),
            .I(N__28585));
    InMux I__6184 (
            .O(N__28590),
            .I(N__28582));
    Span4Mux_s3_h I__6183 (
            .O(N__28585),
            .I(N__28579));
    LocalMux I__6182 (
            .O(N__28582),
            .I(\POWERLED.N_617 ));
    Odrv4 I__6181 (
            .O(N__28579),
            .I(\POWERLED.N_617 ));
    CascadeMux I__6180 (
            .O(N__28574),
            .I(\POWERLED.count_clk_en_cascade_ ));
    CascadeMux I__6179 (
            .O(N__28571),
            .I(N__28568));
    InMux I__6178 (
            .O(N__28568),
            .I(N__28565));
    LocalMux I__6177 (
            .O(N__28565),
            .I(N__28562));
    Odrv4 I__6176 (
            .O(N__28562),
            .I(\POWERLED.un1_count_clk_2_axb_12 ));
    InMux I__6175 (
            .O(N__28559),
            .I(\POWERLED.un1_count_clk_2_cry_12 ));
    InMux I__6174 (
            .O(N__28556),
            .I(\POWERLED.un1_count_clk_2_cry_13_cZ0 ));
    InMux I__6173 (
            .O(N__28553),
            .I(N__28533));
    InMux I__6172 (
            .O(N__28552),
            .I(N__28533));
    InMux I__6171 (
            .O(N__28551),
            .I(N__28533));
    InMux I__6170 (
            .O(N__28550),
            .I(N__28524));
    InMux I__6169 (
            .O(N__28549),
            .I(N__28524));
    InMux I__6168 (
            .O(N__28548),
            .I(N__28524));
    InMux I__6167 (
            .O(N__28547),
            .I(N__28524));
    CascadeMux I__6166 (
            .O(N__28546),
            .I(N__28517));
    InMux I__6165 (
            .O(N__28545),
            .I(N__28509));
    InMux I__6164 (
            .O(N__28544),
            .I(N__28509));
    InMux I__6163 (
            .O(N__28543),
            .I(N__28509));
    InMux I__6162 (
            .O(N__28542),
            .I(N__28502));
    InMux I__6161 (
            .O(N__28541),
            .I(N__28502));
    InMux I__6160 (
            .O(N__28540),
            .I(N__28502));
    LocalMux I__6159 (
            .O(N__28533),
            .I(N__28497));
    LocalMux I__6158 (
            .O(N__28524),
            .I(N__28497));
    InMux I__6157 (
            .O(N__28523),
            .I(N__28484));
    InMux I__6156 (
            .O(N__28522),
            .I(N__28484));
    InMux I__6155 (
            .O(N__28521),
            .I(N__28484));
    InMux I__6154 (
            .O(N__28520),
            .I(N__28484));
    InMux I__6153 (
            .O(N__28517),
            .I(N__28484));
    InMux I__6152 (
            .O(N__28516),
            .I(N__28484));
    LocalMux I__6151 (
            .O(N__28509),
            .I(\POWERLED.func_state_RNI2VV9A_0_0 ));
    LocalMux I__6150 (
            .O(N__28502),
            .I(\POWERLED.func_state_RNI2VV9A_0_0 ));
    Odrv4 I__6149 (
            .O(N__28497),
            .I(\POWERLED.func_state_RNI2VV9A_0_0 ));
    LocalMux I__6148 (
            .O(N__28484),
            .I(\POWERLED.func_state_RNI2VV9A_0_0 ));
    InMux I__6147 (
            .O(N__28475),
            .I(\POWERLED.un1_count_clk_2_cry_14 ));
    InMux I__6146 (
            .O(N__28472),
            .I(N__28469));
    LocalMux I__6145 (
            .O(N__28469),
            .I(N__28466));
    Odrv12 I__6144 (
            .O(N__28466),
            .I(\POWERLED.count_clk_0_15 ));
    InMux I__6143 (
            .O(N__28463),
            .I(N__28460));
    LocalMux I__6142 (
            .O(N__28460),
            .I(N__28456));
    InMux I__6141 (
            .O(N__28459),
            .I(N__28453));
    Odrv12 I__6140 (
            .O(N__28456),
            .I(\POWERLED.count_clk_1_15 ));
    LocalMux I__6139 (
            .O(N__28453),
            .I(\POWERLED.count_clk_1_15 ));
    InMux I__6138 (
            .O(N__28448),
            .I(N__28444));
    InMux I__6137 (
            .O(N__28447),
            .I(N__28441));
    LocalMux I__6136 (
            .O(N__28444),
            .I(\POWERLED.count_clkZ0Z_15 ));
    LocalMux I__6135 (
            .O(N__28441),
            .I(\POWERLED.count_clkZ0Z_15 ));
    InMux I__6134 (
            .O(N__28436),
            .I(N__28433));
    LocalMux I__6133 (
            .O(N__28433),
            .I(N__28430));
    Span4Mux_v I__6132 (
            .O(N__28430),
            .I(N__28425));
    InMux I__6131 (
            .O(N__28429),
            .I(N__28420));
    InMux I__6130 (
            .O(N__28428),
            .I(N__28420));
    Odrv4 I__6129 (
            .O(N__28425),
            .I(\POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ));
    LocalMux I__6128 (
            .O(N__28420),
            .I(\POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ));
    InMux I__6127 (
            .O(N__28415),
            .I(N__28409));
    InMux I__6126 (
            .O(N__28414),
            .I(N__28409));
    LocalMux I__6125 (
            .O(N__28409),
            .I(\POWERLED.count_clkZ0Z_10 ));
    InMux I__6124 (
            .O(N__28406),
            .I(N__28403));
    LocalMux I__6123 (
            .O(N__28403),
            .I(\POWERLED.un1_count_clk_2_axb_10 ));
    InMux I__6122 (
            .O(N__28400),
            .I(N__28397));
    LocalMux I__6121 (
            .O(N__28397),
            .I(\POWERLED.un1_count_clk_2_axb_14 ));
    InMux I__6120 (
            .O(N__28394),
            .I(N__28388));
    InMux I__6119 (
            .O(N__28393),
            .I(N__28388));
    LocalMux I__6118 (
            .O(N__28388),
            .I(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ));
    InMux I__6117 (
            .O(N__28385),
            .I(\POWERLED.un1_count_clk_2_cry_3 ));
    InMux I__6116 (
            .O(N__28382),
            .I(N__28378));
    CascadeMux I__6115 (
            .O(N__28381),
            .I(N__28374));
    LocalMux I__6114 (
            .O(N__28378),
            .I(N__28371));
    InMux I__6113 (
            .O(N__28377),
            .I(N__28368));
    InMux I__6112 (
            .O(N__28374),
            .I(N__28365));
    Odrv4 I__6111 (
            .O(N__28371),
            .I(\POWERLED.count_clkZ0Z_5 ));
    LocalMux I__6110 (
            .O(N__28368),
            .I(\POWERLED.count_clkZ0Z_5 ));
    LocalMux I__6109 (
            .O(N__28365),
            .I(\POWERLED.count_clkZ0Z_5 ));
    InMux I__6108 (
            .O(N__28358),
            .I(N__28352));
    InMux I__6107 (
            .O(N__28357),
            .I(N__28352));
    LocalMux I__6106 (
            .O(N__28352),
            .I(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ));
    InMux I__6105 (
            .O(N__28349),
            .I(\POWERLED.un1_count_clk_2_cry_4 ));
    InMux I__6104 (
            .O(N__28346),
            .I(N__28339));
    InMux I__6103 (
            .O(N__28345),
            .I(N__28339));
    InMux I__6102 (
            .O(N__28344),
            .I(N__28336));
    LocalMux I__6101 (
            .O(N__28339),
            .I(\POWERLED.count_clkZ0Z_6 ));
    LocalMux I__6100 (
            .O(N__28336),
            .I(\POWERLED.count_clkZ0Z_6 ));
    InMux I__6099 (
            .O(N__28331),
            .I(N__28325));
    InMux I__6098 (
            .O(N__28330),
            .I(N__28325));
    LocalMux I__6097 (
            .O(N__28325),
            .I(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ));
    InMux I__6096 (
            .O(N__28322),
            .I(\POWERLED.un1_count_clk_2_cry_5 ));
    InMux I__6095 (
            .O(N__28319),
            .I(N__28315));
    CascadeMux I__6094 (
            .O(N__28318),
            .I(N__28311));
    LocalMux I__6093 (
            .O(N__28315),
            .I(N__28307));
    InMux I__6092 (
            .O(N__28314),
            .I(N__28304));
    InMux I__6091 (
            .O(N__28311),
            .I(N__28301));
    InMux I__6090 (
            .O(N__28310),
            .I(N__28297));
    Span4Mux_s2_h I__6089 (
            .O(N__28307),
            .I(N__28294));
    LocalMux I__6088 (
            .O(N__28304),
            .I(N__28291));
    LocalMux I__6087 (
            .O(N__28301),
            .I(N__28288));
    InMux I__6086 (
            .O(N__28300),
            .I(N__28285));
    LocalMux I__6085 (
            .O(N__28297),
            .I(N__28282));
    Span4Mux_h I__6084 (
            .O(N__28294),
            .I(N__28277));
    Span4Mux_s2_h I__6083 (
            .O(N__28291),
            .I(N__28277));
    Span4Mux_s2_h I__6082 (
            .O(N__28288),
            .I(N__28274));
    LocalMux I__6081 (
            .O(N__28285),
            .I(\POWERLED.count_clkZ0Z_7 ));
    Odrv12 I__6080 (
            .O(N__28282),
            .I(\POWERLED.count_clkZ0Z_7 ));
    Odrv4 I__6079 (
            .O(N__28277),
            .I(\POWERLED.count_clkZ0Z_7 ));
    Odrv4 I__6078 (
            .O(N__28274),
            .I(\POWERLED.count_clkZ0Z_7 ));
    InMux I__6077 (
            .O(N__28265),
            .I(N__28259));
    InMux I__6076 (
            .O(N__28264),
            .I(N__28259));
    LocalMux I__6075 (
            .O(N__28259),
            .I(N__28256));
    Span4Mux_h I__6074 (
            .O(N__28256),
            .I(N__28253));
    Odrv4 I__6073 (
            .O(N__28253),
            .I(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ));
    InMux I__6072 (
            .O(N__28250),
            .I(\POWERLED.un1_count_clk_2_cry_6 ));
    InMux I__6071 (
            .O(N__28247),
            .I(N__28242));
    InMux I__6070 (
            .O(N__28246),
            .I(N__28237));
    InMux I__6069 (
            .O(N__28245),
            .I(N__28237));
    LocalMux I__6068 (
            .O(N__28242),
            .I(N__28234));
    LocalMux I__6067 (
            .O(N__28237),
            .I(\POWERLED.count_clkZ0Z_8 ));
    Odrv4 I__6066 (
            .O(N__28234),
            .I(\POWERLED.count_clkZ0Z_8 ));
    InMux I__6065 (
            .O(N__28229),
            .I(N__28223));
    InMux I__6064 (
            .O(N__28228),
            .I(N__28223));
    LocalMux I__6063 (
            .O(N__28223),
            .I(N__28220));
    Odrv4 I__6062 (
            .O(N__28220),
            .I(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ));
    InMux I__6061 (
            .O(N__28217),
            .I(\POWERLED.un1_count_clk_2_cry_7 ));
    InMux I__6060 (
            .O(N__28214),
            .I(N__28210));
    InMux I__6059 (
            .O(N__28213),
            .I(N__28206));
    LocalMux I__6058 (
            .O(N__28210),
            .I(N__28203));
    InMux I__6057 (
            .O(N__28209),
            .I(N__28200));
    LocalMux I__6056 (
            .O(N__28206),
            .I(N__28193));
    Span4Mux_v I__6055 (
            .O(N__28203),
            .I(N__28193));
    LocalMux I__6054 (
            .O(N__28200),
            .I(N__28193));
    Odrv4 I__6053 (
            .O(N__28193),
            .I(\POWERLED.count_clkZ0Z_9 ));
    InMux I__6052 (
            .O(N__28190),
            .I(N__28186));
    InMux I__6051 (
            .O(N__28189),
            .I(N__28183));
    LocalMux I__6050 (
            .O(N__28186),
            .I(N__28178));
    LocalMux I__6049 (
            .O(N__28183),
            .I(N__28178));
    Odrv4 I__6048 (
            .O(N__28178),
            .I(\POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ));
    InMux I__6047 (
            .O(N__28175),
            .I(bfn_12_6_0_));
    InMux I__6046 (
            .O(N__28172),
            .I(\POWERLED.un1_count_clk_2_cry_9 ));
    InMux I__6045 (
            .O(N__28169),
            .I(N__28163));
    InMux I__6044 (
            .O(N__28168),
            .I(N__28163));
    LocalMux I__6043 (
            .O(N__28163),
            .I(\POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ));
    InMux I__6042 (
            .O(N__28160),
            .I(\POWERLED.un1_count_clk_2_cry_10 ));
    InMux I__6041 (
            .O(N__28157),
            .I(\POWERLED.un1_count_clk_2_cry_11_cZ0 ));
    CascadeMux I__6040 (
            .O(N__28154),
            .I(\POWERLED.count_clkZ0Z_3_cascade_ ));
    CascadeMux I__6039 (
            .O(N__28151),
            .I(\POWERLED.un1_dutycycle_168_0_0_o2_4_cascade_ ));
    InMux I__6038 (
            .O(N__28148),
            .I(N__28142));
    InMux I__6037 (
            .O(N__28147),
            .I(N__28142));
    LocalMux I__6036 (
            .O(N__28142),
            .I(N__28139));
    Odrv4 I__6035 (
            .O(N__28139),
            .I(\POWERLED.count_clk_0_3 ));
    CascadeMux I__6034 (
            .O(N__28136),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_10_0_cascade_ ));
    InMux I__6033 (
            .O(N__28133),
            .I(N__28129));
    InMux I__6032 (
            .O(N__28132),
            .I(N__28126));
    LocalMux I__6031 (
            .O(N__28129),
            .I(N__28123));
    LocalMux I__6030 (
            .O(N__28126),
            .I(N__28120));
    Span4Mux_h I__6029 (
            .O(N__28123),
            .I(N__28117));
    Odrv4 I__6028 (
            .O(N__28120),
            .I(\POWERLED.N_625 ));
    Odrv4 I__6027 (
            .O(N__28117),
            .I(\POWERLED.N_625 ));
    InMux I__6026 (
            .O(N__28112),
            .I(N__28107));
    InMux I__6025 (
            .O(N__28111),
            .I(N__28102));
    InMux I__6024 (
            .O(N__28110),
            .I(N__28102));
    LocalMux I__6023 (
            .O(N__28107),
            .I(N__28099));
    LocalMux I__6022 (
            .O(N__28102),
            .I(N__28096));
    Odrv4 I__6021 (
            .O(N__28099),
            .I(\POWERLED.count_clk_RNIZ0Z_1 ));
    Odrv4 I__6020 (
            .O(N__28096),
            .I(\POWERLED.count_clk_RNIZ0Z_1 ));
    CascadeMux I__6019 (
            .O(N__28091),
            .I(\POWERLED.N_625_cascade_ ));
    InMux I__6018 (
            .O(N__28088),
            .I(N__28085));
    LocalMux I__6017 (
            .O(N__28085),
            .I(N__28082));
    Span4Mux_v I__6016 (
            .O(N__28082),
            .I(N__28079));
    Odrv4 I__6015 (
            .O(N__28079),
            .I(\POWERLED.count_clk_RNIPGQN2_5Z0Z_3 ));
    CascadeMux I__6014 (
            .O(N__28076),
            .I(N__28072));
    CascadeMux I__6013 (
            .O(N__28075),
            .I(N__28067));
    InMux I__6012 (
            .O(N__28072),
            .I(N__28064));
    InMux I__6011 (
            .O(N__28071),
            .I(N__28059));
    InMux I__6010 (
            .O(N__28070),
            .I(N__28059));
    InMux I__6009 (
            .O(N__28067),
            .I(N__28056));
    LocalMux I__6008 (
            .O(N__28064),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__6007 (
            .O(N__28059),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__6006 (
            .O(N__28056),
            .I(\POWERLED.count_clkZ0Z_1 ));
    CascadeMux I__6005 (
            .O(N__28049),
            .I(N__28046));
    InMux I__6004 (
            .O(N__28046),
            .I(N__28041));
    InMux I__6003 (
            .O(N__28045),
            .I(N__28036));
    InMux I__6002 (
            .O(N__28044),
            .I(N__28036));
    LocalMux I__6001 (
            .O(N__28041),
            .I(N__28033));
    LocalMux I__6000 (
            .O(N__28036),
            .I(\POWERLED.count_clkZ0Z_2 ));
    Odrv4 I__5999 (
            .O(N__28033),
            .I(\POWERLED.count_clkZ0Z_2 ));
    InMux I__5998 (
            .O(N__28028),
            .I(N__28022));
    InMux I__5997 (
            .O(N__28027),
            .I(N__28022));
    LocalMux I__5996 (
            .O(N__28022),
            .I(N__28019));
    Odrv4 I__5995 (
            .O(N__28019),
            .I(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ));
    InMux I__5994 (
            .O(N__28016),
            .I(\POWERLED.un1_count_clk_2_cry_1 ));
    CascadeMux I__5993 (
            .O(N__28013),
            .I(N__28010));
    InMux I__5992 (
            .O(N__28010),
            .I(N__28007));
    LocalMux I__5991 (
            .O(N__28007),
            .I(\POWERLED.count_clkZ0Z_3 ));
    InMux I__5990 (
            .O(N__28004),
            .I(N__27995));
    InMux I__5989 (
            .O(N__28003),
            .I(N__27995));
    InMux I__5988 (
            .O(N__28002),
            .I(N__27995));
    LocalMux I__5987 (
            .O(N__27995),
            .I(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ));
    InMux I__5986 (
            .O(N__27992),
            .I(\POWERLED.un1_count_clk_2_cry_2 ));
    CascadeMux I__5985 (
            .O(N__27989),
            .I(N__27984));
    InMux I__5984 (
            .O(N__27988),
            .I(N__27981));
    InMux I__5983 (
            .O(N__27987),
            .I(N__27978));
    InMux I__5982 (
            .O(N__27984),
            .I(N__27975));
    LocalMux I__5981 (
            .O(N__27981),
            .I(\POWERLED.count_clkZ0Z_4 ));
    LocalMux I__5980 (
            .O(N__27978),
            .I(\POWERLED.count_clkZ0Z_4 ));
    LocalMux I__5979 (
            .O(N__27975),
            .I(\POWERLED.count_clkZ0Z_4 ));
    InMux I__5978 (
            .O(N__27968),
            .I(N__27965));
    LocalMux I__5977 (
            .O(N__27965),
            .I(\POWERLED.N_529 ));
    InMux I__5976 (
            .O(N__27962),
            .I(N__27956));
    InMux I__5975 (
            .O(N__27961),
            .I(N__27956));
    LocalMux I__5974 (
            .O(N__27956),
            .I(N__27953));
    Odrv4 I__5973 (
            .O(N__27953),
            .I(\POWERLED.dutycycle_en_12 ));
    InMux I__5972 (
            .O(N__27950),
            .I(N__27947));
    LocalMux I__5971 (
            .O(N__27947),
            .I(\POWERLED.count_clk_0_8 ));
    InMux I__5970 (
            .O(N__27944),
            .I(N__27941));
    LocalMux I__5969 (
            .O(N__27941),
            .I(\POWERLED.count_clk_0_9 ));
    InMux I__5968 (
            .O(N__27938),
            .I(N__27935));
    LocalMux I__5967 (
            .O(N__27935),
            .I(\POWERLED.count_clk_0_2 ));
    InMux I__5966 (
            .O(N__27932),
            .I(N__27929));
    LocalMux I__5965 (
            .O(N__27929),
            .I(N__27926));
    Span4Mux_h I__5964 (
            .O(N__27926),
            .I(N__27923));
    Odrv4 I__5963 (
            .O(N__27923),
            .I(\POWERLED.un1_clk_100khz_40_and_i_0_a2_1_d ));
    CascadeMux I__5962 (
            .O(N__27920),
            .I(\POWERLED.N_526_cascade_ ));
    CascadeMux I__5961 (
            .O(N__27917),
            .I(N__27914));
    InMux I__5960 (
            .O(N__27914),
            .I(N__27908));
    InMux I__5959 (
            .O(N__27913),
            .I(N__27908));
    LocalMux I__5958 (
            .O(N__27908),
            .I(N__27905));
    Odrv12 I__5957 (
            .O(N__27905),
            .I(\POWERLED.dutycycle_RNI36306Z0Z_14 ));
    CascadeMux I__5956 (
            .O(N__27902),
            .I(N__27898));
    CascadeMux I__5955 (
            .O(N__27901),
            .I(N__27894));
    InMux I__5954 (
            .O(N__27898),
            .I(N__27886));
    InMux I__5953 (
            .O(N__27897),
            .I(N__27886));
    InMux I__5952 (
            .O(N__27894),
            .I(N__27881));
    InMux I__5951 (
            .O(N__27893),
            .I(N__27881));
    CascadeMux I__5950 (
            .O(N__27892),
            .I(N__27875));
    InMux I__5949 (
            .O(N__27891),
            .I(N__27872));
    LocalMux I__5948 (
            .O(N__27886),
            .I(N__27867));
    LocalMux I__5947 (
            .O(N__27881),
            .I(N__27867));
    InMux I__5946 (
            .O(N__27880),
            .I(N__27862));
    InMux I__5945 (
            .O(N__27879),
            .I(N__27862));
    InMux I__5944 (
            .O(N__27878),
            .I(N__27856));
    InMux I__5943 (
            .O(N__27875),
            .I(N__27856));
    LocalMux I__5942 (
            .O(N__27872),
            .I(N__27849));
    Span4Mux_s3_v I__5941 (
            .O(N__27867),
            .I(N__27849));
    LocalMux I__5940 (
            .O(N__27862),
            .I(N__27849));
    InMux I__5939 (
            .O(N__27861),
            .I(N__27846));
    LocalMux I__5938 (
            .O(N__27856),
            .I(N__27841));
    Span4Mux_v I__5937 (
            .O(N__27849),
            .I(N__27841));
    LocalMux I__5936 (
            .O(N__27846),
            .I(\POWERLED.func_state_RNI_8Z0Z_1 ));
    Odrv4 I__5935 (
            .O(N__27841),
            .I(\POWERLED.func_state_RNI_8Z0Z_1 ));
    InMux I__5934 (
            .O(N__27836),
            .I(N__27826));
    InMux I__5933 (
            .O(N__27835),
            .I(N__27826));
    InMux I__5932 (
            .O(N__27834),
            .I(N__27820));
    InMux I__5931 (
            .O(N__27833),
            .I(N__27820));
    InMux I__5930 (
            .O(N__27832),
            .I(N__27814));
    InMux I__5929 (
            .O(N__27831),
            .I(N__27814));
    LocalMux I__5928 (
            .O(N__27826),
            .I(N__27811));
    CascadeMux I__5927 (
            .O(N__27825),
            .I(N__27807));
    LocalMux I__5926 (
            .O(N__27820),
            .I(N__27804));
    InMux I__5925 (
            .O(N__27819),
            .I(N__27801));
    LocalMux I__5924 (
            .O(N__27814),
            .I(N__27798));
    Span4Mux_s2_v I__5923 (
            .O(N__27811),
            .I(N__27795));
    InMux I__5922 (
            .O(N__27810),
            .I(N__27792));
    InMux I__5921 (
            .O(N__27807),
            .I(N__27789));
    Span4Mux_h I__5920 (
            .O(N__27804),
            .I(N__27786));
    LocalMux I__5919 (
            .O(N__27801),
            .I(N__27779));
    Span4Mux_s2_v I__5918 (
            .O(N__27798),
            .I(N__27779));
    Span4Mux_h I__5917 (
            .O(N__27795),
            .I(N__27779));
    LocalMux I__5916 (
            .O(N__27792),
            .I(\POWERLED.N_203 ));
    LocalMux I__5915 (
            .O(N__27789),
            .I(\POWERLED.N_203 ));
    Odrv4 I__5914 (
            .O(N__27786),
            .I(\POWERLED.N_203 ));
    Odrv4 I__5913 (
            .O(N__27779),
            .I(\POWERLED.N_203 ));
    InMux I__5912 (
            .O(N__27770),
            .I(N__27764));
    InMux I__5911 (
            .O(N__27769),
            .I(N__27756));
    InMux I__5910 (
            .O(N__27768),
            .I(N__27756));
    InMux I__5909 (
            .O(N__27767),
            .I(N__27756));
    LocalMux I__5908 (
            .O(N__27764),
            .I(N__27751));
    CascadeMux I__5907 (
            .O(N__27763),
            .I(N__27748));
    LocalMux I__5906 (
            .O(N__27756),
            .I(N__27740));
    InMux I__5905 (
            .O(N__27755),
            .I(N__27737));
    InMux I__5904 (
            .O(N__27754),
            .I(N__27734));
    Span4Mux_s3_h I__5903 (
            .O(N__27751),
            .I(N__27731));
    InMux I__5902 (
            .O(N__27748),
            .I(N__27726));
    InMux I__5901 (
            .O(N__27747),
            .I(N__27726));
    InMux I__5900 (
            .O(N__27746),
            .I(N__27721));
    InMux I__5899 (
            .O(N__27745),
            .I(N__27721));
    InMux I__5898 (
            .O(N__27744),
            .I(N__27716));
    InMux I__5897 (
            .O(N__27743),
            .I(N__27716));
    Odrv4 I__5896 (
            .O(N__27740),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__5895 (
            .O(N__27737),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__5894 (
            .O(N__27734),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv4 I__5893 (
            .O(N__27731),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__5892 (
            .O(N__27726),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__5891 (
            .O(N__27721),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__5890 (
            .O(N__27716),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    CascadeMux I__5889 (
            .O(N__27701),
            .I(\POWERLED.N_524_cascade_ ));
    InMux I__5888 (
            .O(N__27698),
            .I(N__27695));
    LocalMux I__5887 (
            .O(N__27695),
            .I(\POWERLED.un1_clk_100khz_47_and_i_1 ));
    IoInMux I__5886 (
            .O(N__27692),
            .I(N__27689));
    LocalMux I__5885 (
            .O(N__27689),
            .I(N__27684));
    CascadeMux I__5884 (
            .O(N__27688),
            .I(N__27681));
    CascadeMux I__5883 (
            .O(N__27687),
            .I(N__27678));
    IoSpan4Mux I__5882 (
            .O(N__27684),
            .I(N__27674));
    InMux I__5881 (
            .O(N__27681),
            .I(N__27667));
    InMux I__5880 (
            .O(N__27678),
            .I(N__27667));
    InMux I__5879 (
            .O(N__27677),
            .I(N__27660));
    Span4Mux_s2_v I__5878 (
            .O(N__27674),
            .I(N__27657));
    InMux I__5877 (
            .O(N__27673),
            .I(N__27654));
    InMux I__5876 (
            .O(N__27672),
            .I(N__27651));
    LocalMux I__5875 (
            .O(N__27667),
            .I(N__27648));
    InMux I__5874 (
            .O(N__27666),
            .I(N__27645));
    CascadeMux I__5873 (
            .O(N__27665),
            .I(N__27641));
    CascadeMux I__5872 (
            .O(N__27664),
            .I(N__27637));
    CascadeMux I__5871 (
            .O(N__27663),
            .I(N__27634));
    LocalMux I__5870 (
            .O(N__27660),
            .I(N__27631));
    Span4Mux_h I__5869 (
            .O(N__27657),
            .I(N__27626));
    LocalMux I__5868 (
            .O(N__27654),
            .I(N__27626));
    LocalMux I__5867 (
            .O(N__27651),
            .I(N__27618));
    Span4Mux_v I__5866 (
            .O(N__27648),
            .I(N__27612));
    LocalMux I__5865 (
            .O(N__27645),
            .I(N__27612));
    InMux I__5864 (
            .O(N__27644),
            .I(N__27609));
    InMux I__5863 (
            .O(N__27641),
            .I(N__27600));
    InMux I__5862 (
            .O(N__27640),
            .I(N__27600));
    InMux I__5861 (
            .O(N__27637),
            .I(N__27600));
    InMux I__5860 (
            .O(N__27634),
            .I(N__27600));
    Span4Mux_s2_v I__5859 (
            .O(N__27631),
            .I(N__27595));
    Span4Mux_h I__5858 (
            .O(N__27626),
            .I(N__27595));
    InMux I__5857 (
            .O(N__27625),
            .I(N__27590));
    InMux I__5856 (
            .O(N__27624),
            .I(N__27590));
    InMux I__5855 (
            .O(N__27623),
            .I(N__27583));
    InMux I__5854 (
            .O(N__27622),
            .I(N__27583));
    InMux I__5853 (
            .O(N__27621),
            .I(N__27583));
    Span4Mux_v I__5852 (
            .O(N__27618),
            .I(N__27579));
    CascadeMux I__5851 (
            .O(N__27617),
            .I(N__27576));
    Span4Mux_v I__5850 (
            .O(N__27612),
            .I(N__27569));
    LocalMux I__5849 (
            .O(N__27609),
            .I(N__27569));
    LocalMux I__5848 (
            .O(N__27600),
            .I(N__27566));
    Span4Mux_v I__5847 (
            .O(N__27595),
            .I(N__27559));
    LocalMux I__5846 (
            .O(N__27590),
            .I(N__27559));
    LocalMux I__5845 (
            .O(N__27583),
            .I(N__27559));
    CascadeMux I__5844 (
            .O(N__27582),
            .I(N__27556));
    Span4Mux_v I__5843 (
            .O(N__27579),
            .I(N__27553));
    InMux I__5842 (
            .O(N__27576),
            .I(N__27546));
    InMux I__5841 (
            .O(N__27575),
            .I(N__27546));
    InMux I__5840 (
            .O(N__27574),
            .I(N__27546));
    Span4Mux_h I__5839 (
            .O(N__27569),
            .I(N__27543));
    Span4Mux_v I__5838 (
            .O(N__27566),
            .I(N__27538));
    Span4Mux_v I__5837 (
            .O(N__27559),
            .I(N__27538));
    InMux I__5836 (
            .O(N__27556),
            .I(N__27535));
    Odrv4 I__5835 (
            .O(N__27553),
            .I(rsmrstn));
    LocalMux I__5834 (
            .O(N__27546),
            .I(rsmrstn));
    Odrv4 I__5833 (
            .O(N__27543),
            .I(rsmrstn));
    Odrv4 I__5832 (
            .O(N__27538),
            .I(rsmrstn));
    LocalMux I__5831 (
            .O(N__27535),
            .I(rsmrstn));
    InMux I__5830 (
            .O(N__27524),
            .I(N__27521));
    LocalMux I__5829 (
            .O(N__27521),
            .I(N__27516));
    InMux I__5828 (
            .O(N__27520),
            .I(N__27513));
    CascadeMux I__5827 (
            .O(N__27519),
            .I(N__27507));
    Span4Mux_v I__5826 (
            .O(N__27516),
            .I(N__27503));
    LocalMux I__5825 (
            .O(N__27513),
            .I(N__27500));
    InMux I__5824 (
            .O(N__27512),
            .I(N__27497));
    InMux I__5823 (
            .O(N__27511),
            .I(N__27492));
    InMux I__5822 (
            .O(N__27510),
            .I(N__27492));
    InMux I__5821 (
            .O(N__27507),
            .I(N__27487));
    InMux I__5820 (
            .O(N__27506),
            .I(N__27487));
    Odrv4 I__5819 (
            .O(N__27503),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    Odrv12 I__5818 (
            .O(N__27500),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__5817 (
            .O(N__27497),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__5816 (
            .O(N__27492),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__5815 (
            .O(N__27487),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    CascadeMux I__5814 (
            .O(N__27476),
            .I(N__27472));
    InMux I__5813 (
            .O(N__27475),
            .I(N__27467));
    InMux I__5812 (
            .O(N__27472),
            .I(N__27467));
    LocalMux I__5811 (
            .O(N__27467),
            .I(N__27464));
    Odrv12 I__5810 (
            .O(N__27464),
            .I(\POWERLED.N_2381_i ));
    CascadeMux I__5809 (
            .O(N__27461),
            .I(N__27453));
    InMux I__5808 (
            .O(N__27460),
            .I(N__27446));
    InMux I__5807 (
            .O(N__27459),
            .I(N__27446));
    InMux I__5806 (
            .O(N__27458),
            .I(N__27443));
    CascadeMux I__5805 (
            .O(N__27457),
            .I(N__27439));
    InMux I__5804 (
            .O(N__27456),
            .I(N__27436));
    InMux I__5803 (
            .O(N__27453),
            .I(N__27431));
    InMux I__5802 (
            .O(N__27452),
            .I(N__27431));
    InMux I__5801 (
            .O(N__27451),
            .I(N__27428));
    LocalMux I__5800 (
            .O(N__27446),
            .I(N__27425));
    LocalMux I__5799 (
            .O(N__27443),
            .I(N__27422));
    InMux I__5798 (
            .O(N__27442),
            .I(N__27419));
    InMux I__5797 (
            .O(N__27439),
            .I(N__27416));
    LocalMux I__5796 (
            .O(N__27436),
            .I(N__27413));
    LocalMux I__5795 (
            .O(N__27431),
            .I(N__27410));
    LocalMux I__5794 (
            .O(N__27428),
            .I(N__27401));
    Span4Mux_v I__5793 (
            .O(N__27425),
            .I(N__27401));
    Span4Mux_v I__5792 (
            .O(N__27422),
            .I(N__27401));
    LocalMux I__5791 (
            .O(N__27419),
            .I(N__27401));
    LocalMux I__5790 (
            .O(N__27416),
            .I(N__27396));
    Span4Mux_s2_h I__5789 (
            .O(N__27413),
            .I(N__27396));
    Span4Mux_v I__5788 (
            .O(N__27410),
            .I(N__27391));
    Span4Mux_v I__5787 (
            .O(N__27401),
            .I(N__27391));
    Span4Mux_v I__5786 (
            .O(N__27396),
            .I(N__27388));
    Odrv4 I__5785 (
            .O(N__27391),
            .I(\POWERLED.N_91_1_N ));
    Odrv4 I__5784 (
            .O(N__27388),
            .I(\POWERLED.N_91_1_N ));
    CascadeMux I__5783 (
            .O(N__27383),
            .I(\POWERLED.N_527_cascade_ ));
    CascadeMux I__5782 (
            .O(N__27380),
            .I(\POWERLED.un1_clk_100khz_48_and_i_1_cascade_ ));
    CascadeMux I__5781 (
            .O(N__27377),
            .I(N__27365));
    CascadeMux I__5780 (
            .O(N__27376),
            .I(N__27361));
    CascadeMux I__5779 (
            .O(N__27375),
            .I(N__27356));
    InMux I__5778 (
            .O(N__27374),
            .I(N__27347));
    InMux I__5777 (
            .O(N__27373),
            .I(N__27347));
    InMux I__5776 (
            .O(N__27372),
            .I(N__27347));
    CascadeMux I__5775 (
            .O(N__27371),
            .I(N__27337));
    InMux I__5774 (
            .O(N__27370),
            .I(N__27328));
    InMux I__5773 (
            .O(N__27369),
            .I(N__27328));
    InMux I__5772 (
            .O(N__27368),
            .I(N__27328));
    InMux I__5771 (
            .O(N__27365),
            .I(N__27328));
    InMux I__5770 (
            .O(N__27364),
            .I(N__27325));
    InMux I__5769 (
            .O(N__27361),
            .I(N__27316));
    InMux I__5768 (
            .O(N__27360),
            .I(N__27316));
    InMux I__5767 (
            .O(N__27359),
            .I(N__27316));
    InMux I__5766 (
            .O(N__27356),
            .I(N__27316));
    InMux I__5765 (
            .O(N__27355),
            .I(N__27313));
    InMux I__5764 (
            .O(N__27354),
            .I(N__27310));
    LocalMux I__5763 (
            .O(N__27347),
            .I(N__27307));
    InMux I__5762 (
            .O(N__27346),
            .I(N__27302));
    InMux I__5761 (
            .O(N__27345),
            .I(N__27302));
    InMux I__5760 (
            .O(N__27344),
            .I(N__27299));
    InMux I__5759 (
            .O(N__27343),
            .I(N__27290));
    InMux I__5758 (
            .O(N__27342),
            .I(N__27290));
    InMux I__5757 (
            .O(N__27341),
            .I(N__27290));
    InMux I__5756 (
            .O(N__27340),
            .I(N__27290));
    InMux I__5755 (
            .O(N__27337),
            .I(N__27287));
    LocalMux I__5754 (
            .O(N__27328),
            .I(N__27280));
    LocalMux I__5753 (
            .O(N__27325),
            .I(N__27280));
    LocalMux I__5752 (
            .O(N__27316),
            .I(N__27280));
    LocalMux I__5751 (
            .O(N__27313),
            .I(N__27275));
    LocalMux I__5750 (
            .O(N__27310),
            .I(N__27275));
    Odrv12 I__5749 (
            .O(N__27307),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__5748 (
            .O(N__27302),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__5747 (
            .O(N__27299),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__5746 (
            .O(N__27290),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__5745 (
            .O(N__27287),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__5744 (
            .O(N__27280),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__5743 (
            .O(N__27275),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    CascadeMux I__5742 (
            .O(N__27260),
            .I(\POWERLED.un1_clk_100khz_30_and_i_0_a2_5_0_0_cascade_ ));
    InMux I__5741 (
            .O(N__27257),
            .I(N__27254));
    LocalMux I__5740 (
            .O(N__27254),
            .I(\POWERLED.dutycycle_eena_2_0_0_tz_1 ));
    CascadeMux I__5739 (
            .O(N__27251),
            .I(\POWERLED.dutycycle_eena_2_d_0_cascade_ ));
    InMux I__5738 (
            .O(N__27248),
            .I(N__27242));
    InMux I__5737 (
            .O(N__27247),
            .I(N__27242));
    LocalMux I__5736 (
            .O(N__27242),
            .I(N__27239));
    Odrv12 I__5735 (
            .O(N__27239),
            .I(\POWERLED.dutycycle_RNIRUFD6Z0Z_9 ));
    InMux I__5734 (
            .O(N__27236),
            .I(N__27229));
    InMux I__5733 (
            .O(N__27235),
            .I(N__27229));
    InMux I__5732 (
            .O(N__27234),
            .I(N__27224));
    LocalMux I__5731 (
            .O(N__27229),
            .I(N__27221));
    InMux I__5730 (
            .O(N__27228),
            .I(N__27216));
    InMux I__5729 (
            .O(N__27227),
            .I(N__27216));
    LocalMux I__5728 (
            .O(N__27224),
            .I(N__27213));
    Span4Mux_s3_v I__5727 (
            .O(N__27221),
            .I(N__27210));
    LocalMux I__5726 (
            .O(N__27216),
            .I(N__27207));
    Span4Mux_h I__5725 (
            .O(N__27213),
            .I(N__27202));
    Span4Mux_h I__5724 (
            .O(N__27210),
            .I(N__27197));
    Span4Mux_h I__5723 (
            .O(N__27207),
            .I(N__27197));
    InMux I__5722 (
            .O(N__27206),
            .I(N__27192));
    InMux I__5721 (
            .O(N__27205),
            .I(N__27192));
    Odrv4 I__5720 (
            .O(N__27202),
            .I(\POWERLED.func_state_RNI2MQDZ0Z_1 ));
    Odrv4 I__5719 (
            .O(N__27197),
            .I(\POWERLED.func_state_RNI2MQDZ0Z_1 ));
    LocalMux I__5718 (
            .O(N__27192),
            .I(\POWERLED.func_state_RNI2MQDZ0Z_1 ));
    CascadeMux I__5717 (
            .O(N__27185),
            .I(N__27181));
    InMux I__5716 (
            .O(N__27184),
            .I(N__27178));
    InMux I__5715 (
            .O(N__27181),
            .I(N__27168));
    LocalMux I__5714 (
            .O(N__27178),
            .I(N__27165));
    InMux I__5713 (
            .O(N__27177),
            .I(N__27160));
    InMux I__5712 (
            .O(N__27176),
            .I(N__27160));
    InMux I__5711 (
            .O(N__27175),
            .I(N__27157));
    InMux I__5710 (
            .O(N__27174),
            .I(N__27152));
    InMux I__5709 (
            .O(N__27173),
            .I(N__27152));
    InMux I__5708 (
            .O(N__27172),
            .I(N__27146));
    InMux I__5707 (
            .O(N__27171),
            .I(N__27146));
    LocalMux I__5706 (
            .O(N__27168),
            .I(N__27141));
    Span4Mux_v I__5705 (
            .O(N__27165),
            .I(N__27141));
    LocalMux I__5704 (
            .O(N__27160),
            .I(N__27138));
    LocalMux I__5703 (
            .O(N__27157),
            .I(N__27133));
    LocalMux I__5702 (
            .O(N__27152),
            .I(N__27133));
    CascadeMux I__5701 (
            .O(N__27151),
            .I(N__27130));
    LocalMux I__5700 (
            .O(N__27146),
            .I(N__27127));
    Span4Mux_h I__5699 (
            .O(N__27141),
            .I(N__27122));
    Span4Mux_h I__5698 (
            .O(N__27138),
            .I(N__27122));
    Span4Mux_h I__5697 (
            .O(N__27133),
            .I(N__27119));
    InMux I__5696 (
            .O(N__27130),
            .I(N__27116));
    Odrv4 I__5695 (
            .O(N__27127),
            .I(RSMRSTn_rep1));
    Odrv4 I__5694 (
            .O(N__27122),
            .I(RSMRSTn_rep1));
    Odrv4 I__5693 (
            .O(N__27119),
            .I(RSMRSTn_rep1));
    LocalMux I__5692 (
            .O(N__27116),
            .I(RSMRSTn_rep1));
    CascadeMux I__5691 (
            .O(N__27107),
            .I(N__27100));
    CascadeMux I__5690 (
            .O(N__27106),
            .I(N__27093));
    CascadeMux I__5689 (
            .O(N__27105),
            .I(N__27090));
    CascadeMux I__5688 (
            .O(N__27104),
            .I(N__27086));
    InMux I__5687 (
            .O(N__27103),
            .I(N__27082));
    InMux I__5686 (
            .O(N__27100),
            .I(N__27079));
    InMux I__5685 (
            .O(N__27099),
            .I(N__27076));
    CascadeMux I__5684 (
            .O(N__27098),
            .I(N__27070));
    CascadeMux I__5683 (
            .O(N__27097),
            .I(N__27067));
    InMux I__5682 (
            .O(N__27096),
            .I(N__27058));
    InMux I__5681 (
            .O(N__27093),
            .I(N__27058));
    InMux I__5680 (
            .O(N__27090),
            .I(N__27058));
    InMux I__5679 (
            .O(N__27089),
            .I(N__27051));
    InMux I__5678 (
            .O(N__27086),
            .I(N__27051));
    InMux I__5677 (
            .O(N__27085),
            .I(N__27051));
    LocalMux I__5676 (
            .O(N__27082),
            .I(N__27046));
    LocalMux I__5675 (
            .O(N__27079),
            .I(N__27046));
    LocalMux I__5674 (
            .O(N__27076),
            .I(N__27043));
    InMux I__5673 (
            .O(N__27075),
            .I(N__27040));
    InMux I__5672 (
            .O(N__27074),
            .I(N__27033));
    InMux I__5671 (
            .O(N__27073),
            .I(N__27033));
    InMux I__5670 (
            .O(N__27070),
            .I(N__27033));
    InMux I__5669 (
            .O(N__27067),
            .I(N__27028));
    InMux I__5668 (
            .O(N__27066),
            .I(N__27028));
    InMux I__5667 (
            .O(N__27065),
            .I(N__27025));
    LocalMux I__5666 (
            .O(N__27058),
            .I(N__27020));
    LocalMux I__5665 (
            .O(N__27051),
            .I(N__27020));
    Span4Mux_v I__5664 (
            .O(N__27046),
            .I(N__27015));
    Span4Mux_v I__5663 (
            .O(N__27043),
            .I(N__27015));
    LocalMux I__5662 (
            .O(N__27040),
            .I(N__27004));
    LocalMux I__5661 (
            .O(N__27033),
            .I(N__27004));
    LocalMux I__5660 (
            .O(N__27028),
            .I(N__27004));
    LocalMux I__5659 (
            .O(N__27025),
            .I(N__27004));
    Span4Mux_s3_v I__5658 (
            .O(N__27020),
            .I(N__27004));
    Odrv4 I__5657 (
            .O(N__27015),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv4 I__5656 (
            .O(N__27004),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    CascadeMux I__5655 (
            .O(N__26999),
            .I(\POWERLED.N_520_cascade_ ));
    CascadeMux I__5654 (
            .O(N__26996),
            .I(N__26993));
    InMux I__5653 (
            .O(N__26993),
            .I(N__26989));
    InMux I__5652 (
            .O(N__26992),
            .I(N__26986));
    LocalMux I__5651 (
            .O(N__26989),
            .I(N__26981));
    LocalMux I__5650 (
            .O(N__26986),
            .I(N__26981));
    Odrv4 I__5649 (
            .O(N__26981),
            .I(\POWERLED.dutycycle_RNIRUFD6Z0Z_12 ));
    InMux I__5648 (
            .O(N__26978),
            .I(N__26970));
    CascadeMux I__5647 (
            .O(N__26977),
            .I(N__26964));
    InMux I__5646 (
            .O(N__26976),
            .I(N__26956));
    InMux I__5645 (
            .O(N__26975),
            .I(N__26956));
    InMux I__5644 (
            .O(N__26974),
            .I(N__26956));
    InMux I__5643 (
            .O(N__26973),
            .I(N__26953));
    LocalMux I__5642 (
            .O(N__26970),
            .I(N__26949));
    InMux I__5641 (
            .O(N__26969),
            .I(N__26942));
    InMux I__5640 (
            .O(N__26968),
            .I(N__26942));
    InMux I__5639 (
            .O(N__26967),
            .I(N__26942));
    InMux I__5638 (
            .O(N__26964),
            .I(N__26939));
    InMux I__5637 (
            .O(N__26963),
            .I(N__26936));
    LocalMux I__5636 (
            .O(N__26956),
            .I(N__26931));
    LocalMux I__5635 (
            .O(N__26953),
            .I(N__26931));
    InMux I__5634 (
            .O(N__26952),
            .I(N__26928));
    Span4Mux_h I__5633 (
            .O(N__26949),
            .I(N__26923));
    LocalMux I__5632 (
            .O(N__26942),
            .I(N__26923));
    LocalMux I__5631 (
            .O(N__26939),
            .I(N__26920));
    LocalMux I__5630 (
            .O(N__26936),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv12 I__5629 (
            .O(N__26931),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__5628 (
            .O(N__26928),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__5627 (
            .O(N__26923),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__5626 (
            .O(N__26920),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    CascadeMux I__5625 (
            .O(N__26909),
            .I(\POWERLED.N_518_cascade_ ));
    InMux I__5624 (
            .O(N__26906),
            .I(N__26903));
    LocalMux I__5623 (
            .O(N__26903),
            .I(\POWERLED.un1_clk_100khz_42_and_i_1 ));
    InMux I__5622 (
            .O(N__26900),
            .I(N__26897));
    LocalMux I__5621 (
            .O(N__26897),
            .I(N__26894));
    Span4Mux_h I__5620 (
            .O(N__26894),
            .I(N__26891));
    Odrv4 I__5619 (
            .O(N__26891),
            .I(\POWERLED.un1_clk_100khz_40_and_i_0_a2_1_0_3_1 ));
    CascadeMux I__5618 (
            .O(N__26888),
            .I(\POWERLED.N_203_cascade_ ));
    CascadeMux I__5617 (
            .O(N__26885),
            .I(\POWERLED.N_521_cascade_ ));
    CascadeMux I__5616 (
            .O(N__26882),
            .I(\POWERLED.un1_clk_100khz_43_and_i_1_cascade_ ));
    InMux I__5615 (
            .O(N__26879),
            .I(N__26876));
    LocalMux I__5614 (
            .O(N__26876),
            .I(\POWERLED.N_523 ));
    CascadeMux I__5613 (
            .O(N__26873),
            .I(\POWERLED.N_503_cascade_ ));
    InMux I__5612 (
            .O(N__26870),
            .I(N__26864));
    InMux I__5611 (
            .O(N__26869),
            .I(N__26864));
    LocalMux I__5610 (
            .O(N__26864),
            .I(N__26861));
    Odrv12 I__5609 (
            .O(N__26861),
            .I(\POWERLED.dutycycle_1_0_0 ));
    InMux I__5608 (
            .O(N__26858),
            .I(N__26855));
    LocalMux I__5607 (
            .O(N__26855),
            .I(\POWERLED.dutycycle_eena ));
    InMux I__5606 (
            .O(N__26852),
            .I(N__26846));
    InMux I__5605 (
            .O(N__26851),
            .I(N__26846));
    LocalMux I__5604 (
            .O(N__26846),
            .I(\POWERLED.dutycycleZ1Z_0 ));
    InMux I__5603 (
            .O(N__26843),
            .I(N__26840));
    LocalMux I__5602 (
            .O(N__26840),
            .I(N__26837));
    Span4Mux_h I__5601 (
            .O(N__26837),
            .I(N__26834));
    Odrv4 I__5600 (
            .O(N__26834),
            .I(\POWERLED.N_510 ));
    CascadeMux I__5599 (
            .O(N__26831),
            .I(\POWERLED.un1_clk_100khz_36_and_i_0_a2_c_cascade_ ));
    InMux I__5598 (
            .O(N__26828),
            .I(N__26825));
    LocalMux I__5597 (
            .O(N__26825),
            .I(N__26817));
    InMux I__5596 (
            .O(N__26824),
            .I(N__26806));
    InMux I__5595 (
            .O(N__26823),
            .I(N__26806));
    InMux I__5594 (
            .O(N__26822),
            .I(N__26806));
    InMux I__5593 (
            .O(N__26821),
            .I(N__26806));
    InMux I__5592 (
            .O(N__26820),
            .I(N__26806));
    Span12Mux_s10_v I__5591 (
            .O(N__26817),
            .I(N__26799));
    LocalMux I__5590 (
            .O(N__26806),
            .I(N__26799));
    InMux I__5589 (
            .O(N__26805),
            .I(N__26796));
    InMux I__5588 (
            .O(N__26804),
            .I(N__26793));
    Odrv12 I__5587 (
            .O(N__26799),
            .I(rsmrst_pwrgd_signal));
    LocalMux I__5586 (
            .O(N__26796),
            .I(rsmrst_pwrgd_signal));
    LocalMux I__5585 (
            .O(N__26793),
            .I(rsmrst_pwrgd_signal));
    InMux I__5584 (
            .O(N__26786),
            .I(N__26783));
    LocalMux I__5583 (
            .O(N__26783),
            .I(\POWERLED.un1_clk_100khz_36_and_i_0_a2_d ));
    InMux I__5582 (
            .O(N__26780),
            .I(N__26777));
    LocalMux I__5581 (
            .O(N__26777),
            .I(\POWERLED.un1_clk_100khz_36_and_i_0_a2_1_0_2 ));
    CascadeMux I__5580 (
            .O(N__26774),
            .I(\POWERLED.un1_clk_100khz_36_and_i_0_a2_1_d_cascade_ ));
    InMux I__5579 (
            .O(N__26771),
            .I(N__26765));
    InMux I__5578 (
            .O(N__26770),
            .I(N__26765));
    LocalMux I__5577 (
            .O(N__26765),
            .I(N__26762));
    Span4Mux_h I__5576 (
            .O(N__26762),
            .I(N__26759));
    Odrv4 I__5575 (
            .O(N__26759),
            .I(\POWERLED.dutycycle_eena_5 ));
    CascadeMux I__5574 (
            .O(N__26756),
            .I(N__26749));
    InMux I__5573 (
            .O(N__26755),
            .I(N__26739));
    CascadeMux I__5572 (
            .O(N__26754),
            .I(N__26736));
    InMux I__5571 (
            .O(N__26753),
            .I(N__26731));
    InMux I__5570 (
            .O(N__26752),
            .I(N__26728));
    InMux I__5569 (
            .O(N__26749),
            .I(N__26721));
    InMux I__5568 (
            .O(N__26748),
            .I(N__26721));
    InMux I__5567 (
            .O(N__26747),
            .I(N__26721));
    InMux I__5566 (
            .O(N__26746),
            .I(N__26718));
    InMux I__5565 (
            .O(N__26745),
            .I(N__26715));
    InMux I__5564 (
            .O(N__26744),
            .I(N__26710));
    InMux I__5563 (
            .O(N__26743),
            .I(N__26710));
    InMux I__5562 (
            .O(N__26742),
            .I(N__26704));
    LocalMux I__5561 (
            .O(N__26739),
            .I(N__26701));
    InMux I__5560 (
            .O(N__26736),
            .I(N__26694));
    InMux I__5559 (
            .O(N__26735),
            .I(N__26694));
    InMux I__5558 (
            .O(N__26734),
            .I(N__26694));
    LocalMux I__5557 (
            .O(N__26731),
            .I(N__26691));
    LocalMux I__5556 (
            .O(N__26728),
            .I(N__26682));
    LocalMux I__5555 (
            .O(N__26721),
            .I(N__26682));
    LocalMux I__5554 (
            .O(N__26718),
            .I(N__26682));
    LocalMux I__5553 (
            .O(N__26715),
            .I(N__26682));
    LocalMux I__5552 (
            .O(N__26710),
            .I(N__26679));
    InMux I__5551 (
            .O(N__26709),
            .I(N__26676));
    InMux I__5550 (
            .O(N__26708),
            .I(N__26671));
    InMux I__5549 (
            .O(N__26707),
            .I(N__26671));
    LocalMux I__5548 (
            .O(N__26704),
            .I(N__26668));
    Span4Mux_v I__5547 (
            .O(N__26701),
            .I(N__26663));
    LocalMux I__5546 (
            .O(N__26694),
            .I(N__26663));
    Span4Mux_v I__5545 (
            .O(N__26691),
            .I(N__26658));
    Span4Mux_v I__5544 (
            .O(N__26682),
            .I(N__26658));
    Span4Mux_v I__5543 (
            .O(N__26679),
            .I(N__26651));
    LocalMux I__5542 (
            .O(N__26676),
            .I(N__26651));
    LocalMux I__5541 (
            .O(N__26671),
            .I(N__26651));
    Span12Mux_v I__5540 (
            .O(N__26668),
            .I(N__26648));
    Span4Mux_v I__5539 (
            .O(N__26663),
            .I(N__26645));
    Span4Mux_h I__5538 (
            .O(N__26658),
            .I(N__26640));
    Span4Mux_v I__5537 (
            .O(N__26651),
            .I(N__26640));
    Odrv12 I__5536 (
            .O(N__26648),
            .I(gpio_fpga_soc_4));
    Odrv4 I__5535 (
            .O(N__26645),
            .I(gpio_fpga_soc_4));
    Odrv4 I__5534 (
            .O(N__26640),
            .I(gpio_fpga_soc_4));
    CascadeMux I__5533 (
            .O(N__26633),
            .I(\POWERLED.N_249_cascade_ ));
    CascadeMux I__5532 (
            .O(N__26630),
            .I(\POWERLED.N_546_cascade_ ));
    InMux I__5531 (
            .O(N__26627),
            .I(N__26624));
    LocalMux I__5530 (
            .O(N__26624),
            .I(N__26620));
    InMux I__5529 (
            .O(N__26623),
            .I(N__26617));
    Span4Mux_h I__5528 (
            .O(N__26620),
            .I(N__26614));
    LocalMux I__5527 (
            .O(N__26617),
            .I(N__26611));
    Odrv4 I__5526 (
            .O(N__26614),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_0 ));
    Odrv12 I__5525 (
            .O(N__26611),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_0 ));
    InMux I__5524 (
            .O(N__26606),
            .I(N__26603));
    LocalMux I__5523 (
            .O(N__26603),
            .I(\POWERLED.N_482 ));
    InMux I__5522 (
            .O(N__26600),
            .I(N__26597));
    LocalMux I__5521 (
            .O(N__26597),
            .I(N__26594));
    Odrv12 I__5520 (
            .O(N__26594),
            .I(\POWERLED.g0_i_m2_rn_1_0 ));
    CascadeMux I__5519 (
            .O(N__26591),
            .I(\POWERLED.dutycycleZ0Z_1_cascade_ ));
    CascadeMux I__5518 (
            .O(N__26588),
            .I(N__26585));
    InMux I__5517 (
            .O(N__26585),
            .I(N__26582));
    LocalMux I__5516 (
            .O(N__26582),
            .I(\POWERLED.dutycycle_eena_0_0 ));
    InMux I__5515 (
            .O(N__26579),
            .I(N__26575));
    InMux I__5514 (
            .O(N__26578),
            .I(N__26572));
    LocalMux I__5513 (
            .O(N__26575),
            .I(N__26569));
    LocalMux I__5512 (
            .O(N__26572),
            .I(\POWERLED.g0_1 ));
    Odrv4 I__5511 (
            .O(N__26569),
            .I(\POWERLED.g0_1 ));
    CascadeMux I__5510 (
            .O(N__26564),
            .I(\POWERLED.dutycycle_eena_0_0_cascade_ ));
    CascadeMux I__5509 (
            .O(N__26561),
            .I(\POWERLED.dutycycle_eena_cascade_ ));
    InMux I__5508 (
            .O(N__26558),
            .I(N__26554));
    CascadeMux I__5507 (
            .O(N__26557),
            .I(N__26549));
    LocalMux I__5506 (
            .O(N__26554),
            .I(N__26544));
    InMux I__5505 (
            .O(N__26553),
            .I(N__26541));
    InMux I__5504 (
            .O(N__26552),
            .I(N__26537));
    InMux I__5503 (
            .O(N__26549),
            .I(N__26532));
    InMux I__5502 (
            .O(N__26548),
            .I(N__26532));
    CascadeMux I__5501 (
            .O(N__26547),
            .I(N__26529));
    Span4Mux_h I__5500 (
            .O(N__26544),
            .I(N__26526));
    LocalMux I__5499 (
            .O(N__26541),
            .I(N__26523));
    InMux I__5498 (
            .O(N__26540),
            .I(N__26519));
    LocalMux I__5497 (
            .O(N__26537),
            .I(N__26516));
    LocalMux I__5496 (
            .O(N__26532),
            .I(N__26513));
    InMux I__5495 (
            .O(N__26529),
            .I(N__26510));
    Span4Mux_h I__5494 (
            .O(N__26526),
            .I(N__26505));
    Span4Mux_h I__5493 (
            .O(N__26523),
            .I(N__26502));
    InMux I__5492 (
            .O(N__26522),
            .I(N__26499));
    LocalMux I__5491 (
            .O(N__26519),
            .I(N__26496));
    Span4Mux_v I__5490 (
            .O(N__26516),
            .I(N__26489));
    Span4Mux_v I__5489 (
            .O(N__26513),
            .I(N__26489));
    LocalMux I__5488 (
            .O(N__26510),
            .I(N__26489));
    InMux I__5487 (
            .O(N__26509),
            .I(N__26484));
    InMux I__5486 (
            .O(N__26508),
            .I(N__26484));
    Odrv4 I__5485 (
            .O(N__26505),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__5484 (
            .O(N__26502),
            .I(\POWERLED.dutycycle ));
    LocalMux I__5483 (
            .O(N__26499),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__5482 (
            .O(N__26496),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__5481 (
            .O(N__26489),
            .I(\POWERLED.dutycycle ));
    LocalMux I__5480 (
            .O(N__26484),
            .I(\POWERLED.dutycycle ));
    CascadeMux I__5479 (
            .O(N__26471),
            .I(N__26467));
    InMux I__5478 (
            .O(N__26470),
            .I(N__26462));
    InMux I__5477 (
            .O(N__26467),
            .I(N__26462));
    LocalMux I__5476 (
            .O(N__26462),
            .I(\POWERLED.g0_i_m2_sn ));
    CascadeMux I__5475 (
            .O(N__26459),
            .I(N__26450));
    CascadeMux I__5474 (
            .O(N__26458),
            .I(N__26447));
    InMux I__5473 (
            .O(N__26457),
            .I(N__26441));
    InMux I__5472 (
            .O(N__26456),
            .I(N__26441));
    InMux I__5471 (
            .O(N__26455),
            .I(N__26436));
    InMux I__5470 (
            .O(N__26454),
            .I(N__26436));
    InMux I__5469 (
            .O(N__26453),
            .I(N__26431));
    InMux I__5468 (
            .O(N__26450),
            .I(N__26431));
    InMux I__5467 (
            .O(N__26447),
            .I(N__26426));
    InMux I__5466 (
            .O(N__26446),
            .I(N__26426));
    LocalMux I__5465 (
            .O(N__26441),
            .I(N__26416));
    LocalMux I__5464 (
            .O(N__26436),
            .I(N__26416));
    LocalMux I__5463 (
            .O(N__26431),
            .I(N__26416));
    LocalMux I__5462 (
            .O(N__26426),
            .I(N__26416));
    InMux I__5461 (
            .O(N__26425),
            .I(N__26413));
    Span4Mux_v I__5460 (
            .O(N__26416),
            .I(N__26410));
    LocalMux I__5459 (
            .O(N__26413),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv4 I__5458 (
            .O(N__26410),
            .I(\POWERLED.func_stateZ0Z_0 ));
    InMux I__5457 (
            .O(N__26405),
            .I(N__26399));
    InMux I__5456 (
            .O(N__26404),
            .I(N__26399));
    LocalMux I__5455 (
            .O(N__26399),
            .I(\POWERLED.g0_i_m2_rn_1 ));
    InMux I__5454 (
            .O(N__26396),
            .I(N__26393));
    LocalMux I__5453 (
            .O(N__26393),
            .I(\POWERLED.dutycycleZ1Z_1 ));
    CascadeMux I__5452 (
            .O(N__26390),
            .I(N__26387));
    InMux I__5451 (
            .O(N__26387),
            .I(N__26380));
    InMux I__5450 (
            .O(N__26386),
            .I(N__26377));
    InMux I__5449 (
            .O(N__26385),
            .I(N__26372));
    InMux I__5448 (
            .O(N__26384),
            .I(N__26372));
    CascadeMux I__5447 (
            .O(N__26383),
            .I(N__26368));
    LocalMux I__5446 (
            .O(N__26380),
            .I(N__26358));
    LocalMux I__5445 (
            .O(N__26377),
            .I(N__26358));
    LocalMux I__5444 (
            .O(N__26372),
            .I(N__26358));
    InMux I__5443 (
            .O(N__26371),
            .I(N__26353));
    InMux I__5442 (
            .O(N__26368),
            .I(N__26353));
    InMux I__5441 (
            .O(N__26367),
            .I(N__26350));
    InMux I__5440 (
            .O(N__26366),
            .I(N__26346));
    CascadeMux I__5439 (
            .O(N__26365),
            .I(N__26343));
    Span4Mux_v I__5438 (
            .O(N__26358),
            .I(N__26339));
    LocalMux I__5437 (
            .O(N__26353),
            .I(N__26334));
    LocalMux I__5436 (
            .O(N__26350),
            .I(N__26334));
    InMux I__5435 (
            .O(N__26349),
            .I(N__26331));
    LocalMux I__5434 (
            .O(N__26346),
            .I(N__26328));
    InMux I__5433 (
            .O(N__26343),
            .I(N__26325));
    InMux I__5432 (
            .O(N__26342),
            .I(N__26322));
    Odrv4 I__5431 (
            .O(N__26339),
            .I(N_247));
    Odrv4 I__5430 (
            .O(N__26334),
            .I(N_247));
    LocalMux I__5429 (
            .O(N__26331),
            .I(N_247));
    Odrv4 I__5428 (
            .O(N__26328),
            .I(N_247));
    LocalMux I__5427 (
            .O(N__26325),
            .I(N_247));
    LocalMux I__5426 (
            .O(N__26322),
            .I(N_247));
    InMux I__5425 (
            .O(N__26309),
            .I(N__26306));
    LocalMux I__5424 (
            .O(N__26306),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_2 ));
    CascadeMux I__5423 (
            .O(N__26303),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_1_cascade_ ));
    InMux I__5422 (
            .O(N__26300),
            .I(N__26297));
    LocalMux I__5421 (
            .O(N__26297),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_4 ));
    InMux I__5420 (
            .O(N__26294),
            .I(N__26288));
    InMux I__5419 (
            .O(N__26293),
            .I(N__26288));
    LocalMux I__5418 (
            .O(N__26288),
            .I(\POWERLED.func_state_RNI_0Z0Z_1 ));
    InMux I__5417 (
            .O(N__26285),
            .I(N__26282));
    LocalMux I__5416 (
            .O(N__26282),
            .I(N__26277));
    InMux I__5415 (
            .O(N__26281),
            .I(N__26272));
    InMux I__5414 (
            .O(N__26280),
            .I(N__26269));
    Span4Mux_v I__5413 (
            .O(N__26277),
            .I(N__26266));
    InMux I__5412 (
            .O(N__26276),
            .I(N__26261));
    InMux I__5411 (
            .O(N__26275),
            .I(N__26261));
    LocalMux I__5410 (
            .O(N__26272),
            .I(N__26256));
    LocalMux I__5409 (
            .O(N__26269),
            .I(N__26256));
    Span4Mux_v I__5408 (
            .O(N__26266),
            .I(N__26253));
    LocalMux I__5407 (
            .O(N__26261),
            .I(N__26250));
    Span4Mux_h I__5406 (
            .O(N__26256),
            .I(N__26247));
    Odrv4 I__5405 (
            .O(N__26253),
            .I(func_state_RNI_4_1));
    Odrv4 I__5404 (
            .O(N__26250),
            .I(func_state_RNI_4_1));
    Odrv4 I__5403 (
            .O(N__26247),
            .I(func_state_RNI_4_1));
    InMux I__5402 (
            .O(N__26240),
            .I(N__26236));
    CascadeMux I__5401 (
            .O(N__26239),
            .I(N__26232));
    LocalMux I__5400 (
            .O(N__26236),
            .I(N__26227));
    InMux I__5399 (
            .O(N__26235),
            .I(N__26224));
    InMux I__5398 (
            .O(N__26232),
            .I(N__26219));
    InMux I__5397 (
            .O(N__26231),
            .I(N__26219));
    InMux I__5396 (
            .O(N__26230),
            .I(N__26216));
    Span4Mux_h I__5395 (
            .O(N__26227),
            .I(N__26213));
    LocalMux I__5394 (
            .O(N__26224),
            .I(N__26210));
    LocalMux I__5393 (
            .O(N__26219),
            .I(N__26205));
    LocalMux I__5392 (
            .O(N__26216),
            .I(N__26205));
    Span4Mux_s1_h I__5391 (
            .O(N__26213),
            .I(N__26200));
    Span4Mux_h I__5390 (
            .O(N__26210),
            .I(N__26200));
    Span4Mux_v I__5389 (
            .O(N__26205),
            .I(N__26197));
    Odrv4 I__5388 (
            .O(N__26200),
            .I(func_state_RNI_0_0));
    Odrv4 I__5387 (
            .O(N__26197),
            .I(func_state_RNI_0_0));
    InMux I__5386 (
            .O(N__26192),
            .I(N__26186));
    InMux I__5385 (
            .O(N__26191),
            .I(N__26186));
    LocalMux I__5384 (
            .O(N__26186),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_0 ));
    CascadeMux I__5383 (
            .O(N__26183),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_0_cascade_ ));
    CascadeMux I__5382 (
            .O(N__26180),
            .I(N__26176));
    InMux I__5381 (
            .O(N__26179),
            .I(N__26171));
    InMux I__5380 (
            .O(N__26176),
            .I(N__26164));
    InMux I__5379 (
            .O(N__26175),
            .I(N__26164));
    InMux I__5378 (
            .O(N__26174),
            .I(N__26164));
    LocalMux I__5377 (
            .O(N__26171),
            .I(N__26161));
    LocalMux I__5376 (
            .O(N__26164),
            .I(N__26158));
    Span4Mux_v I__5375 (
            .O(N__26161),
            .I(N__26155));
    Span4Mux_s3_h I__5374 (
            .O(N__26158),
            .I(N__26152));
    Odrv4 I__5373 (
            .O(N__26155),
            .I(\POWERLED.dutycycle_N_3_mux_0 ));
    Odrv4 I__5372 (
            .O(N__26152),
            .I(\POWERLED.dutycycle_N_3_mux_0 ));
    CascadeMux I__5371 (
            .O(N__26147),
            .I(\POWERLED.N_668_cascade_ ));
    InMux I__5370 (
            .O(N__26144),
            .I(N__26141));
    LocalMux I__5369 (
            .O(N__26141),
            .I(N__26138));
    Odrv4 I__5368 (
            .O(N__26138),
            .I(\POWERLED.N_490 ));
    CascadeMux I__5367 (
            .O(N__26135),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_1_cascade_ ));
    InMux I__5366 (
            .O(N__26132),
            .I(N__26114));
    InMux I__5365 (
            .O(N__26131),
            .I(N__26114));
    InMux I__5364 (
            .O(N__26130),
            .I(N__26107));
    InMux I__5363 (
            .O(N__26129),
            .I(N__26107));
    InMux I__5362 (
            .O(N__26128),
            .I(N__26107));
    InMux I__5361 (
            .O(N__26127),
            .I(N__26102));
    InMux I__5360 (
            .O(N__26126),
            .I(N__26102));
    InMux I__5359 (
            .O(N__26125),
            .I(N__26087));
    InMux I__5358 (
            .O(N__26124),
            .I(N__26087));
    InMux I__5357 (
            .O(N__26123),
            .I(N__26087));
    InMux I__5356 (
            .O(N__26122),
            .I(N__26087));
    InMux I__5355 (
            .O(N__26121),
            .I(N__26080));
    InMux I__5354 (
            .O(N__26120),
            .I(N__26080));
    InMux I__5353 (
            .O(N__26119),
            .I(N__26080));
    LocalMux I__5352 (
            .O(N__26114),
            .I(N__26077));
    LocalMux I__5351 (
            .O(N__26107),
            .I(N__26072));
    LocalMux I__5350 (
            .O(N__26102),
            .I(N__26072));
    InMux I__5349 (
            .O(N__26101),
            .I(N__26059));
    InMux I__5348 (
            .O(N__26100),
            .I(N__26059));
    InMux I__5347 (
            .O(N__26099),
            .I(N__26059));
    InMux I__5346 (
            .O(N__26098),
            .I(N__26059));
    InMux I__5345 (
            .O(N__26097),
            .I(N__26059));
    InMux I__5344 (
            .O(N__26096),
            .I(N__26059));
    LocalMux I__5343 (
            .O(N__26087),
            .I(N__26056));
    LocalMux I__5342 (
            .O(N__26080),
            .I(N__26053));
    Span4Mux_s2_v I__5341 (
            .O(N__26077),
            .I(N__26046));
    Span4Mux_h I__5340 (
            .O(N__26072),
            .I(N__26046));
    LocalMux I__5339 (
            .O(N__26059),
            .I(N__26046));
    Span4Mux_v I__5338 (
            .O(N__26056),
            .I(N__26041));
    Span4Mux_v I__5337 (
            .O(N__26053),
            .I(N__26041));
    Span4Mux_v I__5336 (
            .O(N__26046),
            .I(N__26038));
    Odrv4 I__5335 (
            .O(N__26041),
            .I(\POWERLED.N_123 ));
    Odrv4 I__5334 (
            .O(N__26038),
            .I(\POWERLED.N_123 ));
    InMux I__5333 (
            .O(N__26033),
            .I(N__26030));
    LocalMux I__5332 (
            .O(N__26030),
            .I(N__26026));
    InMux I__5331 (
            .O(N__26029),
            .I(N__26023));
    Span4Mux_h I__5330 (
            .O(N__26026),
            .I(N__26020));
    LocalMux I__5329 (
            .O(N__26023),
            .I(\POWERLED.N_443 ));
    Odrv4 I__5328 (
            .O(N__26020),
            .I(\POWERLED.N_443 ));
    CascadeMux I__5327 (
            .O(N__26015),
            .I(N__26011));
    CascadeMux I__5326 (
            .O(N__26014),
            .I(N__26007));
    InMux I__5325 (
            .O(N__26011),
            .I(N__26004));
    InMux I__5324 (
            .O(N__26010),
            .I(N__25999));
    InMux I__5323 (
            .O(N__26007),
            .I(N__25999));
    LocalMux I__5322 (
            .O(N__26004),
            .I(N__25996));
    LocalMux I__5321 (
            .O(N__25999),
            .I(N__25991));
    Span4Mux_h I__5320 (
            .O(N__25996),
            .I(N__25991));
    Odrv4 I__5319 (
            .O(N__25991),
            .I(\POWERLED.count_off_RNIH9TEZ0Z_10 ));
    InMux I__5318 (
            .O(N__25988),
            .I(N__25985));
    LocalMux I__5317 (
            .O(N__25985),
            .I(N__25982));
    Odrv12 I__5316 (
            .O(N__25982),
            .I(\POWERLED.un1_func_state25_6_0_0_0_2_1 ));
    InMux I__5315 (
            .O(N__25979),
            .I(N__25973));
    InMux I__5314 (
            .O(N__25978),
            .I(N__25973));
    LocalMux I__5313 (
            .O(N__25973),
            .I(\POWERLED.N_668 ));
    InMux I__5312 (
            .O(N__25970),
            .I(N__25966));
    CascadeMux I__5311 (
            .O(N__25969),
            .I(N__25963));
    LocalMux I__5310 (
            .O(N__25966),
            .I(N__25960));
    InMux I__5309 (
            .O(N__25963),
            .I(N__25957));
    Span12Mux_s3_h I__5308 (
            .O(N__25960),
            .I(N__25954));
    LocalMux I__5307 (
            .O(N__25957),
            .I(N__25951));
    Odrv12 I__5306 (
            .O(N__25954),
            .I(\POWERLED.count_off_1_sqmuxa ));
    Odrv12 I__5305 (
            .O(N__25951),
            .I(\POWERLED.count_off_1_sqmuxa ));
    InMux I__5304 (
            .O(N__25946),
            .I(N__25943));
    LocalMux I__5303 (
            .O(N__25943),
            .I(N__25940));
    Odrv4 I__5302 (
            .O(N__25940),
            .I(\POWERLED.un1_dutycycle_172_m0 ));
    CascadeMux I__5301 (
            .O(N__25937),
            .I(\POWERLED.un1_dutycycle_172_m1_ns_1_cascade_ ));
    InMux I__5300 (
            .O(N__25934),
            .I(N__25931));
    LocalMux I__5299 (
            .O(N__25931),
            .I(N__25928));
    Span4Mux_v I__5298 (
            .O(N__25928),
            .I(N__25925));
    Odrv4 I__5297 (
            .O(N__25925),
            .I(\POWERLED.un1_dutycycle_172_m1 ));
    CascadeMux I__5296 (
            .O(N__25922),
            .I(N__25918));
    CascadeMux I__5295 (
            .O(N__25921),
            .I(N__25915));
    InMux I__5294 (
            .O(N__25918),
            .I(N__25912));
    InMux I__5293 (
            .O(N__25915),
            .I(N__25909));
    LocalMux I__5292 (
            .O(N__25912),
            .I(N__25904));
    LocalMux I__5291 (
            .O(N__25909),
            .I(N__25904));
    Span4Mux_v I__5290 (
            .O(N__25904),
            .I(N__25901));
    Odrv4 I__5289 (
            .O(N__25901),
            .I(\POWERLED.func_state_RNI_3Z0Z_1 ));
    CascadeMux I__5288 (
            .O(N__25898),
            .I(\POWERLED.count_clk_RNIZ0Z_0_cascade_ ));
    CascadeMux I__5287 (
            .O(N__25895),
            .I(\POWERLED.count_clkZ0Z_1_cascade_ ));
    InMux I__5286 (
            .O(N__25892),
            .I(N__25889));
    LocalMux I__5285 (
            .O(N__25889),
            .I(\POWERLED.count_clk_0_1 ));
    CascadeMux I__5284 (
            .O(N__25886),
            .I(N__25883));
    InMux I__5283 (
            .O(N__25883),
            .I(N__25880));
    LocalMux I__5282 (
            .O(N__25880),
            .I(N__25877));
    Odrv4 I__5281 (
            .O(N__25877),
            .I(\POWERLED.count_clk_0_11 ));
    InMux I__5280 (
            .O(N__25874),
            .I(N__25868));
    CascadeMux I__5279 (
            .O(N__25873),
            .I(N__25861));
    InMux I__5278 (
            .O(N__25872),
            .I(N__25858));
    InMux I__5277 (
            .O(N__25871),
            .I(N__25855));
    LocalMux I__5276 (
            .O(N__25868),
            .I(N__25852));
    InMux I__5275 (
            .O(N__25867),
            .I(N__25847));
    InMux I__5274 (
            .O(N__25866),
            .I(N__25847));
    InMux I__5273 (
            .O(N__25865),
            .I(N__25844));
    InMux I__5272 (
            .O(N__25864),
            .I(N__25839));
    InMux I__5271 (
            .O(N__25861),
            .I(N__25839));
    LocalMux I__5270 (
            .O(N__25858),
            .I(N__25836));
    LocalMux I__5269 (
            .O(N__25855),
            .I(N__25833));
    Span4Mux_v I__5268 (
            .O(N__25852),
            .I(N__25830));
    LocalMux I__5267 (
            .O(N__25847),
            .I(N__25823));
    LocalMux I__5266 (
            .O(N__25844),
            .I(N__25823));
    LocalMux I__5265 (
            .O(N__25839),
            .I(N__25823));
    Span4Mux_s2_h I__5264 (
            .O(N__25836),
            .I(N__25820));
    Span4Mux_s2_h I__5263 (
            .O(N__25833),
            .I(N__25817));
    Odrv4 I__5262 (
            .O(N__25830),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv4 I__5261 (
            .O(N__25823),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv4 I__5260 (
            .O(N__25820),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv4 I__5259 (
            .O(N__25817),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    CascadeMux I__5258 (
            .O(N__25808),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_8_3_cascade_ ));
    SRMux I__5257 (
            .O(N__25805),
            .I(N__25802));
    LocalMux I__5256 (
            .O(N__25802),
            .I(N__25797));
    SRMux I__5255 (
            .O(N__25801),
            .I(N__25794));
    SRMux I__5254 (
            .O(N__25800),
            .I(N__25791));
    Span4Mux_v I__5253 (
            .O(N__25797),
            .I(N__25786));
    LocalMux I__5252 (
            .O(N__25794),
            .I(N__25786));
    LocalMux I__5251 (
            .O(N__25791),
            .I(N__25783));
    Span4Mux_s2_v I__5250 (
            .O(N__25786),
            .I(N__25778));
    Span4Mux_s1_h I__5249 (
            .O(N__25783),
            .I(N__25778));
    Odrv4 I__5248 (
            .O(N__25778),
            .I(G_30));
    InMux I__5247 (
            .O(N__25775),
            .I(N__25772));
    LocalMux I__5246 (
            .O(N__25772),
            .I(\POWERLED.count_clk_0_4 ));
    InMux I__5245 (
            .O(N__25769),
            .I(N__25766));
    LocalMux I__5244 (
            .O(N__25766),
            .I(\POWERLED.count_clk_0_5 ));
    InMux I__5243 (
            .O(N__25763),
            .I(N__25760));
    LocalMux I__5242 (
            .O(N__25760),
            .I(\POWERLED.count_clk_0_6 ));
    InMux I__5241 (
            .O(N__25757),
            .I(N__25727));
    InMux I__5240 (
            .O(N__25756),
            .I(N__25727));
    InMux I__5239 (
            .O(N__25755),
            .I(N__25718));
    InMux I__5238 (
            .O(N__25754),
            .I(N__25718));
    InMux I__5237 (
            .O(N__25753),
            .I(N__25718));
    InMux I__5236 (
            .O(N__25752),
            .I(N__25718));
    InMux I__5235 (
            .O(N__25751),
            .I(N__25709));
    InMux I__5234 (
            .O(N__25750),
            .I(N__25709));
    InMux I__5233 (
            .O(N__25749),
            .I(N__25709));
    InMux I__5232 (
            .O(N__25748),
            .I(N__25709));
    InMux I__5231 (
            .O(N__25747),
            .I(N__25702));
    InMux I__5230 (
            .O(N__25746),
            .I(N__25702));
    InMux I__5229 (
            .O(N__25745),
            .I(N__25702));
    CascadeMux I__5228 (
            .O(N__25744),
            .I(N__25699));
    InMux I__5227 (
            .O(N__25743),
            .I(N__25694));
    InMux I__5226 (
            .O(N__25742),
            .I(N__25687));
    InMux I__5225 (
            .O(N__25741),
            .I(N__25687));
    InMux I__5224 (
            .O(N__25740),
            .I(N__25687));
    InMux I__5223 (
            .O(N__25739),
            .I(N__25684));
    InMux I__5222 (
            .O(N__25738),
            .I(N__25673));
    InMux I__5221 (
            .O(N__25737),
            .I(N__25673));
    InMux I__5220 (
            .O(N__25736),
            .I(N__25673));
    InMux I__5219 (
            .O(N__25735),
            .I(N__25673));
    InMux I__5218 (
            .O(N__25734),
            .I(N__25673));
    InMux I__5217 (
            .O(N__25733),
            .I(N__25668));
    InMux I__5216 (
            .O(N__25732),
            .I(N__25668));
    LocalMux I__5215 (
            .O(N__25727),
            .I(N__25659));
    LocalMux I__5214 (
            .O(N__25718),
            .I(N__25659));
    LocalMux I__5213 (
            .O(N__25709),
            .I(N__25659));
    LocalMux I__5212 (
            .O(N__25702),
            .I(N__25659));
    InMux I__5211 (
            .O(N__25699),
            .I(N__25648));
    InMux I__5210 (
            .O(N__25698),
            .I(N__25648));
    InMux I__5209 (
            .O(N__25697),
            .I(N__25648));
    LocalMux I__5208 (
            .O(N__25694),
            .I(N__25635));
    LocalMux I__5207 (
            .O(N__25687),
            .I(N__25635));
    LocalMux I__5206 (
            .O(N__25684),
            .I(N__25635));
    LocalMux I__5205 (
            .O(N__25673),
            .I(N__25635));
    LocalMux I__5204 (
            .O(N__25668),
            .I(N__25635));
    Span4Mux_v I__5203 (
            .O(N__25659),
            .I(N__25635));
    InMux I__5202 (
            .O(N__25658),
            .I(N__25631));
    InMux I__5201 (
            .O(N__25657),
            .I(N__25624));
    InMux I__5200 (
            .O(N__25656),
            .I(N__25624));
    InMux I__5199 (
            .O(N__25655),
            .I(N__25624));
    LocalMux I__5198 (
            .O(N__25648),
            .I(N__25621));
    Span4Mux_v I__5197 (
            .O(N__25635),
            .I(N__25616));
    InMux I__5196 (
            .O(N__25634),
            .I(N__25613));
    LocalMux I__5195 (
            .O(N__25631),
            .I(N__25610));
    LocalMux I__5194 (
            .O(N__25624),
            .I(N__25605));
    Span12Mux_s6_h I__5193 (
            .O(N__25621),
            .I(N__25605));
    InMux I__5192 (
            .O(N__25620),
            .I(N__25600));
    InMux I__5191 (
            .O(N__25619),
            .I(N__25600));
    Sp12to4 I__5190 (
            .O(N__25616),
            .I(N__25595));
    LocalMux I__5189 (
            .O(N__25613),
            .I(N__25595));
    Odrv4 I__5188 (
            .O(N__25610),
            .I(clk_100Khz_signalkeep_3));
    Odrv12 I__5187 (
            .O(N__25605),
            .I(clk_100Khz_signalkeep_3));
    LocalMux I__5186 (
            .O(N__25600),
            .I(clk_100Khz_signalkeep_3));
    Odrv12 I__5185 (
            .O(N__25595),
            .I(clk_100Khz_signalkeep_3));
    InMux I__5184 (
            .O(N__25586),
            .I(N__25583));
    LocalMux I__5183 (
            .O(N__25583),
            .I(N__25574));
    InMux I__5182 (
            .O(N__25582),
            .I(N__25569));
    InMux I__5181 (
            .O(N__25581),
            .I(N__25569));
    InMux I__5180 (
            .O(N__25580),
            .I(N__25566));
    InMux I__5179 (
            .O(N__25579),
            .I(N__25561));
    InMux I__5178 (
            .O(N__25578),
            .I(N__25561));
    InMux I__5177 (
            .O(N__25577),
            .I(N__25558));
    Span4Mux_h I__5176 (
            .O(N__25574),
            .I(N__25553));
    LocalMux I__5175 (
            .O(N__25569),
            .I(N__25553));
    LocalMux I__5174 (
            .O(N__25566),
            .I(clk_100Khz_signalkeep_3_rep1));
    LocalMux I__5173 (
            .O(N__25561),
            .I(clk_100Khz_signalkeep_3_rep1));
    LocalMux I__5172 (
            .O(N__25558),
            .I(clk_100Khz_signalkeep_3_rep1));
    Odrv4 I__5171 (
            .O(N__25553),
            .I(clk_100Khz_signalkeep_3_rep1));
    InMux I__5170 (
            .O(N__25544),
            .I(N__25540));
    InMux I__5169 (
            .O(N__25543),
            .I(N__25537));
    LocalMux I__5168 (
            .O(N__25540),
            .I(N__25534));
    LocalMux I__5167 (
            .O(N__25537),
            .I(N__25529));
    Span4Mux_s2_v I__5166 (
            .O(N__25534),
            .I(N__25529));
    Odrv4 I__5165 (
            .O(N__25529),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    InMux I__5164 (
            .O(N__25526),
            .I(\VPP_VDDQ.un1_count_1_cry_8 ));
    CascadeMux I__5163 (
            .O(N__25523),
            .I(N__25520));
    InMux I__5162 (
            .O(N__25520),
            .I(N__25517));
    LocalMux I__5161 (
            .O(N__25517),
            .I(N__25513));
    InMux I__5160 (
            .O(N__25516),
            .I(N__25510));
    Span4Mux_h I__5159 (
            .O(N__25513),
            .I(N__25507));
    LocalMux I__5158 (
            .O(N__25510),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    Odrv4 I__5157 (
            .O(N__25507),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    InMux I__5156 (
            .O(N__25502),
            .I(\VPP_VDDQ.un1_count_1_cry_9 ));
    CascadeMux I__5155 (
            .O(N__25499),
            .I(N__25496));
    InMux I__5154 (
            .O(N__25496),
            .I(N__25493));
    LocalMux I__5153 (
            .O(N__25493),
            .I(N__25489));
    InMux I__5152 (
            .O(N__25492),
            .I(N__25486));
    Span4Mux_s2_v I__5151 (
            .O(N__25489),
            .I(N__25483));
    LocalMux I__5150 (
            .O(N__25486),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    Odrv4 I__5149 (
            .O(N__25483),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    InMux I__5148 (
            .O(N__25478),
            .I(\VPP_VDDQ.un1_count_1_cry_10 ));
    InMux I__5147 (
            .O(N__25475),
            .I(N__25472));
    LocalMux I__5146 (
            .O(N__25472),
            .I(N__25468));
    InMux I__5145 (
            .O(N__25471),
            .I(N__25465));
    Span4Mux_s2_v I__5144 (
            .O(N__25468),
            .I(N__25462));
    LocalMux I__5143 (
            .O(N__25465),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    Odrv4 I__5142 (
            .O(N__25462),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    InMux I__5141 (
            .O(N__25457),
            .I(\VPP_VDDQ.un1_count_1_cry_11 ));
    InMux I__5140 (
            .O(N__25454),
            .I(N__25451));
    LocalMux I__5139 (
            .O(N__25451),
            .I(N__25447));
    InMux I__5138 (
            .O(N__25450),
            .I(N__25444));
    Span4Mux_h I__5137 (
            .O(N__25447),
            .I(N__25441));
    LocalMux I__5136 (
            .O(N__25444),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    Odrv4 I__5135 (
            .O(N__25441),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    InMux I__5134 (
            .O(N__25436),
            .I(\VPP_VDDQ.un1_count_1_cry_12 ));
    InMux I__5133 (
            .O(N__25433),
            .I(N__25390));
    InMux I__5132 (
            .O(N__25432),
            .I(N__25390));
    InMux I__5131 (
            .O(N__25431),
            .I(N__25390));
    InMux I__5130 (
            .O(N__25430),
            .I(N__25390));
    InMux I__5129 (
            .O(N__25429),
            .I(N__25381));
    InMux I__5128 (
            .O(N__25428),
            .I(N__25381));
    InMux I__5127 (
            .O(N__25427),
            .I(N__25381));
    InMux I__5126 (
            .O(N__25426),
            .I(N__25381));
    InMux I__5125 (
            .O(N__25425),
            .I(N__25372));
    InMux I__5124 (
            .O(N__25424),
            .I(N__25372));
    InMux I__5123 (
            .O(N__25423),
            .I(N__25372));
    InMux I__5122 (
            .O(N__25422),
            .I(N__25372));
    InMux I__5121 (
            .O(N__25421),
            .I(N__25363));
    InMux I__5120 (
            .O(N__25420),
            .I(N__25363));
    InMux I__5119 (
            .O(N__25419),
            .I(N__25363));
    InMux I__5118 (
            .O(N__25418),
            .I(N__25363));
    InMux I__5117 (
            .O(N__25417),
            .I(N__25356));
    InMux I__5116 (
            .O(N__25416),
            .I(N__25356));
    InMux I__5115 (
            .O(N__25415),
            .I(N__25356));
    InMux I__5114 (
            .O(N__25414),
            .I(N__25347));
    InMux I__5113 (
            .O(N__25413),
            .I(N__25347));
    InMux I__5112 (
            .O(N__25412),
            .I(N__25347));
    InMux I__5111 (
            .O(N__25411),
            .I(N__25347));
    InMux I__5110 (
            .O(N__25410),
            .I(N__25340));
    InMux I__5109 (
            .O(N__25409),
            .I(N__25340));
    InMux I__5108 (
            .O(N__25408),
            .I(N__25340));
    InMux I__5107 (
            .O(N__25407),
            .I(N__25331));
    InMux I__5106 (
            .O(N__25406),
            .I(N__25331));
    InMux I__5105 (
            .O(N__25405),
            .I(N__25331));
    InMux I__5104 (
            .O(N__25404),
            .I(N__25331));
    InMux I__5103 (
            .O(N__25403),
            .I(N__25328));
    InMux I__5102 (
            .O(N__25402),
            .I(N__25325));
    InMux I__5101 (
            .O(N__25401),
            .I(N__25320));
    InMux I__5100 (
            .O(N__25400),
            .I(N__25320));
    InMux I__5099 (
            .O(N__25399),
            .I(N__25317));
    LocalMux I__5098 (
            .O(N__25390),
            .I(N__25305));
    LocalMux I__5097 (
            .O(N__25381),
            .I(N__25302));
    LocalMux I__5096 (
            .O(N__25372),
            .I(N__25299));
    LocalMux I__5095 (
            .O(N__25363),
            .I(N__25296));
    LocalMux I__5094 (
            .O(N__25356),
            .I(N__25293));
    LocalMux I__5093 (
            .O(N__25347),
            .I(N__25290));
    LocalMux I__5092 (
            .O(N__25340),
            .I(N__25287));
    LocalMux I__5091 (
            .O(N__25331),
            .I(N__25284));
    LocalMux I__5090 (
            .O(N__25328),
            .I(N__25281));
    LocalMux I__5089 (
            .O(N__25325),
            .I(N__25278));
    LocalMux I__5088 (
            .O(N__25320),
            .I(N__25275));
    LocalMux I__5087 (
            .O(N__25317),
            .I(N__25272));
    CEMux I__5086 (
            .O(N__25316),
            .I(N__25229));
    CEMux I__5085 (
            .O(N__25315),
            .I(N__25229));
    CEMux I__5084 (
            .O(N__25314),
            .I(N__25229));
    CEMux I__5083 (
            .O(N__25313),
            .I(N__25229));
    CEMux I__5082 (
            .O(N__25312),
            .I(N__25229));
    CEMux I__5081 (
            .O(N__25311),
            .I(N__25229));
    CEMux I__5080 (
            .O(N__25310),
            .I(N__25229));
    CEMux I__5079 (
            .O(N__25309),
            .I(N__25229));
    CEMux I__5078 (
            .O(N__25308),
            .I(N__25229));
    Glb2LocalMux I__5077 (
            .O(N__25305),
            .I(N__25229));
    Glb2LocalMux I__5076 (
            .O(N__25302),
            .I(N__25229));
    Glb2LocalMux I__5075 (
            .O(N__25299),
            .I(N__25229));
    Glb2LocalMux I__5074 (
            .O(N__25296),
            .I(N__25229));
    Glb2LocalMux I__5073 (
            .O(N__25293),
            .I(N__25229));
    Glb2LocalMux I__5072 (
            .O(N__25290),
            .I(N__25229));
    Glb2LocalMux I__5071 (
            .O(N__25287),
            .I(N__25229));
    Glb2LocalMux I__5070 (
            .O(N__25284),
            .I(N__25229));
    Glb2LocalMux I__5069 (
            .O(N__25281),
            .I(N__25229));
    Glb2LocalMux I__5068 (
            .O(N__25278),
            .I(N__25229));
    Glb2LocalMux I__5067 (
            .O(N__25275),
            .I(N__25229));
    Glb2LocalMux I__5066 (
            .O(N__25272),
            .I(N__25229));
    GlobalMux I__5065 (
            .O(N__25229),
            .I(N__25226));
    gio2CtrlBuf I__5064 (
            .O(N__25226),
            .I(N_92_g));
    InMux I__5063 (
            .O(N__25223),
            .I(N__25219));
    InMux I__5062 (
            .O(N__25222),
            .I(N__25216));
    LocalMux I__5061 (
            .O(N__25219),
            .I(N__25213));
    LocalMux I__5060 (
            .O(N__25216),
            .I(N__25208));
    Span4Mux_s2_v I__5059 (
            .O(N__25213),
            .I(N__25208));
    Odrv4 I__5058 (
            .O(N__25208),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    InMux I__5057 (
            .O(N__25205),
            .I(\VPP_VDDQ.un1_count_1_cry_13 ));
    IoInMux I__5056 (
            .O(N__25202),
            .I(N__25199));
    LocalMux I__5055 (
            .O(N__25199),
            .I(N__25196));
    IoSpan4Mux I__5054 (
            .O(N__25196),
            .I(N__25190));
    InMux I__5053 (
            .O(N__25195),
            .I(N__25187));
    InMux I__5052 (
            .O(N__25194),
            .I(N__25184));
    InMux I__5051 (
            .O(N__25193),
            .I(N__25177));
    IoSpan4Mux I__5050 (
            .O(N__25190),
            .I(N__25174));
    LocalMux I__5049 (
            .O(N__25187),
            .I(N__25169));
    LocalMux I__5048 (
            .O(N__25184),
            .I(N__25169));
    InMux I__5047 (
            .O(N__25183),
            .I(N__25166));
    InMux I__5046 (
            .O(N__25182),
            .I(N__25163));
    IoInMux I__5045 (
            .O(N__25181),
            .I(N__25160));
    InMux I__5044 (
            .O(N__25180),
            .I(N__25157));
    LocalMux I__5043 (
            .O(N__25177),
            .I(N__25154));
    Span4Mux_s0_h I__5042 (
            .O(N__25174),
            .I(N__25151));
    Span4Mux_v I__5041 (
            .O(N__25169),
            .I(N__25148));
    LocalMux I__5040 (
            .O(N__25166),
            .I(N__25143));
    LocalMux I__5039 (
            .O(N__25163),
            .I(N__25143));
    LocalMux I__5038 (
            .O(N__25160),
            .I(N__25140));
    LocalMux I__5037 (
            .O(N__25157),
            .I(N__25137));
    Span12Mux_s2_h I__5036 (
            .O(N__25154),
            .I(N__25134));
    Span4Mux_h I__5035 (
            .O(N__25151),
            .I(N__25127));
    Span4Mux_s2_v I__5034 (
            .O(N__25148),
            .I(N__25127));
    Span4Mux_v I__5033 (
            .O(N__25143),
            .I(N__25127));
    IoSpan4Mux I__5032 (
            .O(N__25140),
            .I(N__25124));
    Span12Mux_v I__5031 (
            .O(N__25137),
            .I(N__25121));
    Span12Mux_v I__5030 (
            .O(N__25134),
            .I(N__25118));
    Span4Mux_h I__5029 (
            .O(N__25127),
            .I(N__25113));
    IoSpan4Mux I__5028 (
            .O(N__25124),
            .I(N__25113));
    Odrv12 I__5027 (
            .O(N__25121),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__5026 (
            .O(N__25118),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5025 (
            .O(N__25113),
            .I(CONSTANT_ONE_NET));
    InMux I__5024 (
            .O(N__25106),
            .I(bfn_11_4_0_));
    CascadeMux I__5023 (
            .O(N__25103),
            .I(N__25100));
    InMux I__5022 (
            .O(N__25100),
            .I(N__25097));
    LocalMux I__5021 (
            .O(N__25097),
            .I(N__25093));
    InMux I__5020 (
            .O(N__25096),
            .I(N__25090));
    Span4Mux_h I__5019 (
            .O(N__25093),
            .I(N__25087));
    LocalMux I__5018 (
            .O(N__25090),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    Odrv4 I__5017 (
            .O(N__25087),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    CEMux I__5016 (
            .O(N__25082),
            .I(N__25079));
    LocalMux I__5015 (
            .O(N__25079),
            .I(N__25076));
    Span4Mux_s2_h I__5014 (
            .O(N__25076),
            .I(N__25073));
    Odrv4 I__5013 (
            .O(N__25073),
            .I(\VPP_VDDQ.N_92_0 ));
    InMux I__5012 (
            .O(N__25070),
            .I(N__25066));
    InMux I__5011 (
            .O(N__25069),
            .I(N__25063));
    LocalMux I__5010 (
            .O(N__25066),
            .I(N__25060));
    LocalMux I__5009 (
            .O(N__25063),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    Odrv4 I__5008 (
            .O(N__25060),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    InMux I__5007 (
            .O(N__25055),
            .I(\VPP_VDDQ.un1_count_1_cry_0 ));
    InMux I__5006 (
            .O(N__25052),
            .I(N__25048));
    InMux I__5005 (
            .O(N__25051),
            .I(N__25045));
    LocalMux I__5004 (
            .O(N__25048),
            .I(N__25042));
    LocalMux I__5003 (
            .O(N__25045),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    Odrv4 I__5002 (
            .O(N__25042),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    InMux I__5001 (
            .O(N__25037),
            .I(\VPP_VDDQ.un1_count_1_cry_1 ));
    InMux I__5000 (
            .O(N__25034),
            .I(N__25030));
    InMux I__4999 (
            .O(N__25033),
            .I(N__25027));
    LocalMux I__4998 (
            .O(N__25030),
            .I(N__25024));
    LocalMux I__4997 (
            .O(N__25027),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    Odrv4 I__4996 (
            .O(N__25024),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    InMux I__4995 (
            .O(N__25019),
            .I(\VPP_VDDQ.un1_count_1_cry_2 ));
    InMux I__4994 (
            .O(N__25016),
            .I(N__25012));
    InMux I__4993 (
            .O(N__25015),
            .I(N__25009));
    LocalMux I__4992 (
            .O(N__25012),
            .I(N__25006));
    LocalMux I__4991 (
            .O(N__25009),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    Odrv4 I__4990 (
            .O(N__25006),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    InMux I__4989 (
            .O(N__25001),
            .I(\VPP_VDDQ.un1_count_1_cry_3 ));
    InMux I__4988 (
            .O(N__24998),
            .I(N__24994));
    InMux I__4987 (
            .O(N__24997),
            .I(N__24991));
    LocalMux I__4986 (
            .O(N__24994),
            .I(N__24988));
    LocalMux I__4985 (
            .O(N__24991),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    Odrv4 I__4984 (
            .O(N__24988),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    InMux I__4983 (
            .O(N__24983),
            .I(\VPP_VDDQ.un1_count_1_cry_4 ));
    InMux I__4982 (
            .O(N__24980),
            .I(N__24976));
    InMux I__4981 (
            .O(N__24979),
            .I(N__24973));
    LocalMux I__4980 (
            .O(N__24976),
            .I(N__24970));
    LocalMux I__4979 (
            .O(N__24973),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    Odrv12 I__4978 (
            .O(N__24970),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    InMux I__4977 (
            .O(N__24965),
            .I(\VPP_VDDQ.un1_count_1_cry_5 ));
    CascadeMux I__4976 (
            .O(N__24962),
            .I(N__24959));
    InMux I__4975 (
            .O(N__24959),
            .I(N__24955));
    InMux I__4974 (
            .O(N__24958),
            .I(N__24952));
    LocalMux I__4973 (
            .O(N__24955),
            .I(N__24949));
    LocalMux I__4972 (
            .O(N__24952),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    Odrv4 I__4971 (
            .O(N__24949),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    InMux I__4970 (
            .O(N__24944),
            .I(\VPP_VDDQ.un1_count_1_cry_6 ));
    InMux I__4969 (
            .O(N__24941),
            .I(N__24937));
    InMux I__4968 (
            .O(N__24940),
            .I(N__24934));
    LocalMux I__4967 (
            .O(N__24937),
            .I(N__24931));
    LocalMux I__4966 (
            .O(N__24934),
            .I(N__24926));
    Span4Mux_s2_v I__4965 (
            .O(N__24931),
            .I(N__24926));
    Odrv4 I__4964 (
            .O(N__24926),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    InMux I__4963 (
            .O(N__24923),
            .I(bfn_11_3_0_));
    InMux I__4962 (
            .O(N__24920),
            .I(N__24914));
    InMux I__4961 (
            .O(N__24919),
            .I(N__24914));
    LocalMux I__4960 (
            .O(N__24914),
            .I(N__24911));
    Odrv12 I__4959 (
            .O(N__24911),
            .I(\POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ));
    CascadeMux I__4958 (
            .O(N__24908),
            .I(N__24905));
    InMux I__4957 (
            .O(N__24905),
            .I(N__24899));
    InMux I__4956 (
            .O(N__24904),
            .I(N__24899));
    LocalMux I__4955 (
            .O(N__24899),
            .I(N__24896));
    Span12Mux_s5_h I__4954 (
            .O(N__24896),
            .I(N__24893));
    Odrv12 I__4953 (
            .O(N__24893),
            .I(\POWERLED.dutycycle_en_4 ));
    CascadeMux I__4952 (
            .O(N__24890),
            .I(N__24887));
    InMux I__4951 (
            .O(N__24887),
            .I(N__24881));
    InMux I__4950 (
            .O(N__24886),
            .I(N__24881));
    LocalMux I__4949 (
            .O(N__24881),
            .I(\POWERLED.dutycycleZ1Z_10 ));
    CascadeMux I__4948 (
            .O(N__24878),
            .I(\POWERLED.dutycycleZ0Z_2_cascade_ ));
    InMux I__4947 (
            .O(N__24875),
            .I(N__24872));
    LocalMux I__4946 (
            .O(N__24872),
            .I(N__24869));
    Odrv4 I__4945 (
            .O(N__24869),
            .I(\POWERLED.un2_count_clk_17_0_0_a2_0_0 ));
    InMux I__4944 (
            .O(N__24866),
            .I(N__24863));
    LocalMux I__4943 (
            .O(N__24863),
            .I(\POWERLED.un1_dutycycle_53_50_0_0 ));
    InMux I__4942 (
            .O(N__24860),
            .I(N__24853));
    InMux I__4941 (
            .O(N__24859),
            .I(N__24850));
    InMux I__4940 (
            .O(N__24858),
            .I(N__24843));
    InMux I__4939 (
            .O(N__24857),
            .I(N__24843));
    InMux I__4938 (
            .O(N__24856),
            .I(N__24843));
    LocalMux I__4937 (
            .O(N__24853),
            .I(N__24840));
    LocalMux I__4936 (
            .O(N__24850),
            .I(\POWERLED.un1_dutycycle_53_4_0 ));
    LocalMux I__4935 (
            .O(N__24843),
            .I(\POWERLED.un1_dutycycle_53_4_0 ));
    Odrv4 I__4934 (
            .O(N__24840),
            .I(\POWERLED.un1_dutycycle_53_4_0 ));
    CascadeMux I__4933 (
            .O(N__24833),
            .I(\POWERLED.un1_dutycycle_53_10_2_cascade_ ));
    InMux I__4932 (
            .O(N__24830),
            .I(N__24827));
    LocalMux I__4931 (
            .O(N__24827),
            .I(N__24824));
    Odrv4 I__4930 (
            .O(N__24824),
            .I(\POWERLED.un1_dutycycle_53_10_3 ));
    InMux I__4929 (
            .O(N__24821),
            .I(N__24818));
    LocalMux I__4928 (
            .O(N__24818),
            .I(\POWERLED.un1_dutycycle_53_9_a1_0 ));
    CascadeMux I__4927 (
            .O(N__24815),
            .I(N__24810));
    CascadeMux I__4926 (
            .O(N__24814),
            .I(N__24806));
    InMux I__4925 (
            .O(N__24813),
            .I(N__24803));
    InMux I__4924 (
            .O(N__24810),
            .I(N__24800));
    CascadeMux I__4923 (
            .O(N__24809),
            .I(N__24797));
    InMux I__4922 (
            .O(N__24806),
            .I(N__24790));
    LocalMux I__4921 (
            .O(N__24803),
            .I(N__24785));
    LocalMux I__4920 (
            .O(N__24800),
            .I(N__24785));
    InMux I__4919 (
            .O(N__24797),
            .I(N__24782));
    InMux I__4918 (
            .O(N__24796),
            .I(N__24779));
    CascadeMux I__4917 (
            .O(N__24795),
            .I(N__24774));
    InMux I__4916 (
            .O(N__24794),
            .I(N__24771));
    InMux I__4915 (
            .O(N__24793),
            .I(N__24768));
    LocalMux I__4914 (
            .O(N__24790),
            .I(N__24762));
    Span4Mux_h I__4913 (
            .O(N__24785),
            .I(N__24762));
    LocalMux I__4912 (
            .O(N__24782),
            .I(N__24757));
    LocalMux I__4911 (
            .O(N__24779),
            .I(N__24757));
    InMux I__4910 (
            .O(N__24778),
            .I(N__24750));
    InMux I__4909 (
            .O(N__24777),
            .I(N__24750));
    InMux I__4908 (
            .O(N__24774),
            .I(N__24750));
    LocalMux I__4907 (
            .O(N__24771),
            .I(N__24743));
    LocalMux I__4906 (
            .O(N__24768),
            .I(N__24740));
    InMux I__4905 (
            .O(N__24767),
            .I(N__24737));
    Span4Mux_v I__4904 (
            .O(N__24762),
            .I(N__24732));
    Span4Mux_h I__4903 (
            .O(N__24757),
            .I(N__24732));
    LocalMux I__4902 (
            .O(N__24750),
            .I(N__24729));
    InMux I__4901 (
            .O(N__24749),
            .I(N__24720));
    InMux I__4900 (
            .O(N__24748),
            .I(N__24720));
    InMux I__4899 (
            .O(N__24747),
            .I(N__24720));
    InMux I__4898 (
            .O(N__24746),
            .I(N__24720));
    Odrv4 I__4897 (
            .O(N__24743),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv12 I__4896 (
            .O(N__24740),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__4895 (
            .O(N__24737),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__4894 (
            .O(N__24732),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__4893 (
            .O(N__24729),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__4892 (
            .O(N__24720),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    CascadeMux I__4891 (
            .O(N__24707),
            .I(N__24697));
    InMux I__4890 (
            .O(N__24706),
            .I(N__24692));
    InMux I__4889 (
            .O(N__24705),
            .I(N__24689));
    InMux I__4888 (
            .O(N__24704),
            .I(N__24682));
    InMux I__4887 (
            .O(N__24703),
            .I(N__24682));
    InMux I__4886 (
            .O(N__24702),
            .I(N__24682));
    InMux I__4885 (
            .O(N__24701),
            .I(N__24679));
    InMux I__4884 (
            .O(N__24700),
            .I(N__24673));
    InMux I__4883 (
            .O(N__24697),
            .I(N__24670));
    InMux I__4882 (
            .O(N__24696),
            .I(N__24665));
    InMux I__4881 (
            .O(N__24695),
            .I(N__24665));
    LocalMux I__4880 (
            .O(N__24692),
            .I(N__24660));
    LocalMux I__4879 (
            .O(N__24689),
            .I(N__24660));
    LocalMux I__4878 (
            .O(N__24682),
            .I(N__24657));
    LocalMux I__4877 (
            .O(N__24679),
            .I(N__24654));
    InMux I__4876 (
            .O(N__24678),
            .I(N__24649));
    InMux I__4875 (
            .O(N__24677),
            .I(N__24649));
    InMux I__4874 (
            .O(N__24676),
            .I(N__24646));
    LocalMux I__4873 (
            .O(N__24673),
            .I(N__24637));
    LocalMux I__4872 (
            .O(N__24670),
            .I(N__24637));
    LocalMux I__4871 (
            .O(N__24665),
            .I(N__24637));
    Span4Mux_v I__4870 (
            .O(N__24660),
            .I(N__24637));
    Span4Mux_v I__4869 (
            .O(N__24657),
            .I(N__24634));
    Odrv4 I__4868 (
            .O(N__24654),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__4867 (
            .O(N__24649),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__4866 (
            .O(N__24646),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__4865 (
            .O(N__24637),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__4864 (
            .O(N__24634),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    CascadeMux I__4863 (
            .O(N__24623),
            .I(N__24620));
    InMux I__4862 (
            .O(N__24620),
            .I(N__24615));
    InMux I__4861 (
            .O(N__24619),
            .I(N__24609));
    CascadeMux I__4860 (
            .O(N__24618),
            .I(N__24600));
    LocalMux I__4859 (
            .O(N__24615),
            .I(N__24596));
    InMux I__4858 (
            .O(N__24614),
            .I(N__24591));
    InMux I__4857 (
            .O(N__24613),
            .I(N__24591));
    InMux I__4856 (
            .O(N__24612),
            .I(N__24588));
    LocalMux I__4855 (
            .O(N__24609),
            .I(N__24585));
    InMux I__4854 (
            .O(N__24608),
            .I(N__24582));
    InMux I__4853 (
            .O(N__24607),
            .I(N__24579));
    InMux I__4852 (
            .O(N__24606),
            .I(N__24574));
    InMux I__4851 (
            .O(N__24605),
            .I(N__24574));
    InMux I__4850 (
            .O(N__24604),
            .I(N__24569));
    InMux I__4849 (
            .O(N__24603),
            .I(N__24569));
    InMux I__4848 (
            .O(N__24600),
            .I(N__24564));
    InMux I__4847 (
            .O(N__24599),
            .I(N__24564));
    Span4Mux_h I__4846 (
            .O(N__24596),
            .I(N__24557));
    LocalMux I__4845 (
            .O(N__24591),
            .I(N__24557));
    LocalMux I__4844 (
            .O(N__24588),
            .I(N__24557));
    Odrv4 I__4843 (
            .O(N__24585),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__4842 (
            .O(N__24582),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__4841 (
            .O(N__24579),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__4840 (
            .O(N__24574),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__4839 (
            .O(N__24569),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__4838 (
            .O(N__24564),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__4837 (
            .O(N__24557),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    CascadeMux I__4836 (
            .O(N__24542),
            .I(N__24539));
    InMux I__4835 (
            .O(N__24539),
            .I(N__24536));
    LocalMux I__4834 (
            .O(N__24536),
            .I(\POWERLED.un1_dutycycle_53_50_3_0 ));
    CascadeMux I__4833 (
            .O(N__24533),
            .I(N__24529));
    InMux I__4832 (
            .O(N__24532),
            .I(N__24526));
    InMux I__4831 (
            .O(N__24529),
            .I(N__24523));
    LocalMux I__4830 (
            .O(N__24526),
            .I(N__24520));
    LocalMux I__4829 (
            .O(N__24523),
            .I(N__24517));
    Span4Mux_s2_v I__4828 (
            .O(N__24520),
            .I(N__24512));
    Span4Mux_s2_v I__4827 (
            .O(N__24517),
            .I(N__24512));
    Odrv4 I__4826 (
            .O(N__24512),
            .I(\VPP_VDDQ.N_64_i ));
    InMux I__4825 (
            .O(N__24509),
            .I(N__24505));
    InMux I__4824 (
            .O(N__24508),
            .I(N__24502));
    LocalMux I__4823 (
            .O(N__24505),
            .I(N__24499));
    LocalMux I__4822 (
            .O(N__24502),
            .I(N__24494));
    Span4Mux_s1_v I__4821 (
            .O(N__24499),
            .I(N__24494));
    Odrv4 I__4820 (
            .O(N__24494),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    InMux I__4819 (
            .O(N__24491),
            .I(N__24488));
    LocalMux I__4818 (
            .O(N__24488),
            .I(\POWERLED.un1_dutycycle_53_45_0 ));
    InMux I__4817 (
            .O(N__24485),
            .I(N__24482));
    LocalMux I__4816 (
            .O(N__24482),
            .I(N__24479));
    Odrv4 I__4815 (
            .O(N__24479),
            .I(\POWERLED.dutycycle_RNIZ0Z_4 ));
    CascadeMux I__4814 (
            .O(N__24476),
            .I(\POWERLED.un1_dutycycle_53_35_1_cascade_ ));
    InMux I__4813 (
            .O(N__24473),
            .I(N__24469));
    InMux I__4812 (
            .O(N__24472),
            .I(N__24464));
    LocalMux I__4811 (
            .O(N__24469),
            .I(N__24461));
    InMux I__4810 (
            .O(N__24468),
            .I(N__24456));
    InMux I__4809 (
            .O(N__24467),
            .I(N__24456));
    LocalMux I__4808 (
            .O(N__24464),
            .I(\POWERLED.un1_dutycycle_53_22 ));
    Odrv4 I__4807 (
            .O(N__24461),
            .I(\POWERLED.un1_dutycycle_53_22 ));
    LocalMux I__4806 (
            .O(N__24456),
            .I(\POWERLED.un1_dutycycle_53_22 ));
    InMux I__4805 (
            .O(N__24449),
            .I(N__24446));
    LocalMux I__4804 (
            .O(N__24446),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_6 ));
    InMux I__4803 (
            .O(N__24443),
            .I(N__24438));
    InMux I__4802 (
            .O(N__24442),
            .I(N__24435));
    InMux I__4801 (
            .O(N__24441),
            .I(N__24431));
    LocalMux I__4800 (
            .O(N__24438),
            .I(N__24428));
    LocalMux I__4799 (
            .O(N__24435),
            .I(N__24422));
    InMux I__4798 (
            .O(N__24434),
            .I(N__24419));
    LocalMux I__4797 (
            .O(N__24431),
            .I(N__24416));
    Span4Mux_s3_v I__4796 (
            .O(N__24428),
            .I(N__24413));
    InMux I__4795 (
            .O(N__24427),
            .I(N__24410));
    InMux I__4794 (
            .O(N__24426),
            .I(N__24407));
    InMux I__4793 (
            .O(N__24425),
            .I(N__24404));
    Span4Mux_s1_v I__4792 (
            .O(N__24422),
            .I(N__24397));
    LocalMux I__4791 (
            .O(N__24419),
            .I(N__24397));
    Span4Mux_h I__4790 (
            .O(N__24416),
            .I(N__24397));
    Odrv4 I__4789 (
            .O(N__24413),
            .I(\POWERLED.dutycycle_RNI_10_8 ));
    LocalMux I__4788 (
            .O(N__24410),
            .I(\POWERLED.dutycycle_RNI_10_8 ));
    LocalMux I__4787 (
            .O(N__24407),
            .I(\POWERLED.dutycycle_RNI_10_8 ));
    LocalMux I__4786 (
            .O(N__24404),
            .I(\POWERLED.dutycycle_RNI_10_8 ));
    Odrv4 I__4785 (
            .O(N__24397),
            .I(\POWERLED.dutycycle_RNI_10_8 ));
    InMux I__4784 (
            .O(N__24386),
            .I(N__24383));
    LocalMux I__4783 (
            .O(N__24383),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_6 ));
    CascadeMux I__4782 (
            .O(N__24380),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_6_cascade_ ));
    InMux I__4781 (
            .O(N__24377),
            .I(N__24371));
    InMux I__4780 (
            .O(N__24376),
            .I(N__24371));
    LocalMux I__4779 (
            .O(N__24371),
            .I(\POWERLED.un1_dutycycle_53_35_1 ));
    CascadeMux I__4778 (
            .O(N__24368),
            .I(N__24365));
    InMux I__4777 (
            .O(N__24365),
            .I(N__24361));
    InMux I__4776 (
            .O(N__24364),
            .I(N__24358));
    LocalMux I__4775 (
            .O(N__24361),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_6 ));
    LocalMux I__4774 (
            .O(N__24358),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_6 ));
    CascadeMux I__4773 (
            .O(N__24353),
            .I(N__24350));
    InMux I__4772 (
            .O(N__24350),
            .I(N__24345));
    InMux I__4771 (
            .O(N__24349),
            .I(N__24340));
    InMux I__4770 (
            .O(N__24348),
            .I(N__24340));
    LocalMux I__4769 (
            .O(N__24345),
            .I(\POWERLED.un1_dutycycle_53_50_a0_0 ));
    LocalMux I__4768 (
            .O(N__24340),
            .I(\POWERLED.un1_dutycycle_53_50_a0_0 ));
    CascadeMux I__4767 (
            .O(N__24335),
            .I(\POWERLED.un1_dutycycle_53_50_a0_0_cascade_ ));
    InMux I__4766 (
            .O(N__24332),
            .I(N__24329));
    LocalMux I__4765 (
            .O(N__24329),
            .I(\POWERLED.un1_dutycycle_53_50_a0_0_0 ));
    InMux I__4764 (
            .O(N__24326),
            .I(N__24323));
    LocalMux I__4763 (
            .O(N__24323),
            .I(\POWERLED.un1_dutycycle_53_9_4_0 ));
    InMux I__4762 (
            .O(N__24320),
            .I(N__24317));
    LocalMux I__4761 (
            .O(N__24317),
            .I(\POWERLED.un1_dutycycle_53_9_4_1 ));
    InMux I__4760 (
            .O(N__24314),
            .I(N__24310));
    InMux I__4759 (
            .O(N__24313),
            .I(N__24307));
    LocalMux I__4758 (
            .O(N__24310),
            .I(N__24302));
    LocalMux I__4757 (
            .O(N__24307),
            .I(N__24302));
    Odrv4 I__4756 (
            .O(N__24302),
            .I(\POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0 ));
    CascadeMux I__4755 (
            .O(N__24299),
            .I(N__24295));
    InMux I__4754 (
            .O(N__24298),
            .I(N__24290));
    InMux I__4753 (
            .O(N__24295),
            .I(N__24290));
    LocalMux I__4752 (
            .O(N__24290),
            .I(N__24287));
    Odrv4 I__4751 (
            .O(N__24287),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    CascadeMux I__4750 (
            .O(N__24284),
            .I(\POWERLED.dutycycleZ0Z_7_cascade_ ));
    CascadeMux I__4749 (
            .O(N__24281),
            .I(\POWERLED.un1_dutycycle_53_9_a0_0_cascade_ ));
    CascadeMux I__4748 (
            .O(N__24278),
            .I(N__24275));
    InMux I__4747 (
            .O(N__24275),
            .I(N__24272));
    LocalMux I__4746 (
            .O(N__24272),
            .I(N__24269));
    Odrv4 I__4745 (
            .O(N__24269),
            .I(\POWERLED.un1_dutycycle_53_10_4 ));
    InMux I__4744 (
            .O(N__24266),
            .I(N__24263));
    LocalMux I__4743 (
            .O(N__24263),
            .I(\POWERLED.un1_dutycycle_53_40_0 ));
    CascadeMux I__4742 (
            .O(N__24260),
            .I(\POWERLED.un1_dutycycle_53_axb_11_1_cascade_ ));
    CascadeMux I__4741 (
            .O(N__24257),
            .I(\POWERLED.un1_dutycycle_53_axb_11_cascade_ ));
    CascadeMux I__4740 (
            .O(N__24254),
            .I(N__24251));
    InMux I__4739 (
            .O(N__24251),
            .I(N__24248));
    LocalMux I__4738 (
            .O(N__24248),
            .I(N__24245));
    Odrv4 I__4737 (
            .O(N__24245),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_14 ));
    CascadeMux I__4736 (
            .O(N__24242),
            .I(\POWERLED.dutycycleZ0Z_5_cascade_ ));
    InMux I__4735 (
            .O(N__24239),
            .I(N__24236));
    LocalMux I__4734 (
            .O(N__24236),
            .I(\POWERLED.dutycycle_RNIF86R3Z0Z_4 ));
    InMux I__4733 (
            .O(N__24233),
            .I(N__24230));
    LocalMux I__4732 (
            .O(N__24230),
            .I(\POWERLED.dutycycle_RNIP1UTZ0Z_4 ));
    CascadeMux I__4731 (
            .O(N__24227),
            .I(\POWERLED.dutycycle_RNIF86R3Z0Z_4_cascade_ ));
    InMux I__4730 (
            .O(N__24224),
            .I(N__24215));
    InMux I__4729 (
            .O(N__24223),
            .I(N__24215));
    InMux I__4728 (
            .O(N__24222),
            .I(N__24215));
    LocalMux I__4727 (
            .O(N__24215),
            .I(\POWERLED.dutycycleZ1Z_4 ));
    CascadeMux I__4726 (
            .O(N__24212),
            .I(\POWERLED.un1_dutycycle_53_31_0_0_cascade_ ));
    InMux I__4725 (
            .O(N__24209),
            .I(N__24206));
    LocalMux I__4724 (
            .O(N__24206),
            .I(\POWERLED.un1_dutycycle_53_9_3 ));
    CascadeMux I__4723 (
            .O(N__24203),
            .I(N__24200));
    InMux I__4722 (
            .O(N__24200),
            .I(N__24197));
    LocalMux I__4721 (
            .O(N__24197),
            .I(N__24194));
    Span4Mux_h I__4720 (
            .O(N__24194),
            .I(N__24191));
    Odrv4 I__4719 (
            .O(N__24191),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_11 ));
    InMux I__4718 (
            .O(N__24188),
            .I(N__24182));
    InMux I__4717 (
            .O(N__24187),
            .I(N__24182));
    LocalMux I__4716 (
            .O(N__24182),
            .I(\POWERLED.dutycycleZ1Z_8 ));
    CascadeMux I__4715 (
            .O(N__24179),
            .I(N__24176));
    InMux I__4714 (
            .O(N__24176),
            .I(N__24170));
    InMux I__4713 (
            .O(N__24175),
            .I(N__24170));
    LocalMux I__4712 (
            .O(N__24170),
            .I(N__24167));
    Odrv4 I__4711 (
            .O(N__24167),
            .I(\POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ));
    InMux I__4710 (
            .O(N__24164),
            .I(N__24158));
    InMux I__4709 (
            .O(N__24163),
            .I(N__24158));
    LocalMux I__4708 (
            .O(N__24158),
            .I(N__24155));
    Span4Mux_v I__4707 (
            .O(N__24155),
            .I(N__24152));
    Odrv4 I__4706 (
            .O(N__24152),
            .I(\POWERLED.dutycycle_RNIRT5H5Z0Z_8 ));
    CascadeMux I__4705 (
            .O(N__24149),
            .I(\POWERLED.dutycycleZ0Z_3_cascade_ ));
    CascadeMux I__4704 (
            .O(N__24146),
            .I(\POWERLED.dutycycle_RNI_10_8_cascade_ ));
    InMux I__4703 (
            .O(N__24143),
            .I(N__24140));
    LocalMux I__4702 (
            .O(N__24140),
            .I(\POWERLED.un1_dutycycle_53_9_4 ));
    InMux I__4701 (
            .O(N__24137),
            .I(N__24131));
    InMux I__4700 (
            .O(N__24136),
            .I(N__24131));
    LocalMux I__4699 (
            .O(N__24131),
            .I(N__24128));
    Span4Mux_v I__4698 (
            .O(N__24128),
            .I(N__24125));
    Odrv4 I__4697 (
            .O(N__24125),
            .I(\POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0 ));
    InMux I__4696 (
            .O(N__24122),
            .I(\POWERLED.un1_dutycycle_94_cry_10 ));
    InMux I__4695 (
            .O(N__24119),
            .I(\POWERLED.un1_dutycycle_94_cry_11_cZ0 ));
    InMux I__4694 (
            .O(N__24116),
            .I(N__24108));
    InMux I__4693 (
            .O(N__24115),
            .I(N__24103));
    InMux I__4692 (
            .O(N__24114),
            .I(N__24103));
    InMux I__4691 (
            .O(N__24113),
            .I(N__24098));
    InMux I__4690 (
            .O(N__24112),
            .I(N__24098));
    InMux I__4689 (
            .O(N__24111),
            .I(N__24095));
    LocalMux I__4688 (
            .O(N__24108),
            .I(N__24090));
    LocalMux I__4687 (
            .O(N__24103),
            .I(N__24085));
    LocalMux I__4686 (
            .O(N__24098),
            .I(N__24085));
    LocalMux I__4685 (
            .O(N__24095),
            .I(N__24082));
    InMux I__4684 (
            .O(N__24094),
            .I(N__24079));
    InMux I__4683 (
            .O(N__24093),
            .I(N__24076));
    Span4Mux_h I__4682 (
            .O(N__24090),
            .I(N__24071));
    Span4Mux_s1_v I__4681 (
            .O(N__24085),
            .I(N__24071));
    Odrv4 I__4680 (
            .O(N__24082),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__4679 (
            .O(N__24079),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__4678 (
            .O(N__24076),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv4 I__4677 (
            .O(N__24071),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    InMux I__4676 (
            .O(N__24062),
            .I(N__24056));
    InMux I__4675 (
            .O(N__24061),
            .I(N__24056));
    LocalMux I__4674 (
            .O(N__24056),
            .I(N__24053));
    Span4Mux_h I__4673 (
            .O(N__24053),
            .I(N__24050));
    Odrv4 I__4672 (
            .O(N__24050),
            .I(\POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ));
    InMux I__4671 (
            .O(N__24047),
            .I(\POWERLED.un1_dutycycle_94_cry_12 ));
    CascadeMux I__4670 (
            .O(N__24044),
            .I(N__24033));
    CascadeMux I__4669 (
            .O(N__24043),
            .I(N__24030));
    CascadeMux I__4668 (
            .O(N__24042),
            .I(N__24026));
    CascadeMux I__4667 (
            .O(N__24041),
            .I(N__24023));
    CascadeMux I__4666 (
            .O(N__24040),
            .I(N__24018));
    CascadeMux I__4665 (
            .O(N__24039),
            .I(N__24015));
    CascadeMux I__4664 (
            .O(N__24038),
            .I(N__24011));
    CascadeMux I__4663 (
            .O(N__24037),
            .I(N__24007));
    CascadeMux I__4662 (
            .O(N__24036),
            .I(N__24004));
    InMux I__4661 (
            .O(N__24033),
            .I(N__23999));
    InMux I__4660 (
            .O(N__24030),
            .I(N__23999));
    InMux I__4659 (
            .O(N__24029),
            .I(N__23994));
    InMux I__4658 (
            .O(N__24026),
            .I(N__23994));
    InMux I__4657 (
            .O(N__24023),
            .I(N__23983));
    InMux I__4656 (
            .O(N__24022),
            .I(N__23983));
    InMux I__4655 (
            .O(N__24021),
            .I(N__23983));
    InMux I__4654 (
            .O(N__24018),
            .I(N__23983));
    InMux I__4653 (
            .O(N__24015),
            .I(N__23983));
    InMux I__4652 (
            .O(N__24014),
            .I(N__23972));
    InMux I__4651 (
            .O(N__24011),
            .I(N__23972));
    InMux I__4650 (
            .O(N__24010),
            .I(N__23972));
    InMux I__4649 (
            .O(N__24007),
            .I(N__23972));
    InMux I__4648 (
            .O(N__24004),
            .I(N__23972));
    LocalMux I__4647 (
            .O(N__23999),
            .I(N__23963));
    LocalMux I__4646 (
            .O(N__23994),
            .I(N__23963));
    LocalMux I__4645 (
            .O(N__23983),
            .I(N__23963));
    LocalMux I__4644 (
            .O(N__23972),
            .I(N__23963));
    Odrv4 I__4643 (
            .O(N__23963),
            .I(\POWERLED.N_435_i ));
    CascadeMux I__4642 (
            .O(N__23960),
            .I(N__23957));
    InMux I__4641 (
            .O(N__23957),
            .I(N__23951));
    InMux I__4640 (
            .O(N__23956),
            .I(N__23951));
    LocalMux I__4639 (
            .O(N__23951),
            .I(N__23948));
    Span4Mux_s3_v I__4638 (
            .O(N__23948),
            .I(N__23945));
    Odrv4 I__4637 (
            .O(N__23945),
            .I(\POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ));
    InMux I__4636 (
            .O(N__23942),
            .I(\POWERLED.un1_dutycycle_94_cry_13_cZ0 ));
    InMux I__4635 (
            .O(N__23939),
            .I(\POWERLED.un1_dutycycle_94_cry_14 ));
    CascadeMux I__4634 (
            .O(N__23936),
            .I(N__23932));
    InMux I__4633 (
            .O(N__23935),
            .I(N__23927));
    InMux I__4632 (
            .O(N__23932),
            .I(N__23927));
    LocalMux I__4631 (
            .O(N__23927),
            .I(N__23924));
    Span4Mux_s2_v I__4630 (
            .O(N__23924),
            .I(N__23921));
    Odrv4 I__4629 (
            .O(N__23921),
            .I(\POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ));
    IoInMux I__4628 (
            .O(N__23918),
            .I(N__23915));
    LocalMux I__4627 (
            .O(N__23915),
            .I(N__23912));
    IoSpan4Mux I__4626 (
            .O(N__23912),
            .I(N__23909));
    Span4Mux_s3_h I__4625 (
            .O(N__23909),
            .I(N__23906));
    Span4Mux_h I__4624 (
            .O(N__23906),
            .I(N__23903));
    Odrv4 I__4623 (
            .O(N__23903),
            .I(vccst_en));
    CascadeMux I__4622 (
            .O(N__23900),
            .I(N__23897));
    InMux I__4621 (
            .O(N__23897),
            .I(N__23894));
    LocalMux I__4620 (
            .O(N__23894),
            .I(N__23891));
    Odrv4 I__4619 (
            .O(N__23891),
            .I(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ));
    CascadeMux I__4618 (
            .O(N__23888),
            .I(\POWERLED.dutycycle_RNIP1UTZ0Z_4_cascade_ ));
    CascadeMux I__4617 (
            .O(N__23885),
            .I(N__23882));
    InMux I__4616 (
            .O(N__23882),
            .I(N__23879));
    LocalMux I__4615 (
            .O(N__23879),
            .I(\POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ));
    InMux I__4614 (
            .O(N__23876),
            .I(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ));
    InMux I__4613 (
            .O(N__23873),
            .I(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ));
    InMux I__4612 (
            .O(N__23870),
            .I(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ));
    InMux I__4611 (
            .O(N__23867),
            .I(\POWERLED.un1_dutycycle_94_cry_4 ));
    InMux I__4610 (
            .O(N__23864),
            .I(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ));
    InMux I__4609 (
            .O(N__23861),
            .I(N__23858));
    LocalMux I__4608 (
            .O(N__23858),
            .I(\POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ));
    InMux I__4607 (
            .O(N__23855),
            .I(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ));
    InMux I__4606 (
            .O(N__23852),
            .I(bfn_9_11_0_));
    InMux I__4605 (
            .O(N__23849),
            .I(N__23843));
    InMux I__4604 (
            .O(N__23848),
            .I(N__23843));
    LocalMux I__4603 (
            .O(N__23843),
            .I(N__23840));
    Odrv4 I__4602 (
            .O(N__23840),
            .I(\POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61 ));
    InMux I__4601 (
            .O(N__23837),
            .I(\POWERLED.un1_dutycycle_94_cry_8 ));
    InMux I__4600 (
            .O(N__23834),
            .I(\POWERLED.un1_dutycycle_94_cry_9 ));
    CascadeMux I__4599 (
            .O(N__23831),
            .I(N__23828));
    InMux I__4598 (
            .O(N__23828),
            .I(N__23825));
    LocalMux I__4597 (
            .O(N__23825),
            .I(\POWERLED.func_state_1_m2s2_i_0_a2_1_0 ));
    CascadeMux I__4596 (
            .O(N__23822),
            .I(\POWERLED.un1_dutycycle_96_0_a3_0_a2_1_cascade_ ));
    InMux I__4595 (
            .O(N__23819),
            .I(N__23816));
    LocalMux I__4594 (
            .O(N__23816),
            .I(N__23812));
    InMux I__4593 (
            .O(N__23815),
            .I(N__23809));
    Odrv4 I__4592 (
            .O(N__23812),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_3 ));
    LocalMux I__4591 (
            .O(N__23809),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_3 ));
    CascadeMux I__4590 (
            .O(N__23804),
            .I(\POWERLED.N_251_cascade_ ));
    InMux I__4589 (
            .O(N__23801),
            .I(N__23798));
    LocalMux I__4588 (
            .O(N__23798),
            .I(N__23795));
    Odrv4 I__4587 (
            .O(N__23795),
            .I(\POWERLED.N_506 ));
    InMux I__4586 (
            .O(N__23792),
            .I(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ));
    CascadeMux I__4585 (
            .O(N__23789),
            .I(\POWERLED.N_448_cascade_ ));
    InMux I__4584 (
            .O(N__23786),
            .I(N__23783));
    LocalMux I__4583 (
            .O(N__23783),
            .I(N__23780));
    Odrv4 I__4582 (
            .O(N__23780),
            .I(\POWERLED.N_656_0 ));
    CascadeMux I__4581 (
            .O(N__23777),
            .I(\POWERLED.N_133_cascade_ ));
    InMux I__4580 (
            .O(N__23774),
            .I(N__23771));
    LocalMux I__4579 (
            .O(N__23771),
            .I(\POWERLED.un1_dutycycle_172_m4 ));
    InMux I__4578 (
            .O(N__23768),
            .I(N__23765));
    LocalMux I__4577 (
            .O(N__23765),
            .I(N__23762));
    Odrv4 I__4576 (
            .O(N__23762),
            .I(\POWERLED.dutycycle_eena_14_c ));
    CascadeMux I__4575 (
            .O(N__23759),
            .I(\POWERLED.N_488_cascade_ ));
    InMux I__4574 (
            .O(N__23756),
            .I(N__23753));
    LocalMux I__4573 (
            .O(N__23753),
            .I(\POWERLED.un1_dutycycle_172_m2 ));
    CascadeMux I__4572 (
            .O(N__23750),
            .I(\POWERLED.un1_clk_100khz_30_and_i_0_0_sx_cascade_ ));
    InMux I__4571 (
            .O(N__23747),
            .I(N__23744));
    LocalMux I__4570 (
            .O(N__23744),
            .I(\POWERLED.un1_dutycycle_164_0_a3_0_a2_0 ));
    CascadeMux I__4569 (
            .O(N__23741),
            .I(\POWERLED.count_clkZ0Z_7_cascade_ ));
    InMux I__4568 (
            .O(N__23738),
            .I(N__23735));
    LocalMux I__4567 (
            .O(N__23735),
            .I(N__23732));
    Odrv4 I__4566 (
            .O(N__23732),
            .I(\POWERLED.un1_func_state25_6_0_o_N_4 ));
    InMux I__4565 (
            .O(N__23729),
            .I(N__23723));
    InMux I__4564 (
            .O(N__23728),
            .I(N__23723));
    LocalMux I__4563 (
            .O(N__23723),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_9_0 ));
    InMux I__4562 (
            .O(N__23720),
            .I(N__23717));
    LocalMux I__4561 (
            .O(N__23717),
            .I(\POWERLED.count_clk_0_7 ));
    CascadeMux I__4560 (
            .O(N__23714),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_5_cascade_ ));
    InMux I__4559 (
            .O(N__23711),
            .I(N__23708));
    LocalMux I__4558 (
            .O(N__23708),
            .I(N__23705));
    Odrv4 I__4557 (
            .O(N__23705),
            .I(\POWERLED.un1_dutycycle_172_m3 ));
    CascadeMux I__4556 (
            .O(N__23702),
            .I(\POWERLED.un1_clk_100khz_52_and_i_0_m2_ns_1_cascade_ ));
    InMux I__4555 (
            .O(N__23699),
            .I(N__23696));
    LocalMux I__4554 (
            .O(N__23696),
            .I(POWERLED_g2_1_0_0));
    InMux I__4553 (
            .O(N__23693),
            .I(N__23690));
    LocalMux I__4552 (
            .O(N__23690),
            .I(N__23687));
    Span4Mux_v I__4551 (
            .O(N__23687),
            .I(N__23684));
    Odrv4 I__4550 (
            .O(N__23684),
            .I(\POWERLED.N_74 ));
    CascadeMux I__4549 (
            .O(N__23681),
            .I(\POWERLED.N_4_0_cascade_ ));
    InMux I__4548 (
            .O(N__23678),
            .I(N__23672));
    InMux I__4547 (
            .O(N__23677),
            .I(N__23672));
    LocalMux I__4546 (
            .O(N__23672),
            .I(\POWERLED.func_state_1_m2_0_0_0 ));
    InMux I__4545 (
            .O(N__23669),
            .I(N__23666));
    LocalMux I__4544 (
            .O(N__23666),
            .I(\POWERLED.g1_0_0 ));
    InMux I__4543 (
            .O(N__23663),
            .I(N__23660));
    LocalMux I__4542 (
            .O(N__23660),
            .I(\POWERLED.func_state_1_m2_N_3_7_1 ));
    InMux I__4541 (
            .O(N__23657),
            .I(N__23649));
    InMux I__4540 (
            .O(N__23656),
            .I(N__23649));
    InMux I__4539 (
            .O(N__23655),
            .I(N__23644));
    InMux I__4538 (
            .O(N__23654),
            .I(N__23644));
    LocalMux I__4537 (
            .O(N__23649),
            .I(clk_100Khz_signalkeep_3_fast));
    LocalMux I__4536 (
            .O(N__23644),
            .I(clk_100Khz_signalkeep_3_fast));
    CascadeMux I__4535 (
            .O(N__23639),
            .I(N__23636));
    InMux I__4534 (
            .O(N__23636),
            .I(N__23633));
    LocalMux I__4533 (
            .O(N__23633),
            .I(\POWERLED.N_671_0 ));
    CascadeMux I__4532 (
            .O(N__23630),
            .I(G_7_i_a4_1_0_cascade_));
    InMux I__4531 (
            .O(N__23627),
            .I(N__23624));
    LocalMux I__4530 (
            .O(N__23624),
            .I(\RSMRST_PWRGD.G_7_i_0 ));
    CascadeMux I__4529 (
            .O(N__23621),
            .I(\POWERLED.N_533_cascade_ ));
    InMux I__4528 (
            .O(N__23618),
            .I(N__23615));
    LocalMux I__4527 (
            .O(N__23615),
            .I(\POWERLED.N_533 ));
    InMux I__4526 (
            .O(N__23612),
            .I(N__23609));
    LocalMux I__4525 (
            .O(N__23609),
            .I(\POWERLED.un1_clk_100khz_51_and_i_3_0_sx ));
    InMux I__4524 (
            .O(N__23606),
            .I(N__23603));
    LocalMux I__4523 (
            .O(N__23603),
            .I(N__23599));
    InMux I__4522 (
            .O(N__23602),
            .I(N__23596));
    Span4Mux_h I__4521 (
            .O(N__23599),
            .I(N__23593));
    LocalMux I__4520 (
            .O(N__23596),
            .I(\POWERLED.count_offZ0Z_4 ));
    Odrv4 I__4519 (
            .O(N__23593),
            .I(\POWERLED.count_offZ0Z_4 ));
    InMux I__4518 (
            .O(N__23588),
            .I(N__23584));
    InMux I__4517 (
            .O(N__23587),
            .I(N__23581));
    LocalMux I__4516 (
            .O(N__23584),
            .I(N__23576));
    LocalMux I__4515 (
            .O(N__23581),
            .I(N__23576));
    Span4Mux_h I__4514 (
            .O(N__23576),
            .I(N__23573));
    Odrv4 I__4513 (
            .O(N__23573),
            .I(\POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ));
    InMux I__4512 (
            .O(N__23570),
            .I(N__23567));
    LocalMux I__4511 (
            .O(N__23567),
            .I(\POWERLED.count_off_0_4 ));
    InMux I__4510 (
            .O(N__23564),
            .I(N__23558));
    InMux I__4509 (
            .O(N__23563),
            .I(N__23558));
    LocalMux I__4508 (
            .O(N__23558),
            .I(N__23555));
    Odrv4 I__4507 (
            .O(N__23555),
            .I(\POWERLED.count_off_RNIZ0Z_1 ));
    InMux I__4506 (
            .O(N__23552),
            .I(N__23549));
    LocalMux I__4505 (
            .O(N__23549),
            .I(\POWERLED.count_off_0_1 ));
    CEMux I__4504 (
            .O(N__23546),
            .I(N__23534));
    CEMux I__4503 (
            .O(N__23545),
            .I(N__23531));
    InMux I__4502 (
            .O(N__23544),
            .I(N__23522));
    InMux I__4501 (
            .O(N__23543),
            .I(N__23522));
    InMux I__4500 (
            .O(N__23542),
            .I(N__23522));
    InMux I__4499 (
            .O(N__23541),
            .I(N__23522));
    CascadeMux I__4498 (
            .O(N__23540),
            .I(N__23515));
    CascadeMux I__4497 (
            .O(N__23539),
            .I(N__23512));
    CEMux I__4496 (
            .O(N__23538),
            .I(N__23508));
    CEMux I__4495 (
            .O(N__23537),
            .I(N__23505));
    LocalMux I__4494 (
            .O(N__23534),
            .I(N__23502));
    LocalMux I__4493 (
            .O(N__23531),
            .I(N__23499));
    LocalMux I__4492 (
            .O(N__23522),
            .I(N__23496));
    InMux I__4491 (
            .O(N__23521),
            .I(N__23491));
    InMux I__4490 (
            .O(N__23520),
            .I(N__23491));
    CEMux I__4489 (
            .O(N__23519),
            .I(N__23480));
    CEMux I__4488 (
            .O(N__23518),
            .I(N__23477));
    InMux I__4487 (
            .O(N__23515),
            .I(N__23474));
    InMux I__4486 (
            .O(N__23512),
            .I(N__23469));
    InMux I__4485 (
            .O(N__23511),
            .I(N__23469));
    LocalMux I__4484 (
            .O(N__23508),
            .I(N__23466));
    LocalMux I__4483 (
            .O(N__23505),
            .I(N__23461));
    Span4Mux_s2_v I__4482 (
            .O(N__23502),
            .I(N__23461));
    Span4Mux_s2_v I__4481 (
            .O(N__23499),
            .I(N__23456));
    Span4Mux_s2_v I__4480 (
            .O(N__23496),
            .I(N__23456));
    LocalMux I__4479 (
            .O(N__23491),
            .I(N__23453));
    InMux I__4478 (
            .O(N__23490),
            .I(N__23442));
    CEMux I__4477 (
            .O(N__23489),
            .I(N__23442));
    InMux I__4476 (
            .O(N__23488),
            .I(N__23442));
    InMux I__4475 (
            .O(N__23487),
            .I(N__23442));
    InMux I__4474 (
            .O(N__23486),
            .I(N__23442));
    InMux I__4473 (
            .O(N__23485),
            .I(N__23435));
    InMux I__4472 (
            .O(N__23484),
            .I(N__23435));
    InMux I__4471 (
            .O(N__23483),
            .I(N__23435));
    LocalMux I__4470 (
            .O(N__23480),
            .I(N__23432));
    LocalMux I__4469 (
            .O(N__23477),
            .I(N__23429));
    LocalMux I__4468 (
            .O(N__23474),
            .I(N__23424));
    LocalMux I__4467 (
            .O(N__23469),
            .I(N__23424));
    Span4Mux_v I__4466 (
            .O(N__23466),
            .I(N__23415));
    Span4Mux_v I__4465 (
            .O(N__23461),
            .I(N__23415));
    Span4Mux_v I__4464 (
            .O(N__23456),
            .I(N__23415));
    Span4Mux_v I__4463 (
            .O(N__23453),
            .I(N__23415));
    LocalMux I__4462 (
            .O(N__23442),
            .I(N__23410));
    LocalMux I__4461 (
            .O(N__23435),
            .I(N__23410));
    Span4Mux_s3_h I__4460 (
            .O(N__23432),
            .I(N__23403));
    Span4Mux_s3_v I__4459 (
            .O(N__23429),
            .I(N__23403));
    Span4Mux_s3_h I__4458 (
            .O(N__23424),
            .I(N__23403));
    Odrv4 I__4457 (
            .O(N__23415),
            .I(\POWERLED.func_state_RNI7LSV8Z0Z_0 ));
    Odrv12 I__4456 (
            .O(N__23410),
            .I(\POWERLED.func_state_RNI7LSV8Z0Z_0 ));
    Odrv4 I__4455 (
            .O(N__23403),
            .I(\POWERLED.func_state_RNI7LSV8Z0Z_0 ));
    InMux I__4454 (
            .O(N__23396),
            .I(N__23393));
    LocalMux I__4453 (
            .O(N__23393),
            .I(N__23388));
    InMux I__4452 (
            .O(N__23392),
            .I(N__23383));
    InMux I__4451 (
            .O(N__23391),
            .I(N__23383));
    Span4Mux_h I__4450 (
            .O(N__23388),
            .I(N__23380));
    LocalMux I__4449 (
            .O(N__23383),
            .I(N__23377));
    Odrv4 I__4448 (
            .O(N__23380),
            .I(\POWERLED.count_offZ0Z_1 ));
    Odrv4 I__4447 (
            .O(N__23377),
            .I(\POWERLED.count_offZ0Z_1 ));
    CascadeMux I__4446 (
            .O(N__23372),
            .I(N_7_cascade_));
    CascadeMux I__4445 (
            .O(N__23369),
            .I(N_8_0_cascade_));
    CascadeMux I__4444 (
            .O(N__23366),
            .I(\POWERLED.g0_5Z0Z_1_cascade_ ));
    CascadeMux I__4443 (
            .O(N__23363),
            .I(\POWERLED.G_30Z0Z_0_cascade_ ));
    InMux I__4442 (
            .O(N__23360),
            .I(N__23356));
    InMux I__4441 (
            .O(N__23359),
            .I(N__23353));
    LocalMux I__4440 (
            .O(N__23356),
            .I(VPP_VDDQ_un6_count));
    LocalMux I__4439 (
            .O(N__23353),
            .I(VPP_VDDQ_un6_count));
    CascadeMux I__4438 (
            .O(N__23348),
            .I(G_30_cascade_));
    InMux I__4437 (
            .O(N__23345),
            .I(N__23342));
    LocalMux I__4436 (
            .O(N__23342),
            .I(N__23335));
    InMux I__4435 (
            .O(N__23341),
            .I(N__23326));
    InMux I__4434 (
            .O(N__23340),
            .I(N__23326));
    InMux I__4433 (
            .O(N__23339),
            .I(N__23326));
    InMux I__4432 (
            .O(N__23338),
            .I(N__23326));
    Span4Mux_v I__4431 (
            .O(N__23335),
            .I(N__23323));
    LocalMux I__4430 (
            .O(N__23326),
            .I(N__23320));
    Span4Mux_h I__4429 (
            .O(N__23323),
            .I(N__23315));
    Span4Mux_s3_h I__4428 (
            .O(N__23320),
            .I(N__23315));
    Odrv4 I__4427 (
            .O(N__23315),
            .I(N_626));
    InMux I__4426 (
            .O(N__23312),
            .I(N__23306));
    InMux I__4425 (
            .O(N__23311),
            .I(N__23306));
    LocalMux I__4424 (
            .O(N__23306),
            .I(N__23303));
    Span4Mux_h I__4423 (
            .O(N__23303),
            .I(N__23298));
    CascadeMux I__4422 (
            .O(N__23302),
            .I(N__23293));
    CascadeMux I__4421 (
            .O(N__23301),
            .I(N__23290));
    Span4Mux_h I__4420 (
            .O(N__23298),
            .I(N__23286));
    InMux I__4419 (
            .O(N__23297),
            .I(N__23283));
    InMux I__4418 (
            .O(N__23296),
            .I(N__23274));
    InMux I__4417 (
            .O(N__23293),
            .I(N__23274));
    InMux I__4416 (
            .O(N__23290),
            .I(N__23274));
    InMux I__4415 (
            .O(N__23289),
            .I(N__23274));
    Odrv4 I__4414 (
            .O(N__23286),
            .I(VPP_VDDQ_curr_state_1));
    LocalMux I__4413 (
            .O(N__23283),
            .I(VPP_VDDQ_curr_state_1));
    LocalMux I__4412 (
            .O(N__23274),
            .I(VPP_VDDQ_curr_state_1));
    CascadeMux I__4411 (
            .O(N__23267),
            .I(N__23264));
    InMux I__4410 (
            .O(N__23264),
            .I(N__23261));
    LocalMux I__4409 (
            .O(N__23261),
            .I(N__23258));
    Span4Mux_h I__4408 (
            .O(N__23258),
            .I(N__23255));
    Span4Mux_h I__4407 (
            .O(N__23255),
            .I(N__23248));
    InMux I__4406 (
            .O(N__23254),
            .I(N__23239));
    InMux I__4405 (
            .O(N__23253),
            .I(N__23239));
    InMux I__4404 (
            .O(N__23252),
            .I(N__23239));
    InMux I__4403 (
            .O(N__23251),
            .I(N__23239));
    Odrv4 I__4402 (
            .O(N__23248),
            .I(VPP_VDDQ_curr_state_0));
    LocalMux I__4401 (
            .O(N__23239),
            .I(VPP_VDDQ_curr_state_0));
    InMux I__4400 (
            .O(N__23234),
            .I(N__23231));
    LocalMux I__4399 (
            .O(N__23231),
            .I(\POWERLED.count_off_0_3 ));
    CascadeMux I__4398 (
            .O(N__23228),
            .I(N__23225));
    InMux I__4397 (
            .O(N__23225),
            .I(N__23219));
    InMux I__4396 (
            .O(N__23224),
            .I(N__23219));
    LocalMux I__4395 (
            .O(N__23219),
            .I(N__23216));
    Span4Mux_h I__4394 (
            .O(N__23216),
            .I(N__23213));
    Odrv4 I__4393 (
            .O(N__23213),
            .I(\POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ));
    InMux I__4392 (
            .O(N__23210),
            .I(N__23207));
    LocalMux I__4391 (
            .O(N__23207),
            .I(N__23204));
    Span4Mux_s3_v I__4390 (
            .O(N__23204),
            .I(N__23201));
    Odrv4 I__4389 (
            .O(N__23201),
            .I(\POWERLED.count_offZ0Z_3 ));
    InMux I__4388 (
            .O(N__23198),
            .I(N__23195));
    LocalMux I__4387 (
            .O(N__23195),
            .I(N__23192));
    Span4Mux_v I__4386 (
            .O(N__23192),
            .I(N__23188));
    InMux I__4385 (
            .O(N__23191),
            .I(N__23185));
    Span4Mux_v I__4384 (
            .O(N__23188),
            .I(N__23182));
    LocalMux I__4383 (
            .O(N__23185),
            .I(N__23179));
    Odrv4 I__4382 (
            .O(N__23182),
            .I(\POWERLED.count_offZ0Z_7 ));
    Odrv12 I__4381 (
            .O(N__23179),
            .I(\POWERLED.count_offZ0Z_7 ));
    CascadeMux I__4380 (
            .O(N__23174),
            .I(\POWERLED.count_offZ0Z_3_cascade_ ));
    InMux I__4379 (
            .O(N__23171),
            .I(N__23168));
    LocalMux I__4378 (
            .O(N__23168),
            .I(N__23164));
    InMux I__4377 (
            .O(N__23167),
            .I(N__23161));
    Span4Mux_v I__4376 (
            .O(N__23164),
            .I(N__23158));
    LocalMux I__4375 (
            .O(N__23161),
            .I(N__23155));
    Span4Mux_v I__4374 (
            .O(N__23158),
            .I(N__23152));
    Span4Mux_v I__4373 (
            .O(N__23155),
            .I(N__23149));
    Odrv4 I__4372 (
            .O(N__23152),
            .I(\POWERLED.count_offZ0Z_8 ));
    Odrv4 I__4371 (
            .O(N__23149),
            .I(\POWERLED.count_offZ0Z_8 ));
    InMux I__4370 (
            .O(N__23144),
            .I(N__23141));
    LocalMux I__4369 (
            .O(N__23141),
            .I(\POWERLED.un34_clk_100khz_10 ));
    InMux I__4368 (
            .O(N__23138),
            .I(N__23135));
    LocalMux I__4367 (
            .O(N__23135),
            .I(N__23132));
    Span12Mux_s5_h I__4366 (
            .O(N__23132),
            .I(N__23129));
    Odrv12 I__4365 (
            .O(N__23129),
            .I(\POWERLED.un34_clk_100khz_11 ));
    CascadeMux I__4364 (
            .O(N__23126),
            .I(\POWERLED.un34_clk_100khz_8_cascade_ ));
    InMux I__4363 (
            .O(N__23123),
            .I(N__23120));
    LocalMux I__4362 (
            .O(N__23120),
            .I(N__23117));
    Odrv4 I__4361 (
            .O(N__23117),
            .I(\POWERLED.un34_clk_100khz_9 ));
    CascadeMux I__4360 (
            .O(N__23114),
            .I(\POWERLED.dutycycleZ0Z_9_cascade_ ));
    CascadeMux I__4359 (
            .O(N__23111),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_11_cascade_ ));
    CascadeMux I__4358 (
            .O(N__23108),
            .I(N__23105));
    InMux I__4357 (
            .O(N__23105),
            .I(N__23102));
    LocalMux I__4356 (
            .O(N__23102),
            .I(\POWERLED.un1_dutycycle_53_2_1 ));
    CascadeMux I__4355 (
            .O(N__23099),
            .I(\POWERLED.un1_dutycycle_53_2_1_cascade_ ));
    InMux I__4354 (
            .O(N__23096),
            .I(N__23090));
    InMux I__4353 (
            .O(N__23095),
            .I(N__23090));
    LocalMux I__4352 (
            .O(N__23090),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_13 ));
    CascadeMux I__4351 (
            .O(N__23087),
            .I(\VPP_VDDQ.un6_count_8_cascade_ ));
    InMux I__4350 (
            .O(N__23084),
            .I(N__23081));
    LocalMux I__4349 (
            .O(N__23081),
            .I(\VPP_VDDQ.un6_count_10 ));
    InMux I__4348 (
            .O(N__23078),
            .I(N__23075));
    LocalMux I__4347 (
            .O(N__23075),
            .I(\VPP_VDDQ.un6_count_11 ));
    InMux I__4346 (
            .O(N__23072),
            .I(N__23069));
    LocalMux I__4345 (
            .O(N__23069),
            .I(\VPP_VDDQ.un6_count_9 ));
    CascadeMux I__4344 (
            .O(N__23066),
            .I(\POWERLED.dutycycle_RNI_12Z0Z_8_cascade_ ));
    CascadeMux I__4343 (
            .O(N__23063),
            .I(N__23060));
    InMux I__4342 (
            .O(N__23060),
            .I(N__23057));
    LocalMux I__4341 (
            .O(N__23057),
            .I(\POWERLED.dutycycle_RNIZ0Z_15 ));
    CascadeMux I__4340 (
            .O(N__23054),
            .I(N__23051));
    InMux I__4339 (
            .O(N__23051),
            .I(N__23045));
    InMux I__4338 (
            .O(N__23050),
            .I(N__23045));
    LocalMux I__4337 (
            .O(N__23045),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    CascadeMux I__4336 (
            .O(N__23042),
            .I(\POWERLED.dutycycleZ0Z_14_cascade_ ));
    CascadeMux I__4335 (
            .O(N__23039),
            .I(\POWERLED.N_2381_i_cascade_ ));
    InMux I__4334 (
            .O(N__23036),
            .I(N__23033));
    LocalMux I__4333 (
            .O(N__23033),
            .I(\POWERLED.un2_count_clk_17_0_0_a2_0_5 ));
    InMux I__4332 (
            .O(N__23030),
            .I(N__23027));
    LocalMux I__4331 (
            .O(N__23027),
            .I(N__23024));
    Odrv4 I__4330 (
            .O(N__23024),
            .I(\POWERLED.dutycycle_RNIZ0Z_13 ));
    CascadeMux I__4329 (
            .O(N__23021),
            .I(N__23017));
    InMux I__4328 (
            .O(N__23020),
            .I(N__23012));
    InMux I__4327 (
            .O(N__23017),
            .I(N__23012));
    LocalMux I__4326 (
            .O(N__23012),
            .I(\POWERLED.dutycycleZ1Z_11 ));
    InMux I__4325 (
            .O(N__23009),
            .I(N__23003));
    InMux I__4324 (
            .O(N__23008),
            .I(N__23003));
    LocalMux I__4323 (
            .O(N__23003),
            .I(N__23000));
    Span4Mux_v I__4322 (
            .O(N__23000),
            .I(N__22997));
    Odrv4 I__4321 (
            .O(N__22997),
            .I(\POWERLED.dutycycle_en_7 ));
    CascadeMux I__4320 (
            .O(N__22994),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_8_cascade_ ));
    CascadeMux I__4319 (
            .O(N__22991),
            .I(\POWERLED.dutycycle_RNIZ0Z_6_cascade_ ));
    InMux I__4318 (
            .O(N__22988),
            .I(N__22985));
    LocalMux I__4317 (
            .O(N__22985),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_7 ));
    InMux I__4316 (
            .O(N__22982),
            .I(N__22979));
    LocalMux I__4315 (
            .O(N__22979),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_8 ));
    CascadeMux I__4314 (
            .O(N__22976),
            .I(N__22973));
    InMux I__4313 (
            .O(N__22973),
            .I(N__22970));
    LocalMux I__4312 (
            .O(N__22970),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_5 ));
    CascadeMux I__4311 (
            .O(N__22967),
            .I(\POWERLED.un1_dutycycle_53_31_a4_1_cascade_ ));
    InMux I__4310 (
            .O(N__22964),
            .I(N__22961));
    LocalMux I__4309 (
            .O(N__22961),
            .I(\POWERLED.un1_dutycycle_53_31_a5_1 ));
    InMux I__4308 (
            .O(N__22958),
            .I(N__22955));
    LocalMux I__4307 (
            .O(N__22955),
            .I(\POWERLED.un1_dutycycle_53_31_a0_2 ));
    CascadeMux I__4306 (
            .O(N__22952),
            .I(N__22949));
    InMux I__4305 (
            .O(N__22949),
            .I(N__22946));
    LocalMux I__4304 (
            .O(N__22946),
            .I(\POWERLED.dutycycle_RNIZ0Z_12 ));
    InMux I__4303 (
            .O(N__22943),
            .I(N__22937));
    InMux I__4302 (
            .O(N__22942),
            .I(N__22937));
    LocalMux I__4301 (
            .O(N__22937),
            .I(\POWERLED.dutycycleZ1Z_14 ));
    CascadeMux I__4300 (
            .O(N__22934),
            .I(N__22931));
    InMux I__4299 (
            .O(N__22931),
            .I(N__22925));
    InMux I__4298 (
            .O(N__22930),
            .I(N__22925));
    LocalMux I__4297 (
            .O(N__22925),
            .I(N__22922));
    Odrv4 I__4296 (
            .O(N__22922),
            .I(\POWERLED.dutycycle_en_10 ));
    CascadeMux I__4295 (
            .O(N__22919),
            .I(N__22916));
    InMux I__4294 (
            .O(N__22916),
            .I(N__22910));
    InMux I__4293 (
            .O(N__22915),
            .I(N__22910));
    LocalMux I__4292 (
            .O(N__22910),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    InMux I__4291 (
            .O(N__22907),
            .I(N__22904));
    LocalMux I__4290 (
            .O(N__22904),
            .I(\POWERLED.un1_dutycycle_53_41_0 ));
    CascadeMux I__4289 (
            .O(N__22901),
            .I(\POWERLED.un1_dutycycle_53_40_0_cascade_ ));
    CascadeMux I__4288 (
            .O(N__22898),
            .I(N__22895));
    InMux I__4287 (
            .O(N__22895),
            .I(N__22892));
    LocalMux I__4286 (
            .O(N__22892),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_13 ));
    CascadeMux I__4285 (
            .O(N__22889),
            .I(N__22885));
    CascadeMux I__4284 (
            .O(N__22888),
            .I(N__22882));
    InMux I__4283 (
            .O(N__22885),
            .I(N__22877));
    InMux I__4282 (
            .O(N__22882),
            .I(N__22877));
    LocalMux I__4281 (
            .O(N__22877),
            .I(\POWERLED.dutycycleZ1Z_9 ));
    CascadeMux I__4280 (
            .O(N__22874),
            .I(\POWERLED.dutycycleZ0Z_4_cascade_ ));
    InMux I__4279 (
            .O(N__22871),
            .I(N__22866));
    InMux I__4278 (
            .O(N__22870),
            .I(N__22863));
    InMux I__4277 (
            .O(N__22869),
            .I(N__22860));
    LocalMux I__4276 (
            .O(N__22866),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__4275 (
            .O(N__22863),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__4274 (
            .O(N__22860),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    CascadeMux I__4273 (
            .O(N__22853),
            .I(N__22850));
    InMux I__4272 (
            .O(N__22850),
            .I(N__22847));
    LocalMux I__4271 (
            .O(N__22847),
            .I(\POWERLED.mult1_un47_sum_l_fx_3 ));
    InMux I__4270 (
            .O(N__22844),
            .I(N__22841));
    LocalMux I__4269 (
            .O(N__22841),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_0 ));
    CascadeMux I__4268 (
            .O(N__22838),
            .I(\POWERLED.dutycycle_RNIZ0Z_3_cascade_ ));
    CascadeMux I__4267 (
            .O(N__22835),
            .I(N__22832));
    InMux I__4266 (
            .O(N__22832),
            .I(N__22829));
    LocalMux I__4265 (
            .O(N__22829),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_8 ));
    CascadeMux I__4264 (
            .O(N__22826),
            .I(N__22823));
    InMux I__4263 (
            .O(N__22823),
            .I(N__22820));
    LocalMux I__4262 (
            .O(N__22820),
            .I(\POWERLED.dutycycle_RNIZ0Z_2 ));
    CascadeMux I__4261 (
            .O(N__22817),
            .I(N__22814));
    InMux I__4260 (
            .O(N__22814),
            .I(N__22808));
    InMux I__4259 (
            .O(N__22813),
            .I(N__22801));
    InMux I__4258 (
            .O(N__22812),
            .I(N__22801));
    InMux I__4257 (
            .O(N__22811),
            .I(N__22801));
    LocalMux I__4256 (
            .O(N__22808),
            .I(N__22798));
    LocalMux I__4255 (
            .O(N__22801),
            .I(N__22795));
    Odrv4 I__4254 (
            .O(N__22798),
            .I(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ));
    Odrv12 I__4253 (
            .O(N__22795),
            .I(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ));
    CascadeMux I__4252 (
            .O(N__22790),
            .I(N__22786));
    InMux I__4251 (
            .O(N__22789),
            .I(N__22780));
    InMux I__4250 (
            .O(N__22786),
            .I(N__22780));
    InMux I__4249 (
            .O(N__22785),
            .I(N__22777));
    LocalMux I__4248 (
            .O(N__22780),
            .I(N__22774));
    LocalMux I__4247 (
            .O(N__22777),
            .I(N__22771));
    Span4Mux_v I__4246 (
            .O(N__22774),
            .I(N__22768));
    Odrv4 I__4245 (
            .O(N__22771),
            .I(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ));
    Odrv4 I__4244 (
            .O(N__22768),
            .I(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ));
    CascadeMux I__4243 (
            .O(N__22763),
            .I(N__22760));
    InMux I__4242 (
            .O(N__22760),
            .I(N__22757));
    LocalMux I__4241 (
            .O(N__22757),
            .I(\POWERLED.mult1_un47_sum_axb_4 ));
    InMux I__4240 (
            .O(N__22754),
            .I(N__22751));
    LocalMux I__4239 (
            .O(N__22751),
            .I(N__22748));
    Odrv4 I__4238 (
            .O(N__22748),
            .I(\POWERLED.mult1_un159_sum_i ));
    CascadeMux I__4237 (
            .O(N__22745),
            .I(N__22741));
    CascadeMux I__4236 (
            .O(N__22744),
            .I(N__22738));
    InMux I__4235 (
            .O(N__22741),
            .I(N__22735));
    InMux I__4234 (
            .O(N__22738),
            .I(N__22732));
    LocalMux I__4233 (
            .O(N__22735),
            .I(N__22729));
    LocalMux I__4232 (
            .O(N__22732),
            .I(N__22724));
    Span4Mux_h I__4231 (
            .O(N__22729),
            .I(N__22724));
    Odrv4 I__4230 (
            .O(N__22724),
            .I(\POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434 ));
    CascadeMux I__4229 (
            .O(N__22721),
            .I(N__22718));
    InMux I__4228 (
            .O(N__22718),
            .I(N__22715));
    LocalMux I__4227 (
            .O(N__22715),
            .I(\POWERLED.un1_dutycycle_53_i_29 ));
    InMux I__4226 (
            .O(N__22712),
            .I(\POWERLED.mult1_un47_sum_cry_2 ));
    CascadeMux I__4225 (
            .O(N__22709),
            .I(N__22706));
    InMux I__4224 (
            .O(N__22706),
            .I(N__22703));
    LocalMux I__4223 (
            .O(N__22703),
            .I(\POWERLED.mult1_un47_sum_cry_4_s ));
    InMux I__4222 (
            .O(N__22700),
            .I(\POWERLED.mult1_un47_sum_cry_3 ));
    CascadeMux I__4221 (
            .O(N__22697),
            .I(N__22694));
    InMux I__4220 (
            .O(N__22694),
            .I(N__22691));
    LocalMux I__4219 (
            .O(N__22691),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_4 ));
    CascadeMux I__4218 (
            .O(N__22688),
            .I(N__22685));
    InMux I__4217 (
            .O(N__22685),
            .I(N__22682));
    LocalMux I__4216 (
            .O(N__22682),
            .I(\POWERLED.mult1_un47_sum_cry_5_s ));
    InMux I__4215 (
            .O(N__22679),
            .I(\POWERLED.mult1_un47_sum_cry_4 ));
    CascadeMux I__4214 (
            .O(N__22676),
            .I(N__22673));
    InMux I__4213 (
            .O(N__22673),
            .I(N__22670));
    LocalMux I__4212 (
            .O(N__22670),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_5 ));
    InMux I__4211 (
            .O(N__22667),
            .I(N__22660));
    InMux I__4210 (
            .O(N__22666),
            .I(N__22660));
    InMux I__4209 (
            .O(N__22665),
            .I(N__22657));
    LocalMux I__4208 (
            .O(N__22660),
            .I(\POWERLED.mult1_un47_sum_cry_6_s ));
    LocalMux I__4207 (
            .O(N__22657),
            .I(\POWERLED.mult1_un47_sum_cry_6_s ));
    InMux I__4206 (
            .O(N__22652),
            .I(\POWERLED.mult1_un47_sum_cry_5 ));
    CascadeMux I__4205 (
            .O(N__22649),
            .I(N__22646));
    InMux I__4204 (
            .O(N__22646),
            .I(N__22643));
    LocalMux I__4203 (
            .O(N__22643),
            .I(\POWERLED.mult1_un54_sum_cry_7_THRU_CO ));
    InMux I__4202 (
            .O(N__22640),
            .I(\POWERLED.mult1_un47_sum_cry_6 ));
    CascadeMux I__4201 (
            .O(N__22637),
            .I(N__22633));
    InMux I__4200 (
            .O(N__22636),
            .I(N__22627));
    InMux I__4199 (
            .O(N__22633),
            .I(N__22627));
    InMux I__4198 (
            .O(N__22632),
            .I(N__22624));
    LocalMux I__4197 (
            .O(N__22627),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    LocalMux I__4196 (
            .O(N__22624),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    CascadeMux I__4195 (
            .O(N__22619),
            .I(\POWERLED.mult1_un54_sum_s_8_cascade_ ));
    CascadeMux I__4194 (
            .O(N__22616),
            .I(N__22612));
    CascadeMux I__4193 (
            .O(N__22615),
            .I(N__22608));
    InMux I__4192 (
            .O(N__22612),
            .I(N__22601));
    InMux I__4191 (
            .O(N__22611),
            .I(N__22601));
    InMux I__4190 (
            .O(N__22608),
            .I(N__22601));
    LocalMux I__4189 (
            .O(N__22601),
            .I(\POWERLED.mult1_un54_sum_i_8 ));
    CascadeMux I__4188 (
            .O(N__22598),
            .I(\POWERLED.N_71_cascade_ ));
    CascadeMux I__4187 (
            .O(N__22595),
            .I(\POWERLED.dutycycleZ0Z_0_cascade_ ));
    CascadeMux I__4186 (
            .O(N__22592),
            .I(N__22589));
    InMux I__4185 (
            .O(N__22589),
            .I(N__22586));
    LocalMux I__4184 (
            .O(N__22586),
            .I(N__22583));
    Span4Mux_h I__4183 (
            .O(N__22583),
            .I(N__22580));
    Odrv4 I__4182 (
            .O(N__22580),
            .I(\POWERLED.mult1_un152_sum_i ));
    CascadeMux I__4181 (
            .O(N__22577),
            .I(\POWERLED.N_426_i_cascade_ ));
    InMux I__4180 (
            .O(N__22574),
            .I(N__22571));
    LocalMux I__4179 (
            .O(N__22571),
            .I(\POWERLED.dutycycle_eena_1 ));
    InMux I__4178 (
            .O(N__22568),
            .I(N__22565));
    LocalMux I__4177 (
            .O(N__22565),
            .I(\POWERLED.N_71 ));
    CascadeMux I__4176 (
            .O(N__22562),
            .I(\POWERLED.dutycycle_eena_1_cascade_ ));
    InMux I__4175 (
            .O(N__22559),
            .I(N__22553));
    InMux I__4174 (
            .O(N__22558),
            .I(N__22553));
    LocalMux I__4173 (
            .O(N__22553),
            .I(\POWERLED.dutycycleZ1Z_2 ));
    CascadeMux I__4172 (
            .O(N__22550),
            .I(N__22544));
    InMux I__4171 (
            .O(N__22549),
            .I(N__22540));
    InMux I__4170 (
            .O(N__22548),
            .I(N__22528));
    InMux I__4169 (
            .O(N__22547),
            .I(N__22528));
    InMux I__4168 (
            .O(N__22544),
            .I(N__22528));
    InMux I__4167 (
            .O(N__22543),
            .I(N__22528));
    LocalMux I__4166 (
            .O(N__22540),
            .I(N__22525));
    InMux I__4165 (
            .O(N__22539),
            .I(N__22514));
    InMux I__4164 (
            .O(N__22538),
            .I(N__22514));
    InMux I__4163 (
            .O(N__22537),
            .I(N__22514));
    LocalMux I__4162 (
            .O(N__22528),
            .I(N__22511));
    Span4Mux_v I__4161 (
            .O(N__22525),
            .I(N__22508));
    CascadeMux I__4160 (
            .O(N__22524),
            .I(N__22505));
    InMux I__4159 (
            .O(N__22523),
            .I(N__22500));
    InMux I__4158 (
            .O(N__22522),
            .I(N__22497));
    InMux I__4157 (
            .O(N__22521),
            .I(N__22494));
    LocalMux I__4156 (
            .O(N__22514),
            .I(N__22491));
    Span4Mux_v I__4155 (
            .O(N__22511),
            .I(N__22486));
    Span4Mux_h I__4154 (
            .O(N__22508),
            .I(N__22486));
    InMux I__4153 (
            .O(N__22505),
            .I(N__22481));
    InMux I__4152 (
            .O(N__22504),
            .I(N__22481));
    InMux I__4151 (
            .O(N__22503),
            .I(N__22478));
    LocalMux I__4150 (
            .O(N__22500),
            .I(N__22475));
    LocalMux I__4149 (
            .O(N__22497),
            .I(COUNTER_un4_counter_7_THRU_CO));
    LocalMux I__4148 (
            .O(N__22494),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv12 I__4147 (
            .O(N__22491),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv4 I__4146 (
            .O(N__22486),
            .I(COUNTER_un4_counter_7_THRU_CO));
    LocalMux I__4145 (
            .O(N__22481),
            .I(COUNTER_un4_counter_7_THRU_CO));
    LocalMux I__4144 (
            .O(N__22478),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv12 I__4143 (
            .O(N__22475),
            .I(COUNTER_un4_counter_7_THRU_CO));
    InMux I__4142 (
            .O(N__22460),
            .I(N__22457));
    LocalMux I__4141 (
            .O(N__22457),
            .I(\POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1GZ0 ));
    InMux I__4140 (
            .O(N__22454),
            .I(N__22448));
    InMux I__4139 (
            .O(N__22453),
            .I(N__22448));
    LocalMux I__4138 (
            .O(N__22448),
            .I(\POWERLED.dutycycleZ1Z_7 ));
    CascadeMux I__4137 (
            .O(N__22445),
            .I(\POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1GZ0_cascade_ ));
    InMux I__4136 (
            .O(N__22442),
            .I(N__22439));
    LocalMux I__4135 (
            .O(N__22439),
            .I(\POWERLED.N_540_1 ));
    InMux I__4134 (
            .O(N__22436),
            .I(N__22433));
    LocalMux I__4133 (
            .O(N__22433),
            .I(\POWERLED.N_542 ));
    InMux I__4132 (
            .O(N__22430),
            .I(N__22427));
    LocalMux I__4131 (
            .O(N__22427),
            .I(N__22423));
    InMux I__4130 (
            .O(N__22426),
            .I(N__22420));
    Odrv4 I__4129 (
            .O(N__22423),
            .I(\POWERLED.N_673 ));
    LocalMux I__4128 (
            .O(N__22420),
            .I(\POWERLED.N_673 ));
    CascadeMux I__4127 (
            .O(N__22415),
            .I(\POWERLED.func_state_1_m2s2_i_0_1_cascade_ ));
    InMux I__4126 (
            .O(N__22412),
            .I(N__22409));
    LocalMux I__4125 (
            .O(N__22409),
            .I(\POWERLED.N_6_1 ));
    CascadeMux I__4124 (
            .O(N__22406),
            .I(\POWERLED.N_74_cascade_ ));
    InMux I__4123 (
            .O(N__22403),
            .I(N__22400));
    LocalMux I__4122 (
            .O(N__22400),
            .I(\POWERLED.func_state_1_m2_ns_1_1 ));
    InMux I__4121 (
            .O(N__22397),
            .I(N__22391));
    InMux I__4120 (
            .O(N__22396),
            .I(N__22391));
    LocalMux I__4119 (
            .O(N__22391),
            .I(\POWERLED.func_state_1_m2_1 ));
    InMux I__4118 (
            .O(N__22388),
            .I(N__22384));
    InMux I__4117 (
            .O(N__22387),
            .I(N__22381));
    LocalMux I__4116 (
            .O(N__22384),
            .I(N__22378));
    LocalMux I__4115 (
            .O(N__22381),
            .I(\POWERLED.func_state_RNIBVNSZ0Z_0 ));
    Odrv4 I__4114 (
            .O(N__22378),
            .I(\POWERLED.func_state_RNIBVNSZ0Z_0 ));
    InMux I__4113 (
            .O(N__22373),
            .I(N__22370));
    LocalMux I__4112 (
            .O(N__22370),
            .I(\POWERLED.N_6_2 ));
    InMux I__4111 (
            .O(N__22367),
            .I(N__22364));
    LocalMux I__4110 (
            .O(N__22364),
            .I(\POWERLED.dutycycle_1_0_iv_i_0_a2_0_1_2 ));
    CascadeMux I__4109 (
            .O(N__22361),
            .I(\POWERLED.dutycycle_1_0_iv_i_0_0_2_cascade_ ));
    InMux I__4108 (
            .O(N__22358),
            .I(N__22355));
    LocalMux I__4107 (
            .O(N__22355),
            .I(\POWERLED.un1_func_state25_6_0_0_0_2 ));
    InMux I__4106 (
            .O(N__22352),
            .I(N__22346));
    InMux I__4105 (
            .O(N__22351),
            .I(N__22346));
    LocalMux I__4104 (
            .O(N__22346),
            .I(N__22343));
    Span4Mux_s2_v I__4103 (
            .O(N__22343),
            .I(N__22340));
    Span4Mux_v I__4102 (
            .O(N__22340),
            .I(N__22337));
    Odrv4 I__4101 (
            .O(N__22337),
            .I(\POWERLED.func_state_RNI5SKJ1Z0Z_1 ));
    CascadeMux I__4100 (
            .O(N__22334),
            .I(N__22327));
    CascadeMux I__4099 (
            .O(N__22333),
            .I(N__22324));
    InMux I__4098 (
            .O(N__22332),
            .I(N__22319));
    InMux I__4097 (
            .O(N__22331),
            .I(N__22312));
    InMux I__4096 (
            .O(N__22330),
            .I(N__22312));
    InMux I__4095 (
            .O(N__22327),
            .I(N__22312));
    InMux I__4094 (
            .O(N__22324),
            .I(N__22305));
    InMux I__4093 (
            .O(N__22323),
            .I(N__22305));
    InMux I__4092 (
            .O(N__22322),
            .I(N__22305));
    LocalMux I__4091 (
            .O(N__22319),
            .I(N__22302));
    LocalMux I__4090 (
            .O(N__22312),
            .I(N__22297));
    LocalMux I__4089 (
            .O(N__22305),
            .I(N__22297));
    Span4Mux_v I__4088 (
            .O(N__22302),
            .I(N__22294));
    Span12Mux_v I__4087 (
            .O(N__22297),
            .I(N__22291));
    Span4Mux_v I__4086 (
            .O(N__22294),
            .I(N__22288));
    Odrv12 I__4085 (
            .O(N__22291),
            .I(vddq_ok));
    Odrv4 I__4084 (
            .O(N__22288),
            .I(vddq_ok));
    CascadeMux I__4083 (
            .O(N__22283),
            .I(func_state_RNI_2_0_cascade_));
    InMux I__4082 (
            .O(N__22280),
            .I(N__22277));
    LocalMux I__4081 (
            .O(N__22277),
            .I(\POWERLED.func_state_1_m0_1_1 ));
    CascadeMux I__4080 (
            .O(N__22274),
            .I(v5s_enn_cascade_));
    InMux I__4079 (
            .O(N__22271),
            .I(N__22268));
    LocalMux I__4078 (
            .O(N__22268),
            .I(\POWERLED.func_state_en_0_0 ));
    InMux I__4077 (
            .O(N__22265),
            .I(N__22259));
    InMux I__4076 (
            .O(N__22264),
            .I(N__22259));
    LocalMux I__4075 (
            .O(N__22259),
            .I(\POWERLED.func_stateZ1Z_0 ));
    CascadeMux I__4074 (
            .O(N__22256),
            .I(\POWERLED.func_state_en_0_0_cascade_ ));
    CascadeMux I__4073 (
            .O(N__22253),
            .I(N__22248));
    CascadeMux I__4072 (
            .O(N__22252),
            .I(N__22245));
    CascadeMux I__4071 (
            .O(N__22251),
            .I(N__22242));
    InMux I__4070 (
            .O(N__22248),
            .I(N__22237));
    InMux I__4069 (
            .O(N__22245),
            .I(N__22237));
    InMux I__4068 (
            .O(N__22242),
            .I(N__22234));
    LocalMux I__4067 (
            .O(N__22237),
            .I(RSMRSTn_fast));
    LocalMux I__4066 (
            .O(N__22234),
            .I(RSMRSTn_fast));
    CascadeMux I__4065 (
            .O(N__22229),
            .I(N__22226));
    InMux I__4064 (
            .O(N__22226),
            .I(N__22223));
    LocalMux I__4063 (
            .O(N__22223),
            .I(N__22220));
    Span4Mux_h I__4062 (
            .O(N__22220),
            .I(N__22217));
    Odrv4 I__4061 (
            .O(N__22217),
            .I(\COUNTER.un4_counter_3_and ));
    CascadeMux I__4060 (
            .O(N__22214),
            .I(N__22211));
    InMux I__4059 (
            .O(N__22211),
            .I(N__22208));
    LocalMux I__4058 (
            .O(N__22208),
            .I(\COUNTER.un4_counter_4_and ));
    CascadeMux I__4057 (
            .O(N__22205),
            .I(N__22202));
    InMux I__4056 (
            .O(N__22202),
            .I(N__22199));
    LocalMux I__4055 (
            .O(N__22199),
            .I(\COUNTER.un4_counter_5_and ));
    CascadeMux I__4054 (
            .O(N__22196),
            .I(N__22193));
    InMux I__4053 (
            .O(N__22193),
            .I(N__22190));
    LocalMux I__4052 (
            .O(N__22190),
            .I(N__22187));
    Span4Mux_h I__4051 (
            .O(N__22187),
            .I(N__22184));
    Odrv4 I__4050 (
            .O(N__22184),
            .I(\COUNTER.un4_counter_6_and ));
    CascadeMux I__4049 (
            .O(N__22181),
            .I(N__22178));
    InMux I__4048 (
            .O(N__22178),
            .I(N__22175));
    LocalMux I__4047 (
            .O(N__22175),
            .I(N__22172));
    Span4Mux_h I__4046 (
            .O(N__22172),
            .I(N__22169));
    Odrv4 I__4045 (
            .O(N__22169),
            .I(\COUNTER.un4_counter_7_and ));
    InMux I__4044 (
            .O(N__22166),
            .I(bfn_8_5_0_));
    CascadeMux I__4043 (
            .O(N__22163),
            .I(\POWERLED.N_673_0_cascade_ ));
    InMux I__4042 (
            .O(N__22160),
            .I(N__22157));
    LocalMux I__4041 (
            .O(N__22157),
            .I(\POWERLED.N_423_0 ));
    InMux I__4040 (
            .O(N__22154),
            .I(N__22148));
    InMux I__4039 (
            .O(N__22153),
            .I(N__22148));
    LocalMux I__4038 (
            .O(N__22148),
            .I(\POWERLED.count_off_1_14 ));
    InMux I__4037 (
            .O(N__22145),
            .I(N__22142));
    LocalMux I__4036 (
            .O(N__22142),
            .I(\POWERLED.count_off_0_14 ));
    InMux I__4035 (
            .O(N__22139),
            .I(N__22133));
    InMux I__4034 (
            .O(N__22138),
            .I(N__22133));
    LocalMux I__4033 (
            .O(N__22133),
            .I(\POWERLED.un3_count_off_1_cry_14_c_RNIPGZ0Z497 ));
    InMux I__4032 (
            .O(N__22130),
            .I(N__22127));
    LocalMux I__4031 (
            .O(N__22127),
            .I(\POWERLED.count_off_0_15 ));
    InMux I__4030 (
            .O(N__22124),
            .I(N__22121));
    LocalMux I__4029 (
            .O(N__22121),
            .I(\POWERLED.count_offZ0Z_15 ));
    InMux I__4028 (
            .O(N__22118),
            .I(N__22114));
    InMux I__4027 (
            .O(N__22117),
            .I(N__22111));
    LocalMux I__4026 (
            .O(N__22114),
            .I(\POWERLED.count_offZ0Z_13 ));
    LocalMux I__4025 (
            .O(N__22111),
            .I(\POWERLED.count_offZ0Z_13 ));
    InMux I__4024 (
            .O(N__22106),
            .I(N__22102));
    InMux I__4023 (
            .O(N__22105),
            .I(N__22099));
    LocalMux I__4022 (
            .O(N__22102),
            .I(\POWERLED.count_offZ0Z_14 ));
    LocalMux I__4021 (
            .O(N__22099),
            .I(\POWERLED.count_offZ0Z_14 ));
    CascadeMux I__4020 (
            .O(N__22094),
            .I(\POWERLED.count_offZ0Z_15_cascade_ ));
    CascadeMux I__4019 (
            .O(N__22091),
            .I(N__22086));
    CascadeMux I__4018 (
            .O(N__22090),
            .I(N__22082));
    InMux I__4017 (
            .O(N__22089),
            .I(N__22079));
    InMux I__4016 (
            .O(N__22086),
            .I(N__22074));
    InMux I__4015 (
            .O(N__22085),
            .I(N__22074));
    InMux I__4014 (
            .O(N__22082),
            .I(N__22071));
    LocalMux I__4013 (
            .O(N__22079),
            .I(\POWERLED.count_offZ0Z_0 ));
    LocalMux I__4012 (
            .O(N__22074),
            .I(\POWERLED.count_offZ0Z_0 ));
    LocalMux I__4011 (
            .O(N__22071),
            .I(\POWERLED.count_offZ0Z_0 ));
    InMux I__4010 (
            .O(N__22064),
            .I(N__22061));
    LocalMux I__4009 (
            .O(N__22061),
            .I(N__22058));
    Span4Mux_h I__4008 (
            .O(N__22058),
            .I(N__22055));
    Odrv4 I__4007 (
            .O(N__22055),
            .I(\POWERLED.count_off_0_6 ));
    InMux I__4006 (
            .O(N__22052),
            .I(N__22049));
    LocalMux I__4005 (
            .O(N__22049),
            .I(N__22045));
    InMux I__4004 (
            .O(N__22048),
            .I(N__22042));
    Odrv4 I__4003 (
            .O(N__22045),
            .I(\POWERLED.count_off_1_6 ));
    LocalMux I__4002 (
            .O(N__22042),
            .I(\POWERLED.count_off_1_6 ));
    InMux I__4001 (
            .O(N__22037),
            .I(N__22033));
    InMux I__4000 (
            .O(N__22036),
            .I(N__22030));
    LocalMux I__3999 (
            .O(N__22033),
            .I(\POWERLED.count_offZ0Z_6 ));
    LocalMux I__3998 (
            .O(N__22030),
            .I(\POWERLED.count_offZ0Z_6 ));
    CascadeMux I__3997 (
            .O(N__22025),
            .I(N__22022));
    InMux I__3996 (
            .O(N__22022),
            .I(N__22019));
    LocalMux I__3995 (
            .O(N__22019),
            .I(N__22016));
    Odrv4 I__3994 (
            .O(N__22016),
            .I(\COUNTER.un4_counter_0_and ));
    CascadeMux I__3993 (
            .O(N__22013),
            .I(N__22010));
    InMux I__3992 (
            .O(N__22010),
            .I(N__22007));
    LocalMux I__3991 (
            .O(N__22007),
            .I(N__22004));
    Odrv12 I__3990 (
            .O(N__22004),
            .I(\COUNTER.un4_counter_1_and ));
    CascadeMux I__3989 (
            .O(N__22001),
            .I(N__21998));
    InMux I__3988 (
            .O(N__21998),
            .I(N__21995));
    LocalMux I__3987 (
            .O(N__21995),
            .I(N__21992));
    Odrv4 I__3986 (
            .O(N__21992),
            .I(\COUNTER.un4_counter_2_and ));
    InMux I__3985 (
            .O(N__21989),
            .I(N__21986));
    LocalMux I__3984 (
            .O(N__21986),
            .I(N__21983));
    Span4Mux_h I__3983 (
            .O(N__21983),
            .I(N__21980));
    Odrv4 I__3982 (
            .O(N__21980),
            .I(\POWERLED.count_off_0_5 ));
    InMux I__3981 (
            .O(N__21977),
            .I(N__21974));
    LocalMux I__3980 (
            .O(N__21974),
            .I(N__21971));
    Span4Mux_s0_v I__3979 (
            .O(N__21971),
            .I(N__21967));
    InMux I__3978 (
            .O(N__21970),
            .I(N__21964));
    Odrv4 I__3977 (
            .O(N__21967),
            .I(\POWERLED.count_off_1_5 ));
    LocalMux I__3976 (
            .O(N__21964),
            .I(\POWERLED.count_off_1_5 ));
    InMux I__3975 (
            .O(N__21959),
            .I(N__21956));
    LocalMux I__3974 (
            .O(N__21956),
            .I(\POWERLED.count_offZ0Z_5 ));
    CascadeMux I__3973 (
            .O(N__21953),
            .I(\POWERLED.count_offZ0Z_5_cascade_ ));
    InMux I__3972 (
            .O(N__21950),
            .I(N__21947));
    LocalMux I__3971 (
            .O(N__21947),
            .I(\POWERLED.count_off_0_0 ));
    InMux I__3970 (
            .O(N__21944),
            .I(N__21941));
    LocalMux I__3969 (
            .O(N__21941),
            .I(\POWERLED.count_off_1_0 ));
    InMux I__3968 (
            .O(N__21938),
            .I(N__21935));
    LocalMux I__3967 (
            .O(N__21935),
            .I(\POWERLED.count_off_0_2 ));
    CascadeMux I__3966 (
            .O(N__21932),
            .I(N__21929));
    InMux I__3965 (
            .O(N__21929),
            .I(N__21923));
    InMux I__3964 (
            .O(N__21928),
            .I(N__21923));
    LocalMux I__3963 (
            .O(N__21923),
            .I(\POWERLED.count_off_1_2 ));
    InMux I__3962 (
            .O(N__21920),
            .I(N__21916));
    InMux I__3961 (
            .O(N__21919),
            .I(N__21913));
    LocalMux I__3960 (
            .O(N__21916),
            .I(\POWERLED.count_offZ0Z_2 ));
    LocalMux I__3959 (
            .O(N__21913),
            .I(\POWERLED.count_offZ0Z_2 ));
    InMux I__3958 (
            .O(N__21908),
            .I(N__21902));
    InMux I__3957 (
            .O(N__21907),
            .I(N__21902));
    LocalMux I__3956 (
            .O(N__21902),
            .I(\POWERLED.count_off_1_13 ));
    InMux I__3955 (
            .O(N__21899),
            .I(N__21896));
    LocalMux I__3954 (
            .O(N__21896),
            .I(\POWERLED.count_off_0_13 ));
    CascadeMux I__3953 (
            .O(N__21893),
            .I(\POWERLED.N_598_cascade_ ));
    CascadeMux I__3952 (
            .O(N__21890),
            .I(\POWERLED.N_450_cascade_ ));
    InMux I__3951 (
            .O(N__21887),
            .I(N__21884));
    LocalMux I__3950 (
            .O(N__21884),
            .I(\POWERLED.N_599 ));
    CascadeMux I__3949 (
            .O(N__21881),
            .I(\POWERLED.N_449_cascade_ ));
    InMux I__3948 (
            .O(N__21878),
            .I(N__21875));
    LocalMux I__3947 (
            .O(N__21875),
            .I(\POWERLED.N_2376_i ));
    CascadeMux I__3946 (
            .O(N__21872),
            .I(\POWERLED.N_2376_i_cascade_ ));
    CascadeMux I__3945 (
            .O(N__21869),
            .I(\POWERLED.count_offZ0Z_0_cascade_ ));
    InMux I__3944 (
            .O(N__21866),
            .I(\POWERLED.un1_dutycycle_53_cry_14 ));
    InMux I__3943 (
            .O(N__21863),
            .I(bfn_7_15_0_));
    InMux I__3942 (
            .O(N__21860),
            .I(\POWERLED.CO2 ));
    CascadeMux I__3941 (
            .O(N__21857),
            .I(N__21854));
    InMux I__3940 (
            .O(N__21854),
            .I(N__21848));
    InMux I__3939 (
            .O(N__21853),
            .I(N__21848));
    LocalMux I__3938 (
            .O(N__21848),
            .I(N__21845));
    Span4Mux_v I__3937 (
            .O(N__21845),
            .I(N__21842));
    Odrv4 I__3936 (
            .O(N__21842),
            .I(\POWERLED.CO2_THRU_CO ));
    CascadeMux I__3935 (
            .O(N__21839),
            .I(N__21836));
    InMux I__3934 (
            .O(N__21836),
            .I(N__21833));
    LocalMux I__3933 (
            .O(N__21833),
            .I(\POWERLED.dutycycle_RNIZ0Z_14 ));
    InMux I__3932 (
            .O(N__21830),
            .I(N__21826));
    InMux I__3931 (
            .O(N__21829),
            .I(N__21823));
    LocalMux I__3930 (
            .O(N__21826),
            .I(\POWERLED.mult1_un68_sum ));
    LocalMux I__3929 (
            .O(N__21823),
            .I(\POWERLED.mult1_un68_sum ));
    InMux I__3928 (
            .O(N__21818),
            .I(N__21815));
    LocalMux I__3927 (
            .O(N__21815),
            .I(\POWERLED.mult1_un68_sum_i ));
    InMux I__3926 (
            .O(N__21812),
            .I(N__21809));
    LocalMux I__3925 (
            .O(N__21809),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_15 ));
    CascadeMux I__3924 (
            .O(N__21806),
            .I(N__21803));
    InMux I__3923 (
            .O(N__21803),
            .I(N__21799));
    InMux I__3922 (
            .O(N__21802),
            .I(N__21796));
    LocalMux I__3921 (
            .O(N__21799),
            .I(N__21793));
    LocalMux I__3920 (
            .O(N__21796),
            .I(\POWERLED.mult1_un82_sum ));
    Odrv4 I__3919 (
            .O(N__21793),
            .I(\POWERLED.mult1_un82_sum ));
    InMux I__3918 (
            .O(N__21788),
            .I(N__21785));
    LocalMux I__3917 (
            .O(N__21785),
            .I(N__21782));
    Odrv4 I__3916 (
            .O(N__21782),
            .I(\POWERLED.mult1_un82_sum_i ));
    InMux I__3915 (
            .O(N__21779),
            .I(N__21775));
    InMux I__3914 (
            .O(N__21778),
            .I(N__21772));
    LocalMux I__3913 (
            .O(N__21775),
            .I(N__21769));
    LocalMux I__3912 (
            .O(N__21772),
            .I(\POWERLED.mult1_un61_sum ));
    Odrv4 I__3911 (
            .O(N__21769),
            .I(\POWERLED.mult1_un61_sum ));
    InMux I__3910 (
            .O(N__21764),
            .I(N__21761));
    LocalMux I__3909 (
            .O(N__21761),
            .I(\POWERLED.mult1_un61_sum_i ));
    InMux I__3908 (
            .O(N__21758),
            .I(N__21754));
    InMux I__3907 (
            .O(N__21757),
            .I(N__21751));
    LocalMux I__3906 (
            .O(N__21754),
            .I(N__21748));
    LocalMux I__3905 (
            .O(N__21751),
            .I(\POWERLED.mult1_un103_sum ));
    Odrv4 I__3904 (
            .O(N__21748),
            .I(\POWERLED.mult1_un103_sum ));
    InMux I__3903 (
            .O(N__21743),
            .I(\POWERLED.un1_dutycycle_53_cry_5 ));
    InMux I__3902 (
            .O(N__21740),
            .I(N__21736));
    InMux I__3901 (
            .O(N__21739),
            .I(N__21733));
    LocalMux I__3900 (
            .O(N__21736),
            .I(N__21730));
    LocalMux I__3899 (
            .O(N__21733),
            .I(N__21727));
    Span4Mux_h I__3898 (
            .O(N__21730),
            .I(N__21724));
    Odrv12 I__3897 (
            .O(N__21727),
            .I(\POWERLED.mult1_un96_sum ));
    Odrv4 I__3896 (
            .O(N__21724),
            .I(\POWERLED.mult1_un96_sum ));
    InMux I__3895 (
            .O(N__21719),
            .I(\POWERLED.un1_dutycycle_53_cry_6 ));
    InMux I__3894 (
            .O(N__21716),
            .I(N__21712));
    InMux I__3893 (
            .O(N__21715),
            .I(N__21709));
    LocalMux I__3892 (
            .O(N__21712),
            .I(N__21704));
    LocalMux I__3891 (
            .O(N__21709),
            .I(N__21704));
    Span4Mux_s2_v I__3890 (
            .O(N__21704),
            .I(N__21701));
    Odrv4 I__3889 (
            .O(N__21701),
            .I(\POWERLED.mult1_un89_sum ));
    InMux I__3888 (
            .O(N__21698),
            .I(bfn_7_14_0_));
    InMux I__3887 (
            .O(N__21695),
            .I(\POWERLED.un1_dutycycle_53_cry_8 ));
    InMux I__3886 (
            .O(N__21692),
            .I(N__21689));
    LocalMux I__3885 (
            .O(N__21689),
            .I(N__21685));
    InMux I__3884 (
            .O(N__21688),
            .I(N__21682));
    Odrv4 I__3883 (
            .O(N__21685),
            .I(\POWERLED.mult1_un75_sum ));
    LocalMux I__3882 (
            .O(N__21682),
            .I(\POWERLED.mult1_un75_sum ));
    InMux I__3881 (
            .O(N__21677),
            .I(\POWERLED.un1_dutycycle_53_cry_9 ));
    InMux I__3880 (
            .O(N__21674),
            .I(\POWERLED.un1_dutycycle_53_cry_10 ));
    InMux I__3879 (
            .O(N__21671),
            .I(\POWERLED.un1_dutycycle_53_cry_11 ));
    InMux I__3878 (
            .O(N__21668),
            .I(N__21665));
    LocalMux I__3877 (
            .O(N__21665),
            .I(N__21662));
    Span4Mux_v I__3876 (
            .O(N__21662),
            .I(N__21659));
    Span4Mux_v I__3875 (
            .O(N__21659),
            .I(N__21655));
    InMux I__3874 (
            .O(N__21658),
            .I(N__21652));
    Span4Mux_h I__3873 (
            .O(N__21655),
            .I(N__21647));
    LocalMux I__3872 (
            .O(N__21652),
            .I(N__21647));
    Odrv4 I__3871 (
            .O(N__21647),
            .I(\POWERLED.mult1_un54_sum ));
    InMux I__3870 (
            .O(N__21644),
            .I(\POWERLED.un1_dutycycle_53_cry_12 ));
    InMux I__3869 (
            .O(N__21641),
            .I(\POWERLED.un1_dutycycle_53_cry_13 ));
    CascadeMux I__3868 (
            .O(N__21638),
            .I(N__21635));
    InMux I__3867 (
            .O(N__21635),
            .I(N__21632));
    LocalMux I__3866 (
            .O(N__21632),
            .I(\POWERLED.mult1_un61_sum_axb_8 ));
    InMux I__3865 (
            .O(N__21629),
            .I(\POWERLED.mult1_un61_sum_cry_7 ));
    CascadeMux I__3864 (
            .O(N__21626),
            .I(N__21622));
    InMux I__3863 (
            .O(N__21625),
            .I(N__21617));
    InMux I__3862 (
            .O(N__21622),
            .I(N__21617));
    LocalMux I__3861 (
            .O(N__21617),
            .I(N__21611));
    InMux I__3860 (
            .O(N__21616),
            .I(N__21608));
    InMux I__3859 (
            .O(N__21615),
            .I(N__21603));
    InMux I__3858 (
            .O(N__21614),
            .I(N__21603));
    Odrv4 I__3857 (
            .O(N__21611),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__3856 (
            .O(N__21608),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__3855 (
            .O(N__21603),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    CascadeMux I__3854 (
            .O(N__21596),
            .I(N__21593));
    InMux I__3853 (
            .O(N__21593),
            .I(N__21590));
    LocalMux I__3852 (
            .O(N__21590),
            .I(\POWERLED.un1_dutycycle_53_i_28 ));
    InMux I__3851 (
            .O(N__21587),
            .I(N__21584));
    LocalMux I__3850 (
            .O(N__21584),
            .I(N__21581));
    Span4Mux_v I__3849 (
            .O(N__21581),
            .I(N__21577));
    InMux I__3848 (
            .O(N__21580),
            .I(N__21574));
    Odrv4 I__3847 (
            .O(N__21577),
            .I(\POWERLED.un1_dutycycle_53_axb_0 ));
    LocalMux I__3846 (
            .O(N__21574),
            .I(\POWERLED.un1_dutycycle_53_axb_0 ));
    InMux I__3845 (
            .O(N__21569),
            .I(N__21566));
    LocalMux I__3844 (
            .O(N__21566),
            .I(N__21562));
    InMux I__3843 (
            .O(N__21565),
            .I(N__21559));
    Odrv4 I__3842 (
            .O(N__21562),
            .I(\POWERLED.mult1_un138_sum ));
    LocalMux I__3841 (
            .O(N__21559),
            .I(\POWERLED.mult1_un138_sum ));
    InMux I__3840 (
            .O(N__21554),
            .I(\POWERLED.un1_dutycycle_53_cry_0 ));
    InMux I__3839 (
            .O(N__21551),
            .I(N__21548));
    LocalMux I__3838 (
            .O(N__21548),
            .I(N__21545));
    Span4Mux_v I__3837 (
            .O(N__21545),
            .I(N__21541));
    InMux I__3836 (
            .O(N__21544),
            .I(N__21538));
    Odrv4 I__3835 (
            .O(N__21541),
            .I(\POWERLED.mult1_un131_sum ));
    LocalMux I__3834 (
            .O(N__21538),
            .I(\POWERLED.mult1_un131_sum ));
    InMux I__3833 (
            .O(N__21533),
            .I(\POWERLED.un1_dutycycle_53_cry_1 ));
    InMux I__3832 (
            .O(N__21530),
            .I(N__21527));
    LocalMux I__3831 (
            .O(N__21527),
            .I(N__21524));
    Span4Mux_v I__3830 (
            .O(N__21524),
            .I(N__21520));
    InMux I__3829 (
            .O(N__21523),
            .I(N__21517));
    Odrv4 I__3828 (
            .O(N__21520),
            .I(\POWERLED.mult1_un124_sum ));
    LocalMux I__3827 (
            .O(N__21517),
            .I(\POWERLED.mult1_un124_sum ));
    InMux I__3826 (
            .O(N__21512),
            .I(\POWERLED.un1_dutycycle_53_cry_2 ));
    InMux I__3825 (
            .O(N__21509),
            .I(N__21506));
    LocalMux I__3824 (
            .O(N__21506),
            .I(N__21503));
    Span4Mux_v I__3823 (
            .O(N__21503),
            .I(N__21499));
    InMux I__3822 (
            .O(N__21502),
            .I(N__21496));
    Span4Mux_v I__3821 (
            .O(N__21499),
            .I(N__21491));
    LocalMux I__3820 (
            .O(N__21496),
            .I(N__21491));
    Span4Mux_v I__3819 (
            .O(N__21491),
            .I(N__21488));
    Odrv4 I__3818 (
            .O(N__21488),
            .I(\POWERLED.mult1_un117_sum ));
    InMux I__3817 (
            .O(N__21485),
            .I(\POWERLED.un1_dutycycle_53_cry_3 ));
    InMux I__3816 (
            .O(N__21482),
            .I(N__21479));
    LocalMux I__3815 (
            .O(N__21479),
            .I(N__21475));
    InMux I__3814 (
            .O(N__21478),
            .I(N__21472));
    Span4Mux_h I__3813 (
            .O(N__21475),
            .I(N__21469));
    LocalMux I__3812 (
            .O(N__21472),
            .I(\POWERLED.mult1_un110_sum ));
    Odrv4 I__3811 (
            .O(N__21469),
            .I(\POWERLED.mult1_un110_sum ));
    InMux I__3810 (
            .O(N__21464),
            .I(\POWERLED.un1_dutycycle_53_cry_4 ));
    InMux I__3809 (
            .O(N__21461),
            .I(\POWERLED.mult1_un54_sum_cry_6 ));
    InMux I__3808 (
            .O(N__21458),
            .I(\POWERLED.mult1_un54_sum_cry_7 ));
    CascadeMux I__3807 (
            .O(N__21455),
            .I(N__21452));
    InMux I__3806 (
            .O(N__21452),
            .I(N__21449));
    LocalMux I__3805 (
            .O(N__21449),
            .I(\POWERLED.mult1_un47_sum_l_fx_6 ));
    InMux I__3804 (
            .O(N__21446),
            .I(N__21443));
    LocalMux I__3803 (
            .O(N__21443),
            .I(N__21440));
    Span4Mux_v I__3802 (
            .O(N__21440),
            .I(N__21437));
    Span4Mux_v I__3801 (
            .O(N__21437),
            .I(N__21434));
    Odrv4 I__3800 (
            .O(N__21434),
            .I(\POWERLED.mult1_un54_sum_i ));
    CascadeMux I__3799 (
            .O(N__21431),
            .I(N__21428));
    InMux I__3798 (
            .O(N__21428),
            .I(N__21425));
    LocalMux I__3797 (
            .O(N__21425),
            .I(N__21422));
    Odrv4 I__3796 (
            .O(N__21422),
            .I(\POWERLED.mult1_un61_sum_cry_3_s ));
    InMux I__3795 (
            .O(N__21419),
            .I(\POWERLED.mult1_un61_sum_cry_2 ));
    CascadeMux I__3794 (
            .O(N__21416),
            .I(N__21413));
    InMux I__3793 (
            .O(N__21413),
            .I(N__21410));
    LocalMux I__3792 (
            .O(N__21410),
            .I(\POWERLED.mult1_un54_sum_cry_3_s ));
    InMux I__3791 (
            .O(N__21407),
            .I(N__21404));
    LocalMux I__3790 (
            .O(N__21404),
            .I(N__21401));
    Odrv4 I__3789 (
            .O(N__21401),
            .I(\POWERLED.mult1_un61_sum_cry_4_s ));
    InMux I__3788 (
            .O(N__21398),
            .I(\POWERLED.mult1_un61_sum_cry_3 ));
    InMux I__3787 (
            .O(N__21395),
            .I(N__21392));
    LocalMux I__3786 (
            .O(N__21392),
            .I(\POWERLED.mult1_un54_sum_cry_4_s ));
    CascadeMux I__3785 (
            .O(N__21389),
            .I(N__21386));
    InMux I__3784 (
            .O(N__21386),
            .I(N__21383));
    LocalMux I__3783 (
            .O(N__21383),
            .I(N__21380));
    Odrv4 I__3782 (
            .O(N__21380),
            .I(\POWERLED.mult1_un61_sum_cry_5_s ));
    InMux I__3781 (
            .O(N__21377),
            .I(\POWERLED.mult1_un61_sum_cry_4 ));
    CascadeMux I__3780 (
            .O(N__21374),
            .I(N__21371));
    InMux I__3779 (
            .O(N__21371),
            .I(N__21368));
    LocalMux I__3778 (
            .O(N__21368),
            .I(\POWERLED.mult1_un54_sum_cry_5_s ));
    InMux I__3777 (
            .O(N__21365),
            .I(N__21362));
    LocalMux I__3776 (
            .O(N__21362),
            .I(N__21359));
    Span4Mux_h I__3775 (
            .O(N__21359),
            .I(N__21356));
    Odrv4 I__3774 (
            .O(N__21356),
            .I(\POWERLED.mult1_un61_sum_cry_6_s ));
    InMux I__3773 (
            .O(N__21353),
            .I(\POWERLED.mult1_un61_sum_cry_5 ));
    InMux I__3772 (
            .O(N__21350),
            .I(N__21347));
    LocalMux I__3771 (
            .O(N__21347),
            .I(\POWERLED.mult1_un54_sum_cry_6_s ));
    InMux I__3770 (
            .O(N__21344),
            .I(N__21341));
    LocalMux I__3769 (
            .O(N__21341),
            .I(N__21338));
    Odrv4 I__3768 (
            .O(N__21338),
            .I(\POWERLED.mult1_un68_sum_axb_8 ));
    InMux I__3767 (
            .O(N__21335),
            .I(\POWERLED.mult1_un61_sum_cry_6 ));
    InMux I__3766 (
            .O(N__21332),
            .I(N__21326));
    InMux I__3765 (
            .O(N__21331),
            .I(N__21326));
    LocalMux I__3764 (
            .O(N__21326),
            .I(N__21323));
    Odrv12 I__3763 (
            .O(N__21323),
            .I(\POWERLED.count_off_1_8 ));
    InMux I__3762 (
            .O(N__21320),
            .I(N__21317));
    LocalMux I__3761 (
            .O(N__21317),
            .I(\POWERLED.count_off_0_8 ));
    InMux I__3760 (
            .O(N__21314),
            .I(\POWERLED.mult1_un54_sum_cry_2 ));
    InMux I__3759 (
            .O(N__21311),
            .I(\POWERLED.mult1_un54_sum_cry_3 ));
    InMux I__3758 (
            .O(N__21308),
            .I(\POWERLED.mult1_un54_sum_cry_4 ));
    InMux I__3757 (
            .O(N__21305),
            .I(\POWERLED.mult1_un54_sum_cry_5 ));
    CascadeMux I__3756 (
            .O(N__21302),
            .I(\POWERLED.N_512_cascade_ ));
    CascadeMux I__3755 (
            .O(N__21299),
            .I(\POWERLED.un1_clk_100khz_39_and_i_1_cascade_ ));
    InMux I__3754 (
            .O(N__21296),
            .I(N__21293));
    LocalMux I__3753 (
            .O(N__21293),
            .I(\POWERLED.N_514 ));
    InMux I__3752 (
            .O(N__21290),
            .I(N__21287));
    LocalMux I__3751 (
            .O(N__21287),
            .I(\POWERLED.N_508 ));
    CascadeMux I__3750 (
            .O(N__21284),
            .I(\POWERLED.un1_clk_100khz_33_and_i_1_cascade_ ));
    InMux I__3749 (
            .O(N__21281),
            .I(N__21275));
    InMux I__3748 (
            .O(N__21280),
            .I(N__21275));
    LocalMux I__3747 (
            .O(N__21275),
            .I(N__21272));
    Span4Mux_v I__3746 (
            .O(N__21272),
            .I(N__21269));
    Odrv4 I__3745 (
            .O(N__21269),
            .I(\POWERLED.count_off_1_7 ));
    InMux I__3744 (
            .O(N__21266),
            .I(N__21263));
    LocalMux I__3743 (
            .O(N__21263),
            .I(\POWERLED.count_off_0_7 ));
    CascadeMux I__3742 (
            .O(N__21260),
            .I(\POWERLED.func_state_1_ss0_i_0_0_1_1_cascade_ ));
    InMux I__3741 (
            .O(N__21257),
            .I(N__21254));
    LocalMux I__3740 (
            .O(N__21254),
            .I(\POWERLED.N_423 ));
    InMux I__3739 (
            .O(N__21251),
            .I(N__21248));
    LocalMux I__3738 (
            .O(N__21248),
            .I(\POWERLED.N_671 ));
    CascadeMux I__3737 (
            .O(N__21245),
            .I(N__21242));
    InMux I__3736 (
            .O(N__21242),
            .I(N__21236));
    InMux I__3735 (
            .O(N__21241),
            .I(N__21236));
    LocalMux I__3734 (
            .O(N__21236),
            .I(N__21233));
    Odrv12 I__3733 (
            .O(N__21233),
            .I(\POWERLED.func_state_enZ0 ));
    CascadeMux I__3732 (
            .O(N__21230),
            .I(N__21226));
    InMux I__3731 (
            .O(N__21229),
            .I(N__21221));
    InMux I__3730 (
            .O(N__21226),
            .I(N__21221));
    LocalMux I__3729 (
            .O(N__21221),
            .I(\POWERLED.func_stateZ0Z_1 ));
    InMux I__3728 (
            .O(N__21218),
            .I(N__21208));
    InMux I__3727 (
            .O(N__21217),
            .I(N__21208));
    InMux I__3726 (
            .O(N__21216),
            .I(N__21199));
    InMux I__3725 (
            .O(N__21215),
            .I(N__21199));
    InMux I__3724 (
            .O(N__21214),
            .I(N__21199));
    InMux I__3723 (
            .O(N__21213),
            .I(N__21199));
    LocalMux I__3722 (
            .O(N__21208),
            .I(N__21190));
    LocalMux I__3721 (
            .O(N__21199),
            .I(N__21190));
    InMux I__3720 (
            .O(N__21198),
            .I(N__21183));
    InMux I__3719 (
            .O(N__21197),
            .I(N__21183));
    InMux I__3718 (
            .O(N__21196),
            .I(N__21183));
    InMux I__3717 (
            .O(N__21195),
            .I(N__21180));
    Odrv4 I__3716 (
            .O(N__21190),
            .I(RSMRST_PWRGD_curr_state_0));
    LocalMux I__3715 (
            .O(N__21183),
            .I(RSMRST_PWRGD_curr_state_0));
    LocalMux I__3714 (
            .O(N__21180),
            .I(RSMRST_PWRGD_curr_state_0));
    InMux I__3713 (
            .O(N__21173),
            .I(N__21170));
    LocalMux I__3712 (
            .O(N__21170),
            .I(N__21164));
    InMux I__3711 (
            .O(N__21169),
            .I(N__21161));
    InMux I__3710 (
            .O(N__21168),
            .I(N__21156));
    InMux I__3709 (
            .O(N__21167),
            .I(N__21156));
    Span4Mux_s1_v I__3708 (
            .O(N__21164),
            .I(N__21153));
    LocalMux I__3707 (
            .O(N__21161),
            .I(N__21145));
    LocalMux I__3706 (
            .O(N__21156),
            .I(N__21140));
    Span4Mux_v I__3705 (
            .O(N__21153),
            .I(N__21140));
    InMux I__3704 (
            .O(N__21152),
            .I(N__21129));
    InMux I__3703 (
            .O(N__21151),
            .I(N__21129));
    InMux I__3702 (
            .O(N__21150),
            .I(N__21129));
    InMux I__3701 (
            .O(N__21149),
            .I(N__21129));
    InMux I__3700 (
            .O(N__21148),
            .I(N__21129));
    Span4Mux_h I__3699 (
            .O(N__21145),
            .I(N__21124));
    Span4Mux_h I__3698 (
            .O(N__21140),
            .I(N__21124));
    LocalMux I__3697 (
            .O(N__21129),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    Odrv4 I__3696 (
            .O(N__21124),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__3695 (
            .O(N__21119),
            .I(VCCST_EN_i_1_cascade_));
    CascadeMux I__3694 (
            .O(N__21116),
            .I(\POWERLED.un1_func_state25_6_0_o_N_5_cascade_ ));
    InMux I__3693 (
            .O(N__21113),
            .I(N__21110));
    LocalMux I__3692 (
            .O(N__21110),
            .I(\POWERLED.N_432 ));
    InMux I__3691 (
            .O(N__21107),
            .I(N__21104));
    LocalMux I__3690 (
            .O(N__21104),
            .I(\POWERLED.un1_func_state25_6_0_o_N_7_2 ));
    InMux I__3689 (
            .O(N__21101),
            .I(\POWERLED.un3_count_off_1_cry_14 ));
    InMux I__3688 (
            .O(N__21098),
            .I(N__21094));
    InMux I__3687 (
            .O(N__21097),
            .I(N__21091));
    LocalMux I__3686 (
            .O(N__21094),
            .I(N__21088));
    LocalMux I__3685 (
            .O(N__21091),
            .I(\POWERLED.count_off_1_12 ));
    Odrv4 I__3684 (
            .O(N__21088),
            .I(\POWERLED.count_off_1_12 ));
    InMux I__3683 (
            .O(N__21083),
            .I(N__21080));
    LocalMux I__3682 (
            .O(N__21080),
            .I(N__21077));
    Odrv4 I__3681 (
            .O(N__21077),
            .I(\POWERLED.count_off_0_12 ));
    InMux I__3680 (
            .O(N__21074),
            .I(N__21070));
    InMux I__3679 (
            .O(N__21073),
            .I(N__21067));
    LocalMux I__3678 (
            .O(N__21070),
            .I(\COUNTER.counterZ0Z_19 ));
    LocalMux I__3677 (
            .O(N__21067),
            .I(\COUNTER.counterZ0Z_19 ));
    InMux I__3676 (
            .O(N__21062),
            .I(N__21058));
    InMux I__3675 (
            .O(N__21061),
            .I(N__21055));
    LocalMux I__3674 (
            .O(N__21058),
            .I(\COUNTER.counterZ0Z_17 ));
    LocalMux I__3673 (
            .O(N__21055),
            .I(\COUNTER.counterZ0Z_17 ));
    CascadeMux I__3672 (
            .O(N__21050),
            .I(N__21046));
    InMux I__3671 (
            .O(N__21049),
            .I(N__21043));
    InMux I__3670 (
            .O(N__21046),
            .I(N__21040));
    LocalMux I__3669 (
            .O(N__21043),
            .I(\COUNTER.counterZ0Z_18 ));
    LocalMux I__3668 (
            .O(N__21040),
            .I(\COUNTER.counterZ0Z_18 ));
    InMux I__3667 (
            .O(N__21035),
            .I(N__21031));
    InMux I__3666 (
            .O(N__21034),
            .I(N__21028));
    LocalMux I__3665 (
            .O(N__21031),
            .I(\COUNTER.counterZ0Z_16 ));
    LocalMux I__3664 (
            .O(N__21028),
            .I(\COUNTER.counterZ0Z_16 ));
    InMux I__3663 (
            .O(N__21023),
            .I(N__21019));
    InMux I__3662 (
            .O(N__21022),
            .I(N__21016));
    LocalMux I__3661 (
            .O(N__21019),
            .I(\COUNTER.counterZ0Z_23 ));
    LocalMux I__3660 (
            .O(N__21016),
            .I(\COUNTER.counterZ0Z_23 ));
    InMux I__3659 (
            .O(N__21011),
            .I(N__21007));
    InMux I__3658 (
            .O(N__21010),
            .I(N__21004));
    LocalMux I__3657 (
            .O(N__21007),
            .I(\COUNTER.counterZ0Z_20 ));
    LocalMux I__3656 (
            .O(N__21004),
            .I(\COUNTER.counterZ0Z_20 ));
    CascadeMux I__3655 (
            .O(N__20999),
            .I(N__20995));
    InMux I__3654 (
            .O(N__20998),
            .I(N__20992));
    InMux I__3653 (
            .O(N__20995),
            .I(N__20989));
    LocalMux I__3652 (
            .O(N__20992),
            .I(\COUNTER.counterZ0Z_21 ));
    LocalMux I__3651 (
            .O(N__20989),
            .I(\COUNTER.counterZ0Z_21 ));
    InMux I__3650 (
            .O(N__20984),
            .I(N__20980));
    InMux I__3649 (
            .O(N__20983),
            .I(N__20977));
    LocalMux I__3648 (
            .O(N__20980),
            .I(\COUNTER.counterZ0Z_22 ));
    LocalMux I__3647 (
            .O(N__20977),
            .I(\COUNTER.counterZ0Z_22 ));
    CascadeMux I__3646 (
            .O(N__20972),
            .I(N__20969));
    InMux I__3645 (
            .O(N__20969),
            .I(N__20966));
    LocalMux I__3644 (
            .O(N__20966),
            .I(N__20963));
    Odrv4 I__3643 (
            .O(N__20963),
            .I(N_555));
    SRMux I__3642 (
            .O(N__20960),
            .I(N__20956));
    SRMux I__3641 (
            .O(N__20959),
            .I(N__20952));
    LocalMux I__3640 (
            .O(N__20956),
            .I(N__20949));
    SRMux I__3639 (
            .O(N__20955),
            .I(N__20946));
    LocalMux I__3638 (
            .O(N__20952),
            .I(N__20942));
    Span4Mux_s1_v I__3637 (
            .O(N__20949),
            .I(N__20937));
    LocalMux I__3636 (
            .O(N__20946),
            .I(N__20937));
    InMux I__3635 (
            .O(N__20945),
            .I(N__20934));
    Span4Mux_v I__3634 (
            .O(N__20942),
            .I(N__20931));
    Span4Mux_h I__3633 (
            .O(N__20937),
            .I(N__20926));
    LocalMux I__3632 (
            .O(N__20934),
            .I(N__20926));
    Span4Mux_h I__3631 (
            .O(N__20931),
            .I(N__20921));
    Span4Mux_v I__3630 (
            .O(N__20926),
            .I(N__20921));
    Odrv4 I__3629 (
            .O(N__20921),
            .I(G_14));
    InMux I__3628 (
            .O(N__20918),
            .I(N__20914));
    CascadeMux I__3627 (
            .O(N__20917),
            .I(N__20911));
    LocalMux I__3626 (
            .O(N__20914),
            .I(N__20907));
    InMux I__3625 (
            .O(N__20911),
            .I(N__20902));
    InMux I__3624 (
            .O(N__20910),
            .I(N__20902));
    Span4Mux_h I__3623 (
            .O(N__20907),
            .I(N__20897));
    LocalMux I__3622 (
            .O(N__20902),
            .I(N__20897));
    Sp12to4 I__3621 (
            .O(N__20897),
            .I(N__20894));
    Span12Mux_v I__3620 (
            .O(N__20894),
            .I(N__20891));
    Odrv12 I__3619 (
            .O(N__20891),
            .I(N_662));
    InMux I__3618 (
            .O(N__20888),
            .I(\POWERLED.un3_count_off_1_cry_6 ));
    InMux I__3617 (
            .O(N__20885),
            .I(\POWERLED.un3_count_off_1_cry_7 ));
    InMux I__3616 (
            .O(N__20882),
            .I(N__20879));
    LocalMux I__3615 (
            .O(N__20879),
            .I(N__20876));
    Odrv4 I__3614 (
            .O(N__20876),
            .I(\POWERLED.count_offZ0Z_9 ));
    InMux I__3613 (
            .O(N__20873),
            .I(N__20867));
    InMux I__3612 (
            .O(N__20872),
            .I(N__20867));
    LocalMux I__3611 (
            .O(N__20867),
            .I(N__20864));
    Odrv4 I__3610 (
            .O(N__20864),
            .I(\POWERLED.count_off_1_9 ));
    InMux I__3609 (
            .O(N__20861),
            .I(bfn_7_4_0_));
    CascadeMux I__3608 (
            .O(N__20858),
            .I(N__20855));
    InMux I__3607 (
            .O(N__20855),
            .I(N__20851));
    InMux I__3606 (
            .O(N__20854),
            .I(N__20848));
    LocalMux I__3605 (
            .O(N__20851),
            .I(N__20845));
    LocalMux I__3604 (
            .O(N__20848),
            .I(\POWERLED.count_offZ0Z_10 ));
    Odrv4 I__3603 (
            .O(N__20845),
            .I(\POWERLED.count_offZ0Z_10 ));
    InMux I__3602 (
            .O(N__20840),
            .I(N__20834));
    InMux I__3601 (
            .O(N__20839),
            .I(N__20834));
    LocalMux I__3600 (
            .O(N__20834),
            .I(N__20831));
    Odrv4 I__3599 (
            .O(N__20831),
            .I(\POWERLED.count_off_1_10 ));
    InMux I__3598 (
            .O(N__20828),
            .I(\POWERLED.un3_count_off_1_cry_9 ));
    InMux I__3597 (
            .O(N__20825),
            .I(N__20821));
    InMux I__3596 (
            .O(N__20824),
            .I(N__20818));
    LocalMux I__3595 (
            .O(N__20821),
            .I(N__20815));
    LocalMux I__3594 (
            .O(N__20818),
            .I(\POWERLED.count_offZ0Z_11 ));
    Odrv4 I__3593 (
            .O(N__20815),
            .I(\POWERLED.count_offZ0Z_11 ));
    InMux I__3592 (
            .O(N__20810),
            .I(N__20804));
    InMux I__3591 (
            .O(N__20809),
            .I(N__20804));
    LocalMux I__3590 (
            .O(N__20804),
            .I(N__20801));
    Odrv4 I__3589 (
            .O(N__20801),
            .I(\POWERLED.count_off_1_11 ));
    InMux I__3588 (
            .O(N__20798),
            .I(\POWERLED.un3_count_off_1_cry_10 ));
    InMux I__3587 (
            .O(N__20795),
            .I(N__20791));
    InMux I__3586 (
            .O(N__20794),
            .I(N__20788));
    LocalMux I__3585 (
            .O(N__20791),
            .I(N__20785));
    LocalMux I__3584 (
            .O(N__20788),
            .I(\POWERLED.count_offZ0Z_12 ));
    Odrv4 I__3583 (
            .O(N__20785),
            .I(\POWERLED.count_offZ0Z_12 ));
    InMux I__3582 (
            .O(N__20780),
            .I(\POWERLED.un3_count_off_1_cry_11 ));
    InMux I__3581 (
            .O(N__20777),
            .I(\POWERLED.un3_count_off_1_cry_12 ));
    InMux I__3580 (
            .O(N__20774),
            .I(\POWERLED.un3_count_off_1_cry_13 ));
    InMux I__3579 (
            .O(N__20771),
            .I(N__20768));
    LocalMux I__3578 (
            .O(N__20768),
            .I(\POWERLED.count_off_0_10 ));
    InMux I__3577 (
            .O(N__20765),
            .I(N__20762));
    LocalMux I__3576 (
            .O(N__20762),
            .I(\POWERLED.count_off_0_11 ));
    InMux I__3575 (
            .O(N__20759),
            .I(\POWERLED.un3_count_off_1_cry_1_cZ0 ));
    InMux I__3574 (
            .O(N__20756),
            .I(\POWERLED.un3_count_off_1_cry_2 ));
    InMux I__3573 (
            .O(N__20753),
            .I(\POWERLED.un3_count_off_1_cry_3 ));
    InMux I__3572 (
            .O(N__20750),
            .I(\POWERLED.un3_count_off_1_cry_4 ));
    InMux I__3571 (
            .O(N__20747),
            .I(\POWERLED.un3_count_off_1_cry_5 ));
    CascadeMux I__3570 (
            .O(N__20744),
            .I(N__20739));
    InMux I__3569 (
            .O(N__20743),
            .I(N__20735));
    InMux I__3568 (
            .O(N__20742),
            .I(N__20730));
    InMux I__3567 (
            .O(N__20739),
            .I(N__20730));
    InMux I__3566 (
            .O(N__20738),
            .I(N__20727));
    LocalMux I__3565 (
            .O(N__20735),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__3564 (
            .O(N__20730),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__3563 (
            .O(N__20727),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    CascadeMux I__3562 (
            .O(N__20720),
            .I(N__20717));
    InMux I__3561 (
            .O(N__20717),
            .I(N__20714));
    LocalMux I__3560 (
            .O(N__20714),
            .I(\POWERLED.mult1_un75_sum_cry_5_s ));
    InMux I__3559 (
            .O(N__20711),
            .I(N__20708));
    LocalMux I__3558 (
            .O(N__20708),
            .I(\POWERLED.mult1_un82_sum_cry_6_s ));
    InMux I__3557 (
            .O(N__20705),
            .I(\POWERLED.mult1_un82_sum_cry_5 ));
    InMux I__3556 (
            .O(N__20702),
            .I(N__20699));
    LocalMux I__3555 (
            .O(N__20699),
            .I(\POWERLED.mult1_un75_sum_cry_6_s ));
    CascadeMux I__3554 (
            .O(N__20696),
            .I(N__20692));
    CascadeMux I__3553 (
            .O(N__20695),
            .I(N__20688));
    InMux I__3552 (
            .O(N__20692),
            .I(N__20681));
    InMux I__3551 (
            .O(N__20691),
            .I(N__20681));
    InMux I__3550 (
            .O(N__20688),
            .I(N__20681));
    LocalMux I__3549 (
            .O(N__20681),
            .I(\POWERLED.mult1_un75_sum_i_0_8 ));
    CascadeMux I__3548 (
            .O(N__20678),
            .I(N__20675));
    InMux I__3547 (
            .O(N__20675),
            .I(N__20672));
    LocalMux I__3546 (
            .O(N__20672),
            .I(\POWERLED.mult1_un89_sum_axb_8 ));
    InMux I__3545 (
            .O(N__20669),
            .I(\POWERLED.mult1_un82_sum_cry_6 ));
    CascadeMux I__3544 (
            .O(N__20666),
            .I(N__20663));
    InMux I__3543 (
            .O(N__20663),
            .I(N__20660));
    LocalMux I__3542 (
            .O(N__20660),
            .I(\POWERLED.mult1_un82_sum_axb_8 ));
    InMux I__3541 (
            .O(N__20657),
            .I(\POWERLED.mult1_un82_sum_cry_7 ));
    CascadeMux I__3540 (
            .O(N__20654),
            .I(N__20650));
    InMux I__3539 (
            .O(N__20653),
            .I(N__20642));
    InMux I__3538 (
            .O(N__20650),
            .I(N__20642));
    InMux I__3537 (
            .O(N__20649),
            .I(N__20639));
    InMux I__3536 (
            .O(N__20648),
            .I(N__20634));
    InMux I__3535 (
            .O(N__20647),
            .I(N__20634));
    LocalMux I__3534 (
            .O(N__20642),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__3533 (
            .O(N__20639),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__3532 (
            .O(N__20634),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    InMux I__3531 (
            .O(N__20627),
            .I(N__20624));
    LocalMux I__3530 (
            .O(N__20624),
            .I(\POWERLED.mult1_un75_sum_i ));
    InMux I__3529 (
            .O(N__20621),
            .I(N__20618));
    LocalMux I__3528 (
            .O(N__20618),
            .I(\POWERLED.count_off_0_9 ));
    CascadeMux I__3527 (
            .O(N__20615),
            .I(\POWERLED.count_offZ0Z_9_cascade_ ));
    InMux I__3526 (
            .O(N__20612),
            .I(N__20609));
    LocalMux I__3525 (
            .O(N__20609),
            .I(\POWERLED.mult1_un68_sum_cry_4_s ));
    InMux I__3524 (
            .O(N__20606),
            .I(\POWERLED.mult1_un75_sum_cry_4 ));
    InMux I__3523 (
            .O(N__20603),
            .I(N__20600));
    LocalMux I__3522 (
            .O(N__20600),
            .I(N__20596));
    CascadeMux I__3521 (
            .O(N__20599),
            .I(N__20592));
    Span4Mux_s2_v I__3520 (
            .O(N__20596),
            .I(N__20588));
    InMux I__3519 (
            .O(N__20595),
            .I(N__20583));
    InMux I__3518 (
            .O(N__20592),
            .I(N__20583));
    InMux I__3517 (
            .O(N__20591),
            .I(N__20580));
    Odrv4 I__3516 (
            .O(N__20588),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__3515 (
            .O(N__20583),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__3514 (
            .O(N__20580),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    CascadeMux I__3513 (
            .O(N__20573),
            .I(N__20570));
    InMux I__3512 (
            .O(N__20570),
            .I(N__20567));
    LocalMux I__3511 (
            .O(N__20567),
            .I(\POWERLED.mult1_un68_sum_cry_5_s ));
    InMux I__3510 (
            .O(N__20564),
            .I(\POWERLED.mult1_un75_sum_cry_5 ));
    InMux I__3509 (
            .O(N__20561),
            .I(N__20558));
    LocalMux I__3508 (
            .O(N__20558),
            .I(\POWERLED.mult1_un68_sum_cry_6_s ));
    CascadeMux I__3507 (
            .O(N__20555),
            .I(N__20551));
    CascadeMux I__3506 (
            .O(N__20554),
            .I(N__20547));
    InMux I__3505 (
            .O(N__20551),
            .I(N__20540));
    InMux I__3504 (
            .O(N__20550),
            .I(N__20540));
    InMux I__3503 (
            .O(N__20547),
            .I(N__20540));
    LocalMux I__3502 (
            .O(N__20540),
            .I(\POWERLED.mult1_un68_sum_i_0_8 ));
    InMux I__3501 (
            .O(N__20537),
            .I(\POWERLED.mult1_un75_sum_cry_6 ));
    CascadeMux I__3500 (
            .O(N__20534),
            .I(N__20531));
    InMux I__3499 (
            .O(N__20531),
            .I(N__20528));
    LocalMux I__3498 (
            .O(N__20528),
            .I(\POWERLED.mult1_un75_sum_axb_8 ));
    InMux I__3497 (
            .O(N__20525),
            .I(\POWERLED.mult1_un75_sum_cry_7 ));
    CascadeMux I__3496 (
            .O(N__20522),
            .I(\POWERLED.mult1_un75_sum_s_8_cascade_ ));
    CascadeMux I__3495 (
            .O(N__20519),
            .I(N__20516));
    InMux I__3494 (
            .O(N__20516),
            .I(N__20513));
    LocalMux I__3493 (
            .O(N__20513),
            .I(\POWERLED.mult1_un82_sum_cry_3_s ));
    InMux I__3492 (
            .O(N__20510),
            .I(\POWERLED.mult1_un82_sum_cry_2 ));
    CascadeMux I__3491 (
            .O(N__20507),
            .I(N__20504));
    InMux I__3490 (
            .O(N__20504),
            .I(N__20501));
    LocalMux I__3489 (
            .O(N__20501),
            .I(\POWERLED.mult1_un75_sum_cry_3_s ));
    InMux I__3488 (
            .O(N__20498),
            .I(N__20495));
    LocalMux I__3487 (
            .O(N__20495),
            .I(\POWERLED.mult1_un82_sum_cry_4_s ));
    InMux I__3486 (
            .O(N__20492),
            .I(\POWERLED.mult1_un82_sum_cry_3 ));
    InMux I__3485 (
            .O(N__20489),
            .I(N__20486));
    LocalMux I__3484 (
            .O(N__20486),
            .I(\POWERLED.mult1_un75_sum_cry_4_s ));
    CascadeMux I__3483 (
            .O(N__20483),
            .I(N__20480));
    InMux I__3482 (
            .O(N__20480),
            .I(N__20477));
    LocalMux I__3481 (
            .O(N__20477),
            .I(\POWERLED.mult1_un82_sum_cry_5_s ));
    InMux I__3480 (
            .O(N__20474),
            .I(\POWERLED.mult1_un82_sum_cry_4 ));
    InMux I__3479 (
            .O(N__20471),
            .I(\POWERLED.mult1_un68_sum_cry_3 ));
    InMux I__3478 (
            .O(N__20468),
            .I(\POWERLED.mult1_un68_sum_cry_4 ));
    InMux I__3477 (
            .O(N__20465),
            .I(\POWERLED.mult1_un68_sum_cry_5 ));
    CascadeMux I__3476 (
            .O(N__20462),
            .I(N__20458));
    CascadeMux I__3475 (
            .O(N__20461),
            .I(N__20454));
    InMux I__3474 (
            .O(N__20458),
            .I(N__20447));
    InMux I__3473 (
            .O(N__20457),
            .I(N__20447));
    InMux I__3472 (
            .O(N__20454),
            .I(N__20447));
    LocalMux I__3471 (
            .O(N__20447),
            .I(\POWERLED.mult1_un61_sum_i_0_8 ));
    InMux I__3470 (
            .O(N__20444),
            .I(\POWERLED.mult1_un68_sum_cry_6 ));
    InMux I__3469 (
            .O(N__20441),
            .I(\POWERLED.mult1_un68_sum_cry_7 ));
    CascadeMux I__3468 (
            .O(N__20438),
            .I(\POWERLED.mult1_un68_sum_s_8_cascade_ ));
    InMux I__3467 (
            .O(N__20435),
            .I(\POWERLED.mult1_un75_sum_cry_2 ));
    CascadeMux I__3466 (
            .O(N__20432),
            .I(N__20429));
    InMux I__3465 (
            .O(N__20429),
            .I(N__20426));
    LocalMux I__3464 (
            .O(N__20426),
            .I(\POWERLED.mult1_un68_sum_cry_3_s ));
    InMux I__3463 (
            .O(N__20423),
            .I(\POWERLED.mult1_un75_sum_cry_3 ));
    InMux I__3462 (
            .O(N__20420),
            .I(N__20417));
    LocalMux I__3461 (
            .O(N__20417),
            .I(N__20414));
    Odrv4 I__3460 (
            .O(N__20414),
            .I(\POWERLED.mult1_un131_sum_i ));
    CascadeMux I__3459 (
            .O(N__20411),
            .I(N__20408));
    InMux I__3458 (
            .O(N__20408),
            .I(N__20405));
    LocalMux I__3457 (
            .O(N__20405),
            .I(N__20402));
    Odrv4 I__3456 (
            .O(N__20402),
            .I(\POWERLED.mult1_un145_sum_i ));
    InMux I__3455 (
            .O(N__20399),
            .I(N__20396));
    LocalMux I__3454 (
            .O(N__20396),
            .I(N__20393));
    Span4Mux_h I__3453 (
            .O(N__20393),
            .I(N__20390));
    Odrv4 I__3452 (
            .O(N__20390),
            .I(\POWERLED.mult1_un103_sum_i ));
    InMux I__3451 (
            .O(N__20387),
            .I(N__20384));
    LocalMux I__3450 (
            .O(N__20384),
            .I(N__20381));
    Odrv4 I__3449 (
            .O(N__20381),
            .I(\POWERLED.mult1_un124_sum_i ));
    InMux I__3448 (
            .O(N__20378),
            .I(N__20375));
    LocalMux I__3447 (
            .O(N__20375),
            .I(N__20372));
    Span4Mux_v I__3446 (
            .O(N__20372),
            .I(N__20369));
    Odrv4 I__3445 (
            .O(N__20369),
            .I(\POWERLED.mult1_un110_sum_i ));
    InMux I__3444 (
            .O(N__20366),
            .I(N__20363));
    LocalMux I__3443 (
            .O(N__20363),
            .I(N__20360));
    Span4Mux_s3_v I__3442 (
            .O(N__20360),
            .I(N__20357));
    Odrv4 I__3441 (
            .O(N__20357),
            .I(\POWERLED.mult1_un61_sum_i_8 ));
    InMux I__3440 (
            .O(N__20354),
            .I(\POWERLED.mult1_un68_sum_cry_2 ));
    CascadeMux I__3439 (
            .O(N__20351),
            .I(N__20348));
    InMux I__3438 (
            .O(N__20348),
            .I(N__20345));
    LocalMux I__3437 (
            .O(N__20345),
            .I(\POWERLED.mult1_un159_sum_cry_2_s ));
    InMux I__3436 (
            .O(N__20342),
            .I(\POWERLED.mult1_un159_sum_cry_1 ));
    InMux I__3435 (
            .O(N__20339),
            .I(N__20336));
    LocalMux I__3434 (
            .O(N__20336),
            .I(\POWERLED.mult1_un152_sum_cry_3_s ));
    CascadeMux I__3433 (
            .O(N__20333),
            .I(N__20330));
    InMux I__3432 (
            .O(N__20330),
            .I(N__20327));
    LocalMux I__3431 (
            .O(N__20327),
            .I(\POWERLED.mult1_un159_sum_cry_3_s ));
    InMux I__3430 (
            .O(N__20324),
            .I(\POWERLED.mult1_un159_sum_cry_2 ));
    InMux I__3429 (
            .O(N__20321),
            .I(N__20318));
    LocalMux I__3428 (
            .O(N__20318),
            .I(\POWERLED.mult1_un152_sum_cry_4_s ));
    InMux I__3427 (
            .O(N__20315),
            .I(N__20312));
    LocalMux I__3426 (
            .O(N__20312),
            .I(\POWERLED.mult1_un159_sum_cry_4_s ));
    InMux I__3425 (
            .O(N__20309),
            .I(\POWERLED.mult1_un159_sum_cry_3 ));
    InMux I__3424 (
            .O(N__20306),
            .I(N__20303));
    LocalMux I__3423 (
            .O(N__20303),
            .I(\POWERLED.mult1_un152_sum_cry_5_s ));
    InMux I__3422 (
            .O(N__20300),
            .I(N__20297));
    LocalMux I__3421 (
            .O(N__20297),
            .I(\POWERLED.mult1_un159_sum_cry_5_s ));
    InMux I__3420 (
            .O(N__20294),
            .I(\POWERLED.mult1_un159_sum_cry_4 ));
    InMux I__3419 (
            .O(N__20291),
            .I(N__20288));
    LocalMux I__3418 (
            .O(N__20288),
            .I(\POWERLED.mult1_un152_sum_cry_6_s ));
    InMux I__3417 (
            .O(N__20285),
            .I(N__20282));
    LocalMux I__3416 (
            .O(N__20282),
            .I(\POWERLED.mult1_un166_sum_axb_6 ));
    InMux I__3415 (
            .O(N__20279),
            .I(\POWERLED.mult1_un159_sum_cry_5 ));
    InMux I__3414 (
            .O(N__20276),
            .I(N__20273));
    LocalMux I__3413 (
            .O(N__20273),
            .I(\POWERLED.mult1_un159_sum_axb_7 ));
    InMux I__3412 (
            .O(N__20270),
            .I(\POWERLED.mult1_un159_sum_cry_6 ));
    InMux I__3411 (
            .O(N__20267),
            .I(N__20263));
    CascadeMux I__3410 (
            .O(N__20266),
            .I(N__20260));
    LocalMux I__3409 (
            .O(N__20263),
            .I(N__20254));
    InMux I__3408 (
            .O(N__20260),
            .I(N__20247));
    InMux I__3407 (
            .O(N__20259),
            .I(N__20247));
    InMux I__3406 (
            .O(N__20258),
            .I(N__20247));
    InMux I__3405 (
            .O(N__20257),
            .I(N__20244));
    Odrv4 I__3404 (
            .O(N__20254),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__3403 (
            .O(N__20247),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__3402 (
            .O(N__20244),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    CascadeMux I__3401 (
            .O(N__20237),
            .I(N__20232));
    CascadeMux I__3400 (
            .O(N__20236),
            .I(N__20229));
    InMux I__3399 (
            .O(N__20235),
            .I(N__20224));
    InMux I__3398 (
            .O(N__20232),
            .I(N__20221));
    InMux I__3397 (
            .O(N__20229),
            .I(N__20216));
    InMux I__3396 (
            .O(N__20228),
            .I(N__20216));
    InMux I__3395 (
            .O(N__20227),
            .I(N__20213));
    LocalMux I__3394 (
            .O(N__20224),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__3393 (
            .O(N__20221),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__3392 (
            .O(N__20216),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__3391 (
            .O(N__20213),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    CascadeMux I__3390 (
            .O(N__20204),
            .I(N__20200));
    CascadeMux I__3389 (
            .O(N__20203),
            .I(N__20197));
    InMux I__3388 (
            .O(N__20200),
            .I(N__20193));
    InMux I__3387 (
            .O(N__20197),
            .I(N__20188));
    InMux I__3386 (
            .O(N__20196),
            .I(N__20188));
    LocalMux I__3385 (
            .O(N__20193),
            .I(\POWERLED.mult1_un152_sum_i_0_8 ));
    LocalMux I__3384 (
            .O(N__20188),
            .I(\POWERLED.mult1_un152_sum_i_0_8 ));
    CascadeMux I__3383 (
            .O(N__20183),
            .I(N__20180));
    InMux I__3382 (
            .O(N__20180),
            .I(N__20177));
    LocalMux I__3381 (
            .O(N__20177),
            .I(N__20174));
    Odrv4 I__3380 (
            .O(N__20174),
            .I(\POWERLED.mult1_un138_sum_i ));
    InMux I__3379 (
            .O(N__20171),
            .I(\POWERLED.mult1_un152_sum_cry_2 ));
    InMux I__3378 (
            .O(N__20168),
            .I(N__20165));
    LocalMux I__3377 (
            .O(N__20165),
            .I(\POWERLED.mult1_un145_sum_cry_3_s ));
    InMux I__3376 (
            .O(N__20162),
            .I(\POWERLED.mult1_un152_sum_cry_3 ));
    CascadeMux I__3375 (
            .O(N__20159),
            .I(N__20156));
    InMux I__3374 (
            .O(N__20156),
            .I(N__20153));
    LocalMux I__3373 (
            .O(N__20153),
            .I(\POWERLED.mult1_un145_sum_cry_4_s ));
    InMux I__3372 (
            .O(N__20150),
            .I(\POWERLED.mult1_un152_sum_cry_4 ));
    InMux I__3371 (
            .O(N__20147),
            .I(N__20144));
    LocalMux I__3370 (
            .O(N__20144),
            .I(\POWERLED.mult1_un145_sum_cry_5_s ));
    InMux I__3369 (
            .O(N__20141),
            .I(N__20137));
    CascadeMux I__3368 (
            .O(N__20140),
            .I(N__20134));
    LocalMux I__3367 (
            .O(N__20137),
            .I(N__20129));
    InMux I__3366 (
            .O(N__20134),
            .I(N__20124));
    InMux I__3365 (
            .O(N__20133),
            .I(N__20124));
    InMux I__3364 (
            .O(N__20132),
            .I(N__20121));
    Odrv4 I__3363 (
            .O(N__20129),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__3362 (
            .O(N__20124),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__3361 (
            .O(N__20121),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    InMux I__3360 (
            .O(N__20114),
            .I(\POWERLED.mult1_un152_sum_cry_5 ));
    CascadeMux I__3359 (
            .O(N__20111),
            .I(N__20107));
    InMux I__3358 (
            .O(N__20110),
            .I(N__20099));
    InMux I__3357 (
            .O(N__20107),
            .I(N__20099));
    InMux I__3356 (
            .O(N__20106),
            .I(N__20099));
    LocalMux I__3355 (
            .O(N__20099),
            .I(\POWERLED.mult1_un145_sum_i_0_8 ));
    CascadeMux I__3354 (
            .O(N__20096),
            .I(N__20093));
    InMux I__3353 (
            .O(N__20093),
            .I(N__20090));
    LocalMux I__3352 (
            .O(N__20090),
            .I(N__20087));
    Odrv4 I__3351 (
            .O(N__20087),
            .I(\POWERLED.mult1_un145_sum_cry_6_s ));
    InMux I__3350 (
            .O(N__20084),
            .I(\POWERLED.mult1_un152_sum_cry_6 ));
    InMux I__3349 (
            .O(N__20081),
            .I(N__20078));
    LocalMux I__3348 (
            .O(N__20078),
            .I(\POWERLED.mult1_un152_sum_axb_8 ));
    InMux I__3347 (
            .O(N__20075),
            .I(\POWERLED.mult1_un152_sum_cry_7 ));
    InMux I__3346 (
            .O(N__20072),
            .I(N__20068));
    CascadeMux I__3345 (
            .O(N__20071),
            .I(N__20064));
    LocalMux I__3344 (
            .O(N__20068),
            .I(N__20059));
    InMux I__3343 (
            .O(N__20067),
            .I(N__20056));
    InMux I__3342 (
            .O(N__20064),
            .I(N__20051));
    InMux I__3341 (
            .O(N__20063),
            .I(N__20051));
    InMux I__3340 (
            .O(N__20062),
            .I(N__20048));
    Odrv12 I__3339 (
            .O(N__20059),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__3338 (
            .O(N__20056),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__3337 (
            .O(N__20051),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__3336 (
            .O(N__20048),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    CascadeMux I__3335 (
            .O(N__20039),
            .I(N__20034));
    CascadeMux I__3334 (
            .O(N__20038),
            .I(N__20031));
    CascadeMux I__3333 (
            .O(N__20037),
            .I(N__20028));
    InMux I__3332 (
            .O(N__20034),
            .I(N__20025));
    InMux I__3331 (
            .O(N__20031),
            .I(N__20020));
    InMux I__3330 (
            .O(N__20028),
            .I(N__20020));
    LocalMux I__3329 (
            .O(N__20025),
            .I(\POWERLED.mult1_un131_sum_i_0_8 ));
    LocalMux I__3328 (
            .O(N__20020),
            .I(\POWERLED.mult1_un131_sum_i_0_8 ));
    InMux I__3327 (
            .O(N__20015),
            .I(N__20012));
    LocalMux I__3326 (
            .O(N__20012),
            .I(\POWERLED.mult1_un138_sum_cry_3_s ));
    InMux I__3325 (
            .O(N__20009),
            .I(\POWERLED.mult1_un138_sum_cry_2 ));
    InMux I__3324 (
            .O(N__20006),
            .I(N__20003));
    LocalMux I__3323 (
            .O(N__20003),
            .I(\POWERLED.mult1_un131_sum_cry_3_s ));
    CascadeMux I__3322 (
            .O(N__20000),
            .I(N__19997));
    InMux I__3321 (
            .O(N__19997),
            .I(N__19994));
    LocalMux I__3320 (
            .O(N__19994),
            .I(\POWERLED.mult1_un138_sum_cry_4_s ));
    InMux I__3319 (
            .O(N__19991),
            .I(\POWERLED.mult1_un138_sum_cry_3 ));
    CascadeMux I__3318 (
            .O(N__19988),
            .I(N__19985));
    InMux I__3317 (
            .O(N__19985),
            .I(N__19982));
    LocalMux I__3316 (
            .O(N__19982),
            .I(\POWERLED.mult1_un131_sum_cry_4_s ));
    InMux I__3315 (
            .O(N__19979),
            .I(N__19976));
    LocalMux I__3314 (
            .O(N__19976),
            .I(\POWERLED.mult1_un138_sum_cry_5_s ));
    InMux I__3313 (
            .O(N__19973),
            .I(\POWERLED.mult1_un138_sum_cry_4 ));
    InMux I__3312 (
            .O(N__19970),
            .I(N__19967));
    LocalMux I__3311 (
            .O(N__19967),
            .I(\POWERLED.mult1_un131_sum_cry_5_s ));
    CascadeMux I__3310 (
            .O(N__19964),
            .I(N__19961));
    InMux I__3309 (
            .O(N__19961),
            .I(N__19958));
    LocalMux I__3308 (
            .O(N__19958),
            .I(\POWERLED.mult1_un138_sum_cry_6_s ));
    InMux I__3307 (
            .O(N__19955),
            .I(\POWERLED.mult1_un138_sum_cry_5 ));
    InMux I__3306 (
            .O(N__19952),
            .I(N__19949));
    LocalMux I__3305 (
            .O(N__19949),
            .I(\POWERLED.mult1_un131_sum_cry_6_s ));
    InMux I__3304 (
            .O(N__19946),
            .I(N__19943));
    LocalMux I__3303 (
            .O(N__19943),
            .I(\POWERLED.mult1_un145_sum_axb_8 ));
    InMux I__3302 (
            .O(N__19940),
            .I(\POWERLED.mult1_un138_sum_cry_6 ));
    InMux I__3301 (
            .O(N__19937),
            .I(N__19934));
    LocalMux I__3300 (
            .O(N__19934),
            .I(\POWERLED.mult1_un138_sum_axb_8 ));
    InMux I__3299 (
            .O(N__19931),
            .I(\POWERLED.mult1_un138_sum_cry_7 ));
    InMux I__3298 (
            .O(N__19928),
            .I(N__19925));
    LocalMux I__3297 (
            .O(N__19925),
            .I(N__19921));
    CascadeMux I__3296 (
            .O(N__19924),
            .I(N__19918));
    Span4Mux_v I__3295 (
            .O(N__19921),
            .I(N__19913));
    InMux I__3294 (
            .O(N__19918),
            .I(N__19908));
    InMux I__3293 (
            .O(N__19917),
            .I(N__19908));
    InMux I__3292 (
            .O(N__19916),
            .I(N__19905));
    Odrv4 I__3291 (
            .O(N__19913),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__3290 (
            .O(N__19908),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__3289 (
            .O(N__19905),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    CascadeMux I__3288 (
            .O(N__19898),
            .I(\POWERLED.mult1_un138_sum_s_8_cascade_ ));
    CascadeMux I__3287 (
            .O(N__19895),
            .I(N__19891));
    InMux I__3286 (
            .O(N__19894),
            .I(N__19883));
    InMux I__3285 (
            .O(N__19891),
            .I(N__19883));
    InMux I__3284 (
            .O(N__19890),
            .I(N__19883));
    LocalMux I__3283 (
            .O(N__19883),
            .I(\POWERLED.mult1_un138_sum_i_0_8 ));
    InMux I__3282 (
            .O(N__19880),
            .I(N__19877));
    LocalMux I__3281 (
            .O(N__19877),
            .I(\VPP_VDDQ.un1_count_2_1_axb_6 ));
    InMux I__3280 (
            .O(N__19874),
            .I(N__19871));
    LocalMux I__3279 (
            .O(N__19871),
            .I(\VPP_VDDQ.count_2_0_4 ));
    InMux I__3278 (
            .O(N__19868),
            .I(N__19862));
    InMux I__3277 (
            .O(N__19867),
            .I(N__19862));
    LocalMux I__3276 (
            .O(N__19862),
            .I(\VPP_VDDQ.count_2_1_4 ));
    InMux I__3275 (
            .O(N__19859),
            .I(N__19856));
    LocalMux I__3274 (
            .O(N__19856),
            .I(\VPP_VDDQ.count_2Z0Z_4 ));
    InMux I__3273 (
            .O(N__19853),
            .I(N__19847));
    InMux I__3272 (
            .O(N__19852),
            .I(N__19847));
    LocalMux I__3271 (
            .O(N__19847),
            .I(\VPP_VDDQ.count_2Z0Z_6 ));
    CascadeMux I__3270 (
            .O(N__19844),
            .I(\VPP_VDDQ.count_2Z0Z_4_cascade_ ));
    InMux I__3269 (
            .O(N__19841),
            .I(N__19832));
    InMux I__3268 (
            .O(N__19840),
            .I(N__19832));
    InMux I__3267 (
            .O(N__19839),
            .I(N__19832));
    LocalMux I__3266 (
            .O(N__19832),
            .I(\VPP_VDDQ.count_2_1_6 ));
    InMux I__3265 (
            .O(N__19829),
            .I(N__19826));
    LocalMux I__3264 (
            .O(N__19826),
            .I(N__19823));
    Span4Mux_v I__3263 (
            .O(N__19823),
            .I(N__19820));
    Odrv4 I__3262 (
            .O(N__19820),
            .I(\VPP_VDDQ.un9_clk_100khz_0 ));
    InMux I__3261 (
            .O(N__19817),
            .I(N__19814));
    LocalMux I__3260 (
            .O(N__19814),
            .I(\VPP_VDDQ.count_2_0_2 ));
    InMux I__3259 (
            .O(N__19811),
            .I(N__19805));
    InMux I__3258 (
            .O(N__19810),
            .I(N__19805));
    LocalMux I__3257 (
            .O(N__19805),
            .I(\VPP_VDDQ.count_2_1_2 ));
    InMux I__3256 (
            .O(N__19802),
            .I(N__19789));
    InMux I__3255 (
            .O(N__19801),
            .I(N__19789));
    InMux I__3254 (
            .O(N__19800),
            .I(N__19789));
    CEMux I__3253 (
            .O(N__19799),
            .I(N__19789));
    CEMux I__3252 (
            .O(N__19798),
            .I(N__19786));
    LocalMux I__3251 (
            .O(N__19789),
            .I(N__19767));
    LocalMux I__3250 (
            .O(N__19786),
            .I(N__19767));
    InMux I__3249 (
            .O(N__19785),
            .I(N__19754));
    InMux I__3248 (
            .O(N__19784),
            .I(N__19754));
    InMux I__3247 (
            .O(N__19783),
            .I(N__19754));
    InMux I__3246 (
            .O(N__19782),
            .I(N__19754));
    CEMux I__3245 (
            .O(N__19781),
            .I(N__19750));
    CEMux I__3244 (
            .O(N__19780),
            .I(N__19747));
    InMux I__3243 (
            .O(N__19779),
            .I(N__19738));
    InMux I__3242 (
            .O(N__19778),
            .I(N__19738));
    InMux I__3241 (
            .O(N__19777),
            .I(N__19738));
    CEMux I__3240 (
            .O(N__19776),
            .I(N__19738));
    InMux I__3239 (
            .O(N__19775),
            .I(N__19729));
    InMux I__3238 (
            .O(N__19774),
            .I(N__19729));
    InMux I__3237 (
            .O(N__19773),
            .I(N__19729));
    InMux I__3236 (
            .O(N__19772),
            .I(N__19729));
    Span4Mux_h I__3235 (
            .O(N__19767),
            .I(N__19726));
    InMux I__3234 (
            .O(N__19766),
            .I(N__19717));
    CEMux I__3233 (
            .O(N__19765),
            .I(N__19717));
    InMux I__3232 (
            .O(N__19764),
            .I(N__19717));
    InMux I__3231 (
            .O(N__19763),
            .I(N__19717));
    LocalMux I__3230 (
            .O(N__19754),
            .I(N__19714));
    InMux I__3229 (
            .O(N__19753),
            .I(N__19711));
    LocalMux I__3228 (
            .O(N__19750),
            .I(N__19706));
    LocalMux I__3227 (
            .O(N__19747),
            .I(N__19706));
    LocalMux I__3226 (
            .O(N__19738),
            .I(N__19701));
    LocalMux I__3225 (
            .O(N__19729),
            .I(N__19701));
    Span4Mux_s3_h I__3224 (
            .O(N__19726),
            .I(N__19694));
    LocalMux I__3223 (
            .O(N__19717),
            .I(N__19694));
    Span4Mux_h I__3222 (
            .O(N__19714),
            .I(N__19694));
    LocalMux I__3221 (
            .O(N__19711),
            .I(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0 ));
    Odrv4 I__3220 (
            .O(N__19706),
            .I(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0 ));
    Odrv4 I__3219 (
            .O(N__19701),
            .I(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0 ));
    Odrv4 I__3218 (
            .O(N__19694),
            .I(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0 ));
    InMux I__3217 (
            .O(N__19685),
            .I(N__19682));
    LocalMux I__3216 (
            .O(N__19682),
            .I(\VPP_VDDQ.count_2Z0Z_2 ));
    InMux I__3215 (
            .O(N__19679),
            .I(N__19676));
    LocalMux I__3214 (
            .O(N__19676),
            .I(N__19673));
    Span4Mux_v I__3213 (
            .O(N__19673),
            .I(N__19669));
    InMux I__3212 (
            .O(N__19672),
            .I(N__19666));
    Odrv4 I__3211 (
            .O(N__19669),
            .I(\VPP_VDDQ.count_2Z0Z_5 ));
    LocalMux I__3210 (
            .O(N__19666),
            .I(\VPP_VDDQ.count_2Z0Z_5 ));
    InMux I__3209 (
            .O(N__19661),
            .I(N__19658));
    LocalMux I__3208 (
            .O(N__19658),
            .I(N__19654));
    CascadeMux I__3207 (
            .O(N__19657),
            .I(N__19651));
    Span12Mux_s8_h I__3206 (
            .O(N__19654),
            .I(N__19648));
    InMux I__3205 (
            .O(N__19651),
            .I(N__19645));
    Odrv12 I__3204 (
            .O(N__19648),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    LocalMux I__3203 (
            .O(N__19645),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    CascadeMux I__3202 (
            .O(N__19640),
            .I(\VPP_VDDQ.count_2Z0Z_2_cascade_ ));
    InMux I__3201 (
            .O(N__19637),
            .I(N__19634));
    LocalMux I__3200 (
            .O(N__19634),
            .I(N__19631));
    Span4Mux_v I__3199 (
            .O(N__19631),
            .I(N__19627));
    InMux I__3198 (
            .O(N__19630),
            .I(N__19624));
    Odrv4 I__3197 (
            .O(N__19627),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    LocalMux I__3196 (
            .O(N__19624),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    InMux I__3195 (
            .O(N__19619),
            .I(N__19616));
    LocalMux I__3194 (
            .O(N__19616),
            .I(N__19613));
    Span4Mux_h I__3193 (
            .O(N__19613),
            .I(N__19610));
    Odrv4 I__3192 (
            .O(N__19610),
            .I(\VPP_VDDQ.un9_clk_100khz_9 ));
    InMux I__3191 (
            .O(N__19607),
            .I(\COUNTER.counter_1_cry_22 ));
    InMux I__3190 (
            .O(N__19604),
            .I(N__19600));
    InMux I__3189 (
            .O(N__19603),
            .I(N__19597));
    LocalMux I__3188 (
            .O(N__19600),
            .I(\COUNTER.counterZ0Z_24 ));
    LocalMux I__3187 (
            .O(N__19597),
            .I(\COUNTER.counterZ0Z_24 ));
    InMux I__3186 (
            .O(N__19592),
            .I(\COUNTER.counter_1_cry_23 ));
    InMux I__3185 (
            .O(N__19589),
            .I(N__19585));
    InMux I__3184 (
            .O(N__19588),
            .I(N__19582));
    LocalMux I__3183 (
            .O(N__19585),
            .I(\COUNTER.counterZ0Z_25 ));
    LocalMux I__3182 (
            .O(N__19582),
            .I(\COUNTER.counterZ0Z_25 ));
    InMux I__3181 (
            .O(N__19577),
            .I(bfn_6_7_0_));
    CascadeMux I__3180 (
            .O(N__19574),
            .I(N__19570));
    InMux I__3179 (
            .O(N__19573),
            .I(N__19567));
    InMux I__3178 (
            .O(N__19570),
            .I(N__19564));
    LocalMux I__3177 (
            .O(N__19567),
            .I(\COUNTER.counterZ0Z_26 ));
    LocalMux I__3176 (
            .O(N__19564),
            .I(\COUNTER.counterZ0Z_26 ));
    InMux I__3175 (
            .O(N__19559),
            .I(\COUNTER.counter_1_cry_25 ));
    InMux I__3174 (
            .O(N__19556),
            .I(N__19552));
    InMux I__3173 (
            .O(N__19555),
            .I(N__19549));
    LocalMux I__3172 (
            .O(N__19552),
            .I(\COUNTER.counterZ0Z_27 ));
    LocalMux I__3171 (
            .O(N__19549),
            .I(\COUNTER.counterZ0Z_27 ));
    InMux I__3170 (
            .O(N__19544),
            .I(\COUNTER.counter_1_cry_26 ));
    CascadeMux I__3169 (
            .O(N__19541),
            .I(N__19538));
    InMux I__3168 (
            .O(N__19538),
            .I(N__19534));
    InMux I__3167 (
            .O(N__19537),
            .I(N__19531));
    LocalMux I__3166 (
            .O(N__19534),
            .I(N__19528));
    LocalMux I__3165 (
            .O(N__19531),
            .I(\COUNTER.counterZ0Z_28 ));
    Odrv12 I__3164 (
            .O(N__19528),
            .I(\COUNTER.counterZ0Z_28 ));
    InMux I__3163 (
            .O(N__19523),
            .I(\COUNTER.counter_1_cry_27 ));
    InMux I__3162 (
            .O(N__19520),
            .I(N__19516));
    InMux I__3161 (
            .O(N__19519),
            .I(N__19513));
    LocalMux I__3160 (
            .O(N__19516),
            .I(N__19510));
    LocalMux I__3159 (
            .O(N__19513),
            .I(\COUNTER.counterZ0Z_29 ));
    Odrv12 I__3158 (
            .O(N__19510),
            .I(\COUNTER.counterZ0Z_29 ));
    InMux I__3157 (
            .O(N__19505),
            .I(\COUNTER.counter_1_cry_28 ));
    InMux I__3156 (
            .O(N__19502),
            .I(N__19498));
    InMux I__3155 (
            .O(N__19501),
            .I(N__19495));
    LocalMux I__3154 (
            .O(N__19498),
            .I(N__19492));
    LocalMux I__3153 (
            .O(N__19495),
            .I(\COUNTER.counterZ0Z_30 ));
    Odrv12 I__3152 (
            .O(N__19492),
            .I(\COUNTER.counterZ0Z_30 ));
    InMux I__3151 (
            .O(N__19487),
            .I(\COUNTER.counter_1_cry_29 ));
    InMux I__3150 (
            .O(N__19484),
            .I(\COUNTER.counter_1_cry_30 ));
    InMux I__3149 (
            .O(N__19481),
            .I(N__19477));
    InMux I__3148 (
            .O(N__19480),
            .I(N__19474));
    LocalMux I__3147 (
            .O(N__19477),
            .I(N__19471));
    LocalMux I__3146 (
            .O(N__19474),
            .I(\COUNTER.counterZ0Z_31 ));
    Odrv12 I__3145 (
            .O(N__19471),
            .I(\COUNTER.counterZ0Z_31 ));
    InMux I__3144 (
            .O(N__19466),
            .I(N__19462));
    InMux I__3143 (
            .O(N__19465),
            .I(N__19459));
    LocalMux I__3142 (
            .O(N__19462),
            .I(\COUNTER.counterZ0Z_14 ));
    LocalMux I__3141 (
            .O(N__19459),
            .I(\COUNTER.counterZ0Z_14 ));
    InMux I__3140 (
            .O(N__19454),
            .I(\COUNTER.counter_1_cry_13 ));
    InMux I__3139 (
            .O(N__19451),
            .I(N__19447));
    InMux I__3138 (
            .O(N__19450),
            .I(N__19444));
    LocalMux I__3137 (
            .O(N__19447),
            .I(\COUNTER.counterZ0Z_15 ));
    LocalMux I__3136 (
            .O(N__19444),
            .I(\COUNTER.counterZ0Z_15 ));
    InMux I__3135 (
            .O(N__19439),
            .I(\COUNTER.counter_1_cry_14 ));
    InMux I__3134 (
            .O(N__19436),
            .I(\COUNTER.counter_1_cry_15 ));
    InMux I__3133 (
            .O(N__19433),
            .I(bfn_6_6_0_));
    InMux I__3132 (
            .O(N__19430),
            .I(\COUNTER.counter_1_cry_17 ));
    InMux I__3131 (
            .O(N__19427),
            .I(\COUNTER.counter_1_cry_18 ));
    InMux I__3130 (
            .O(N__19424),
            .I(\COUNTER.counter_1_cry_19 ));
    InMux I__3129 (
            .O(N__19421),
            .I(\COUNTER.counter_1_cry_20 ));
    InMux I__3128 (
            .O(N__19418),
            .I(\COUNTER.counter_1_cry_21 ));
    CascadeMux I__3127 (
            .O(N__19415),
            .I(N__19411));
    InMux I__3126 (
            .O(N__19414),
            .I(N__19407));
    InMux I__3125 (
            .O(N__19411),
            .I(N__19404));
    InMux I__3124 (
            .O(N__19410),
            .I(N__19401));
    LocalMux I__3123 (
            .O(N__19407),
            .I(\COUNTER.counterZ0Z_6 ));
    LocalMux I__3122 (
            .O(N__19404),
            .I(\COUNTER.counterZ0Z_6 ));
    LocalMux I__3121 (
            .O(N__19401),
            .I(\COUNTER.counterZ0Z_6 ));
    InMux I__3120 (
            .O(N__19394),
            .I(N__19391));
    LocalMux I__3119 (
            .O(N__19391),
            .I(\COUNTER.counter_1_cry_5_THRU_CO ));
    InMux I__3118 (
            .O(N__19388),
            .I(\COUNTER.counter_1_cry_5 ));
    InMux I__3117 (
            .O(N__19385),
            .I(N__19381));
    InMux I__3116 (
            .O(N__19384),
            .I(N__19378));
    LocalMux I__3115 (
            .O(N__19381),
            .I(\COUNTER.counterZ0Z_7 ));
    LocalMux I__3114 (
            .O(N__19378),
            .I(\COUNTER.counterZ0Z_7 ));
    InMux I__3113 (
            .O(N__19373),
            .I(\COUNTER.counter_1_cry_6 ));
    InMux I__3112 (
            .O(N__19370),
            .I(N__19366));
    InMux I__3111 (
            .O(N__19369),
            .I(N__19363));
    LocalMux I__3110 (
            .O(N__19366),
            .I(\COUNTER.counterZ0Z_8 ));
    LocalMux I__3109 (
            .O(N__19363),
            .I(\COUNTER.counterZ0Z_8 ));
    InMux I__3108 (
            .O(N__19358),
            .I(\COUNTER.counter_1_cry_7 ));
    InMux I__3107 (
            .O(N__19355),
            .I(N__19351));
    InMux I__3106 (
            .O(N__19354),
            .I(N__19348));
    LocalMux I__3105 (
            .O(N__19351),
            .I(\COUNTER.counterZ0Z_9 ));
    LocalMux I__3104 (
            .O(N__19348),
            .I(\COUNTER.counterZ0Z_9 ));
    InMux I__3103 (
            .O(N__19343),
            .I(bfn_6_5_0_));
    CascadeMux I__3102 (
            .O(N__19340),
            .I(N__19336));
    InMux I__3101 (
            .O(N__19339),
            .I(N__19333));
    InMux I__3100 (
            .O(N__19336),
            .I(N__19330));
    LocalMux I__3099 (
            .O(N__19333),
            .I(\COUNTER.counterZ0Z_10 ));
    LocalMux I__3098 (
            .O(N__19330),
            .I(\COUNTER.counterZ0Z_10 ));
    InMux I__3097 (
            .O(N__19325),
            .I(\COUNTER.counter_1_cry_9 ));
    InMux I__3096 (
            .O(N__19322),
            .I(N__19318));
    InMux I__3095 (
            .O(N__19321),
            .I(N__19315));
    LocalMux I__3094 (
            .O(N__19318),
            .I(\COUNTER.counterZ0Z_11 ));
    LocalMux I__3093 (
            .O(N__19315),
            .I(\COUNTER.counterZ0Z_11 ));
    InMux I__3092 (
            .O(N__19310),
            .I(\COUNTER.counter_1_cry_10 ));
    CascadeMux I__3091 (
            .O(N__19307),
            .I(N__19303));
    InMux I__3090 (
            .O(N__19306),
            .I(N__19300));
    InMux I__3089 (
            .O(N__19303),
            .I(N__19297));
    LocalMux I__3088 (
            .O(N__19300),
            .I(\COUNTER.counterZ0Z_12 ));
    LocalMux I__3087 (
            .O(N__19297),
            .I(\COUNTER.counterZ0Z_12 ));
    InMux I__3086 (
            .O(N__19292),
            .I(\COUNTER.counter_1_cry_11 ));
    InMux I__3085 (
            .O(N__19289),
            .I(N__19285));
    InMux I__3084 (
            .O(N__19288),
            .I(N__19282));
    LocalMux I__3083 (
            .O(N__19285),
            .I(\COUNTER.counterZ0Z_13 ));
    LocalMux I__3082 (
            .O(N__19282),
            .I(\COUNTER.counterZ0Z_13 ));
    InMux I__3081 (
            .O(N__19277),
            .I(\COUNTER.counter_1_cry_12 ));
    InMux I__3080 (
            .O(N__19274),
            .I(N__19270));
    InMux I__3079 (
            .O(N__19273),
            .I(N__19267));
    LocalMux I__3078 (
            .O(N__19270),
            .I(N__19264));
    LocalMux I__3077 (
            .O(N__19267),
            .I(\HDA_STRAP.countZ0Z_1 ));
    Odrv4 I__3076 (
            .O(N__19264),
            .I(\HDA_STRAP.countZ0Z_1 ));
    InMux I__3075 (
            .O(N__19259),
            .I(N__19255));
    CascadeMux I__3074 (
            .O(N__19258),
            .I(N__19251));
    LocalMux I__3073 (
            .O(N__19255),
            .I(N__19248));
    InMux I__3072 (
            .O(N__19254),
            .I(N__19243));
    InMux I__3071 (
            .O(N__19251),
            .I(N__19243));
    Span4Mux_s0_v I__3070 (
            .O(N__19248),
            .I(N__19240));
    LocalMux I__3069 (
            .O(N__19243),
            .I(\HDA_STRAP.countZ0Z_0 ));
    Odrv4 I__3068 (
            .O(N__19240),
            .I(\HDA_STRAP.countZ0Z_0 ));
    InMux I__3067 (
            .O(N__19235),
            .I(N__19231));
    InMux I__3066 (
            .O(N__19234),
            .I(N__19228));
    LocalMux I__3065 (
            .O(N__19231),
            .I(N__19225));
    LocalMux I__3064 (
            .O(N__19228),
            .I(\HDA_STRAP.countZ0Z_17 ));
    Odrv4 I__3063 (
            .O(N__19225),
            .I(\HDA_STRAP.countZ0Z_17 ));
    InMux I__3062 (
            .O(N__19220),
            .I(N__19217));
    LocalMux I__3061 (
            .O(N__19217),
            .I(\HDA_STRAP.un4_count_9 ));
    InMux I__3060 (
            .O(N__19214),
            .I(N__19202));
    InMux I__3059 (
            .O(N__19213),
            .I(N__19202));
    CascadeMux I__3058 (
            .O(N__19212),
            .I(N__19199));
    InMux I__3057 (
            .O(N__19211),
            .I(N__19186));
    InMux I__3056 (
            .O(N__19210),
            .I(N__19186));
    InMux I__3055 (
            .O(N__19209),
            .I(N__19186));
    InMux I__3054 (
            .O(N__19208),
            .I(N__19186));
    InMux I__3053 (
            .O(N__19207),
            .I(N__19186));
    LocalMux I__3052 (
            .O(N__19202),
            .I(N__19183));
    InMux I__3051 (
            .O(N__19199),
            .I(N__19180));
    InMux I__3050 (
            .O(N__19198),
            .I(N__19175));
    InMux I__3049 (
            .O(N__19197),
            .I(N__19175));
    LocalMux I__3048 (
            .O(N__19186),
            .I(N__19170));
    Span4Mux_v I__3047 (
            .O(N__19183),
            .I(N__19170));
    LocalMux I__3046 (
            .O(N__19180),
            .I(\HDA_STRAP.un4_count ));
    LocalMux I__3045 (
            .O(N__19175),
            .I(\HDA_STRAP.un4_count ));
    Odrv4 I__3044 (
            .O(N__19170),
            .I(\HDA_STRAP.un4_count ));
    CascadeMux I__3043 (
            .O(N__19163),
            .I(N__19157));
    CascadeMux I__3042 (
            .O(N__19162),
            .I(N__19154));
    CascadeMux I__3041 (
            .O(N__19161),
            .I(N__19151));
    CascadeMux I__3040 (
            .O(N__19160),
            .I(N__19147));
    InMux I__3039 (
            .O(N__19157),
            .I(N__19141));
    InMux I__3038 (
            .O(N__19154),
            .I(N__19135));
    InMux I__3037 (
            .O(N__19151),
            .I(N__19135));
    InMux I__3036 (
            .O(N__19150),
            .I(N__19132));
    InMux I__3035 (
            .O(N__19147),
            .I(N__19127));
    InMux I__3034 (
            .O(N__19146),
            .I(N__19127));
    CascadeMux I__3033 (
            .O(N__19145),
            .I(N__19124));
    CascadeMux I__3032 (
            .O(N__19144),
            .I(N__19121));
    LocalMux I__3031 (
            .O(N__19141),
            .I(N__19117));
    InMux I__3030 (
            .O(N__19140),
            .I(N__19114));
    LocalMux I__3029 (
            .O(N__19135),
            .I(N__19111));
    LocalMux I__3028 (
            .O(N__19132),
            .I(N__19106));
    LocalMux I__3027 (
            .O(N__19127),
            .I(N__19106));
    InMux I__3026 (
            .O(N__19124),
            .I(N__19099));
    InMux I__3025 (
            .O(N__19121),
            .I(N__19099));
    InMux I__3024 (
            .O(N__19120),
            .I(N__19099));
    Span4Mux_s1_v I__3023 (
            .O(N__19117),
            .I(N__19096));
    LocalMux I__3022 (
            .O(N__19114),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ));
    Odrv12 I__3021 (
            .O(N__19111),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ));
    Odrv12 I__3020 (
            .O(N__19106),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ));
    LocalMux I__3019 (
            .O(N__19099),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ));
    Odrv4 I__3018 (
            .O(N__19096),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ));
    CascadeMux I__3017 (
            .O(N__19085),
            .I(N__19082));
    InMux I__3016 (
            .O(N__19082),
            .I(N__19079));
    LocalMux I__3015 (
            .O(N__19079),
            .I(\HDA_STRAP.un1_count_1_cry_15_THRU_CO ));
    InMux I__3014 (
            .O(N__19076),
            .I(N__19071));
    InMux I__3013 (
            .O(N__19075),
            .I(N__19066));
    InMux I__3012 (
            .O(N__19074),
            .I(N__19066));
    LocalMux I__3011 (
            .O(N__19071),
            .I(\HDA_STRAP.countZ0Z_16 ));
    LocalMux I__3010 (
            .O(N__19066),
            .I(\HDA_STRAP.countZ0Z_16 ));
    InMux I__3009 (
            .O(N__19061),
            .I(N__19055));
    InMux I__3008 (
            .O(N__19060),
            .I(N__19052));
    InMux I__3007 (
            .O(N__19059),
            .I(N__19047));
    InMux I__3006 (
            .O(N__19058),
            .I(N__19047));
    LocalMux I__3005 (
            .O(N__19055),
            .I(\COUNTER.counterZ0Z_0 ));
    LocalMux I__3004 (
            .O(N__19052),
            .I(\COUNTER.counterZ0Z_0 ));
    LocalMux I__3003 (
            .O(N__19047),
            .I(\COUNTER.counterZ0Z_0 ));
    CascadeMux I__3002 (
            .O(N__19040),
            .I(N__19035));
    CascadeMux I__3001 (
            .O(N__19039),
            .I(N__19032));
    InMux I__3000 (
            .O(N__19038),
            .I(N__19029));
    InMux I__2999 (
            .O(N__19035),
            .I(N__19026));
    InMux I__2998 (
            .O(N__19032),
            .I(N__19023));
    LocalMux I__2997 (
            .O(N__19029),
            .I(\COUNTER.counterZ0Z_1 ));
    LocalMux I__2996 (
            .O(N__19026),
            .I(\COUNTER.counterZ0Z_1 ));
    LocalMux I__2995 (
            .O(N__19023),
            .I(\COUNTER.counterZ0Z_1 ));
    CascadeMux I__2994 (
            .O(N__19016),
            .I(N__19011));
    InMux I__2993 (
            .O(N__19015),
            .I(N__19008));
    InMux I__2992 (
            .O(N__19014),
            .I(N__19003));
    InMux I__2991 (
            .O(N__19011),
            .I(N__19003));
    LocalMux I__2990 (
            .O(N__19008),
            .I(\COUNTER.counterZ0Z_2 ));
    LocalMux I__2989 (
            .O(N__19003),
            .I(\COUNTER.counterZ0Z_2 ));
    InMux I__2988 (
            .O(N__18998),
            .I(N__18995));
    LocalMux I__2987 (
            .O(N__18995),
            .I(N__18992));
    Odrv12 I__2986 (
            .O(N__18992),
            .I(\COUNTER.counter_1_cry_1_THRU_CO ));
    InMux I__2985 (
            .O(N__18989),
            .I(\COUNTER.counter_1_cry_1 ));
    InMux I__2984 (
            .O(N__18986),
            .I(N__18981));
    InMux I__2983 (
            .O(N__18985),
            .I(N__18978));
    InMux I__2982 (
            .O(N__18984),
            .I(N__18975));
    LocalMux I__2981 (
            .O(N__18981),
            .I(\COUNTER.counterZ0Z_3 ));
    LocalMux I__2980 (
            .O(N__18978),
            .I(\COUNTER.counterZ0Z_3 ));
    LocalMux I__2979 (
            .O(N__18975),
            .I(\COUNTER.counterZ0Z_3 ));
    InMux I__2978 (
            .O(N__18968),
            .I(N__18965));
    LocalMux I__2977 (
            .O(N__18965),
            .I(\COUNTER.counter_1_cry_2_THRU_CO ));
    InMux I__2976 (
            .O(N__18962),
            .I(\COUNTER.counter_1_cry_2 ));
    InMux I__2975 (
            .O(N__18959),
            .I(N__18954));
    InMux I__2974 (
            .O(N__18958),
            .I(N__18949));
    InMux I__2973 (
            .O(N__18957),
            .I(N__18949));
    LocalMux I__2972 (
            .O(N__18954),
            .I(\COUNTER.counterZ0Z_4 ));
    LocalMux I__2971 (
            .O(N__18949),
            .I(\COUNTER.counterZ0Z_4 ));
    InMux I__2970 (
            .O(N__18944),
            .I(N__18941));
    LocalMux I__2969 (
            .O(N__18941),
            .I(\COUNTER.counter_1_cry_3_THRU_CO ));
    InMux I__2968 (
            .O(N__18938),
            .I(\COUNTER.counter_1_cry_3 ));
    InMux I__2967 (
            .O(N__18935),
            .I(N__18930));
    InMux I__2966 (
            .O(N__18934),
            .I(N__18925));
    InMux I__2965 (
            .O(N__18933),
            .I(N__18925));
    LocalMux I__2964 (
            .O(N__18930),
            .I(\COUNTER.counterZ0Z_5 ));
    LocalMux I__2963 (
            .O(N__18925),
            .I(\COUNTER.counterZ0Z_5 ));
    InMux I__2962 (
            .O(N__18920),
            .I(N__18917));
    LocalMux I__2961 (
            .O(N__18917),
            .I(\COUNTER.counter_1_cry_4_THRU_CO ));
    InMux I__2960 (
            .O(N__18914),
            .I(\COUNTER.counter_1_cry_4 ));
    InMux I__2959 (
            .O(N__18911),
            .I(N__18906));
    InMux I__2958 (
            .O(N__18910),
            .I(N__18903));
    InMux I__2957 (
            .O(N__18909),
            .I(N__18900));
    LocalMux I__2956 (
            .O(N__18906),
            .I(N__18895));
    LocalMux I__2955 (
            .O(N__18903),
            .I(N__18895));
    LocalMux I__2954 (
            .O(N__18900),
            .I(\HDA_STRAP.countZ0Z_8 ));
    Odrv4 I__2953 (
            .O(N__18895),
            .I(\HDA_STRAP.countZ0Z_8 ));
    InMux I__2952 (
            .O(N__18890),
            .I(N__18886));
    InMux I__2951 (
            .O(N__18889),
            .I(N__18883));
    LocalMux I__2950 (
            .O(N__18886),
            .I(\HDA_STRAP.countZ0Z_14 ));
    LocalMux I__2949 (
            .O(N__18883),
            .I(\HDA_STRAP.countZ0Z_14 ));
    CascadeMux I__2948 (
            .O(N__18878),
            .I(N__18875));
    InMux I__2947 (
            .O(N__18875),
            .I(N__18870));
    InMux I__2946 (
            .O(N__18874),
            .I(N__18867));
    InMux I__2945 (
            .O(N__18873),
            .I(N__18864));
    LocalMux I__2944 (
            .O(N__18870),
            .I(N__18861));
    LocalMux I__2943 (
            .O(N__18867),
            .I(\HDA_STRAP.countZ0Z_6 ));
    LocalMux I__2942 (
            .O(N__18864),
            .I(\HDA_STRAP.countZ0Z_6 ));
    Odrv12 I__2941 (
            .O(N__18861),
            .I(\HDA_STRAP.countZ0Z_6 ));
    InMux I__2940 (
            .O(N__18854),
            .I(N__18850));
    InMux I__2939 (
            .O(N__18853),
            .I(N__18847));
    LocalMux I__2938 (
            .O(N__18850),
            .I(\HDA_STRAP.countZ0Z_15 ));
    LocalMux I__2937 (
            .O(N__18847),
            .I(\HDA_STRAP.countZ0Z_15 ));
    InMux I__2936 (
            .O(N__18842),
            .I(N__18838));
    InMux I__2935 (
            .O(N__18841),
            .I(N__18835));
    LocalMux I__2934 (
            .O(N__18838),
            .I(\HDA_STRAP.countZ0Z_4 ));
    LocalMux I__2933 (
            .O(N__18835),
            .I(\HDA_STRAP.countZ0Z_4 ));
    InMux I__2932 (
            .O(N__18830),
            .I(N__18826));
    InMux I__2931 (
            .O(N__18829),
            .I(N__18823));
    LocalMux I__2930 (
            .O(N__18826),
            .I(\HDA_STRAP.countZ0Z_2 ));
    LocalMux I__2929 (
            .O(N__18823),
            .I(\HDA_STRAP.countZ0Z_2 ));
    CascadeMux I__2928 (
            .O(N__18818),
            .I(N__18815));
    InMux I__2927 (
            .O(N__18815),
            .I(N__18811));
    InMux I__2926 (
            .O(N__18814),
            .I(N__18808));
    LocalMux I__2925 (
            .O(N__18811),
            .I(\HDA_STRAP.countZ0Z_3 ));
    LocalMux I__2924 (
            .O(N__18808),
            .I(\HDA_STRAP.countZ0Z_3 ));
    InMux I__2923 (
            .O(N__18803),
            .I(N__18799));
    InMux I__2922 (
            .O(N__18802),
            .I(N__18796));
    LocalMux I__2921 (
            .O(N__18799),
            .I(\HDA_STRAP.countZ0Z_5 ));
    LocalMux I__2920 (
            .O(N__18796),
            .I(\HDA_STRAP.countZ0Z_5 ));
    InMux I__2919 (
            .O(N__18791),
            .I(N__18787));
    InMux I__2918 (
            .O(N__18790),
            .I(N__18784));
    LocalMux I__2917 (
            .O(N__18787),
            .I(N__18778));
    LocalMux I__2916 (
            .O(N__18784),
            .I(N__18778));
    InMux I__2915 (
            .O(N__18783),
            .I(N__18775));
    Span4Mux_s1_v I__2914 (
            .O(N__18778),
            .I(N__18772));
    LocalMux I__2913 (
            .O(N__18775),
            .I(\HDA_STRAP.countZ0Z_11 ));
    Odrv4 I__2912 (
            .O(N__18772),
            .I(\HDA_STRAP.countZ0Z_11 ));
    InMux I__2911 (
            .O(N__18767),
            .I(N__18762));
    InMux I__2910 (
            .O(N__18766),
            .I(N__18759));
    InMux I__2909 (
            .O(N__18765),
            .I(N__18756));
    LocalMux I__2908 (
            .O(N__18762),
            .I(N__18753));
    LocalMux I__2907 (
            .O(N__18759),
            .I(\HDA_STRAP.countZ0Z_10 ));
    LocalMux I__2906 (
            .O(N__18756),
            .I(\HDA_STRAP.countZ0Z_10 ));
    Odrv4 I__2905 (
            .O(N__18753),
            .I(\HDA_STRAP.countZ0Z_10 ));
    InMux I__2904 (
            .O(N__18746),
            .I(N__18743));
    LocalMux I__2903 (
            .O(N__18743),
            .I(\HDA_STRAP.un4_count_12 ));
    CascadeMux I__2902 (
            .O(N__18740),
            .I(\HDA_STRAP.un4_count_13_cascade_ ));
    InMux I__2901 (
            .O(N__18737),
            .I(N__18734));
    LocalMux I__2900 (
            .O(N__18734),
            .I(\HDA_STRAP.un4_count_10 ));
    InMux I__2899 (
            .O(N__18731),
            .I(N__18727));
    InMux I__2898 (
            .O(N__18730),
            .I(N__18724));
    LocalMux I__2897 (
            .O(N__18727),
            .I(\HDA_STRAP.countZ0Z_9 ));
    LocalMux I__2896 (
            .O(N__18724),
            .I(\HDA_STRAP.countZ0Z_9 ));
    InMux I__2895 (
            .O(N__18719),
            .I(N__18715));
    InMux I__2894 (
            .O(N__18718),
            .I(N__18712));
    LocalMux I__2893 (
            .O(N__18715),
            .I(\HDA_STRAP.countZ0Z_12 ));
    LocalMux I__2892 (
            .O(N__18712),
            .I(\HDA_STRAP.countZ0Z_12 ));
    CascadeMux I__2891 (
            .O(N__18707),
            .I(N__18703));
    InMux I__2890 (
            .O(N__18706),
            .I(N__18700));
    InMux I__2889 (
            .O(N__18703),
            .I(N__18697));
    LocalMux I__2888 (
            .O(N__18700),
            .I(\HDA_STRAP.countZ0Z_13 ));
    LocalMux I__2887 (
            .O(N__18697),
            .I(\HDA_STRAP.countZ0Z_13 ));
    InMux I__2886 (
            .O(N__18692),
            .I(N__18688));
    InMux I__2885 (
            .O(N__18691),
            .I(N__18685));
    LocalMux I__2884 (
            .O(N__18688),
            .I(\HDA_STRAP.countZ0Z_7 ));
    LocalMux I__2883 (
            .O(N__18685),
            .I(\HDA_STRAP.countZ0Z_7 ));
    InMux I__2882 (
            .O(N__18680),
            .I(N__18677));
    LocalMux I__2881 (
            .O(N__18677),
            .I(\HDA_STRAP.un4_count_11 ));
    CascadeMux I__2880 (
            .O(N__18674),
            .I(N__18671));
    InMux I__2879 (
            .O(N__18671),
            .I(N__18668));
    LocalMux I__2878 (
            .O(N__18668),
            .I(\POWERLED.mult1_un89_sum_cry_5_s ));
    InMux I__2877 (
            .O(N__18665),
            .I(\POWERLED.mult1_un89_sum_cry_4 ));
    InMux I__2876 (
            .O(N__18662),
            .I(N__18659));
    LocalMux I__2875 (
            .O(N__18659),
            .I(\POWERLED.mult1_un89_sum_cry_6_s ));
    InMux I__2874 (
            .O(N__18656),
            .I(\POWERLED.mult1_un89_sum_cry_5 ));
    CascadeMux I__2873 (
            .O(N__18653),
            .I(N__18650));
    InMux I__2872 (
            .O(N__18650),
            .I(N__18647));
    LocalMux I__2871 (
            .O(N__18647),
            .I(\POWERLED.mult1_un96_sum_axb_8 ));
    InMux I__2870 (
            .O(N__18644),
            .I(\POWERLED.mult1_un89_sum_cry_6 ));
    InMux I__2869 (
            .O(N__18641),
            .I(\POWERLED.mult1_un89_sum_cry_7 ));
    CascadeMux I__2868 (
            .O(N__18638),
            .I(N__18633));
    InMux I__2867 (
            .O(N__18637),
            .I(N__18629));
    InMux I__2866 (
            .O(N__18636),
            .I(N__18624));
    InMux I__2865 (
            .O(N__18633),
            .I(N__18624));
    InMux I__2864 (
            .O(N__18632),
            .I(N__18621));
    LocalMux I__2863 (
            .O(N__18629),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__2862 (
            .O(N__18624),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__2861 (
            .O(N__18621),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    CascadeMux I__2860 (
            .O(N__18614),
            .I(\POWERLED.mult1_un89_sum_s_8_cascade_ ));
    CascadeMux I__2859 (
            .O(N__18611),
            .I(N__18607));
    CascadeMux I__2858 (
            .O(N__18610),
            .I(N__18603));
    InMux I__2857 (
            .O(N__18607),
            .I(N__18596));
    InMux I__2856 (
            .O(N__18606),
            .I(N__18596));
    InMux I__2855 (
            .O(N__18603),
            .I(N__18596));
    LocalMux I__2854 (
            .O(N__18596),
            .I(\POWERLED.mult1_un89_sum_i_0_8 ));
    CascadeMux I__2853 (
            .O(N__18593),
            .I(N__18590));
    InMux I__2852 (
            .O(N__18590),
            .I(N__18587));
    LocalMux I__2851 (
            .O(N__18587),
            .I(\POWERLED.mult1_un75_sum_i_8 ));
    CascadeMux I__2850 (
            .O(N__18584),
            .I(N__18580));
    CascadeMux I__2849 (
            .O(N__18583),
            .I(N__18576));
    InMux I__2848 (
            .O(N__18580),
            .I(N__18569));
    InMux I__2847 (
            .O(N__18579),
            .I(N__18569));
    InMux I__2846 (
            .O(N__18576),
            .I(N__18569));
    LocalMux I__2845 (
            .O(N__18569),
            .I(\POWERLED.mult1_un82_sum_i_0_8 ));
    InMux I__2844 (
            .O(N__18566),
            .I(N__18563));
    LocalMux I__2843 (
            .O(N__18563),
            .I(N__18560));
    Odrv4 I__2842 (
            .O(N__18560),
            .I(\POWERLED.mult1_un89_sum_i ));
    InMux I__2841 (
            .O(N__18557),
            .I(N__18554));
    LocalMux I__2840 (
            .O(N__18554),
            .I(\POWERLED.mult1_un82_sum_i_8 ));
    InMux I__2839 (
            .O(N__18551),
            .I(\POWERLED.mult1_un96_sum_cry_3 ));
    CascadeMux I__2838 (
            .O(N__18548),
            .I(N__18545));
    InMux I__2837 (
            .O(N__18545),
            .I(N__18542));
    LocalMux I__2836 (
            .O(N__18542),
            .I(\POWERLED.mult1_un96_sum_cry_5_s ));
    InMux I__2835 (
            .O(N__18539),
            .I(\POWERLED.mult1_un96_sum_cry_4 ));
    InMux I__2834 (
            .O(N__18536),
            .I(N__18533));
    LocalMux I__2833 (
            .O(N__18533),
            .I(\POWERLED.mult1_un96_sum_cry_6_s ));
    InMux I__2832 (
            .O(N__18530),
            .I(\POWERLED.mult1_un96_sum_cry_5 ));
    CascadeMux I__2831 (
            .O(N__18527),
            .I(N__18524));
    InMux I__2830 (
            .O(N__18524),
            .I(N__18521));
    LocalMux I__2829 (
            .O(N__18521),
            .I(\POWERLED.mult1_un103_sum_axb_8 ));
    InMux I__2828 (
            .O(N__18518),
            .I(\POWERLED.mult1_un96_sum_cry_6 ));
    InMux I__2827 (
            .O(N__18515),
            .I(\POWERLED.mult1_un96_sum_cry_7 ));
    InMux I__2826 (
            .O(N__18512),
            .I(N__18509));
    LocalMux I__2825 (
            .O(N__18509),
            .I(N__18505));
    CascadeMux I__2824 (
            .O(N__18508),
            .I(N__18501));
    Span4Mux_h I__2823 (
            .O(N__18505),
            .I(N__18496));
    InMux I__2822 (
            .O(N__18504),
            .I(N__18491));
    InMux I__2821 (
            .O(N__18501),
            .I(N__18491));
    InMux I__2820 (
            .O(N__18500),
            .I(N__18488));
    InMux I__2819 (
            .O(N__18499),
            .I(N__18485));
    Odrv4 I__2818 (
            .O(N__18496),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__2817 (
            .O(N__18491),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__2816 (
            .O(N__18488),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__2815 (
            .O(N__18485),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    InMux I__2814 (
            .O(N__18476),
            .I(N__18473));
    LocalMux I__2813 (
            .O(N__18473),
            .I(\POWERLED.mult1_un131_sum_i_8 ));
    CascadeMux I__2812 (
            .O(N__18470),
            .I(N__18467));
    InMux I__2811 (
            .O(N__18467),
            .I(N__18464));
    LocalMux I__2810 (
            .O(N__18464),
            .I(\POWERLED.mult1_un89_sum_cry_3_s ));
    InMux I__2809 (
            .O(N__18461),
            .I(\POWERLED.mult1_un89_sum_cry_2 ));
    InMux I__2808 (
            .O(N__18458),
            .I(N__18455));
    LocalMux I__2807 (
            .O(N__18455),
            .I(\POWERLED.mult1_un89_sum_cry_4_s ));
    InMux I__2806 (
            .O(N__18452),
            .I(\POWERLED.mult1_un89_sum_cry_3 ));
    InMux I__2805 (
            .O(N__18449),
            .I(N__18446));
    LocalMux I__2804 (
            .O(N__18446),
            .I(\POWERLED.mult1_un138_sum_i_8 ));
    InMux I__2803 (
            .O(N__18443),
            .I(N__18440));
    LocalMux I__2802 (
            .O(N__18440),
            .I(\POWERLED.un85_clk_100khz_1 ));
    InMux I__2801 (
            .O(N__18437),
            .I(N__18434));
    LocalMux I__2800 (
            .O(N__18434),
            .I(N__18431));
    Odrv4 I__2799 (
            .O(N__18431),
            .I(\POWERLED.mult1_un96_sum_i ));
    CascadeMux I__2798 (
            .O(N__18428),
            .I(N__18424));
    CascadeMux I__2797 (
            .O(N__18427),
            .I(N__18420));
    InMux I__2796 (
            .O(N__18424),
            .I(N__18413));
    InMux I__2795 (
            .O(N__18423),
            .I(N__18413));
    InMux I__2794 (
            .O(N__18420),
            .I(N__18413));
    LocalMux I__2793 (
            .O(N__18413),
            .I(\POWERLED.mult1_un96_sum_i_0_8 ));
    CascadeMux I__2792 (
            .O(N__18410),
            .I(N__18405));
    InMux I__2791 (
            .O(N__18409),
            .I(N__18401));
    InMux I__2790 (
            .O(N__18408),
            .I(N__18396));
    InMux I__2789 (
            .O(N__18405),
            .I(N__18396));
    InMux I__2788 (
            .O(N__18404),
            .I(N__18393));
    LocalMux I__2787 (
            .O(N__18401),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__2786 (
            .O(N__18396),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__2785 (
            .O(N__18393),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    CascadeMux I__2784 (
            .O(N__18386),
            .I(N__18383));
    InMux I__2783 (
            .O(N__18383),
            .I(N__18380));
    LocalMux I__2782 (
            .O(N__18380),
            .I(N__18377));
    Odrv4 I__2781 (
            .O(N__18377),
            .I(\POWERLED.mult1_un103_sum_i_8 ));
    InMux I__2780 (
            .O(N__18374),
            .I(N__18368));
    CascadeMux I__2779 (
            .O(N__18373),
            .I(N__18365));
    CascadeMux I__2778 (
            .O(N__18372),
            .I(N__18362));
    InMux I__2777 (
            .O(N__18371),
            .I(N__18358));
    LocalMux I__2776 (
            .O(N__18368),
            .I(N__18355));
    InMux I__2775 (
            .O(N__18365),
            .I(N__18352));
    InMux I__2774 (
            .O(N__18362),
            .I(N__18347));
    InMux I__2773 (
            .O(N__18361),
            .I(N__18347));
    LocalMux I__2772 (
            .O(N__18358),
            .I(N__18344));
    Odrv4 I__2771 (
            .O(N__18355),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__2770 (
            .O(N__18352),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__2769 (
            .O(N__18347),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    Odrv4 I__2768 (
            .O(N__18344),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    InMux I__2767 (
            .O(N__18335),
            .I(N__18332));
    LocalMux I__2766 (
            .O(N__18332),
            .I(\POWERLED.mult1_un124_sum_i_8 ));
    CascadeMux I__2765 (
            .O(N__18329),
            .I(N__18326));
    InMux I__2764 (
            .O(N__18326),
            .I(N__18323));
    LocalMux I__2763 (
            .O(N__18323),
            .I(\POWERLED.mult1_un96_sum_cry_3_s ));
    InMux I__2762 (
            .O(N__18320),
            .I(\POWERLED.mult1_un96_sum_cry_2 ));
    InMux I__2761 (
            .O(N__18317),
            .I(N__18314));
    LocalMux I__2760 (
            .O(N__18314),
            .I(\POWERLED.mult1_un96_sum_cry_4_s ));
    CascadeMux I__2759 (
            .O(N__18311),
            .I(N__18307));
    CascadeMux I__2758 (
            .O(N__18310),
            .I(N__18303));
    InMux I__2757 (
            .O(N__18307),
            .I(N__18296));
    InMux I__2756 (
            .O(N__18306),
            .I(N__18296));
    InMux I__2755 (
            .O(N__18303),
            .I(N__18296));
    LocalMux I__2754 (
            .O(N__18296),
            .I(G_2150));
    InMux I__2753 (
            .O(N__18293),
            .I(\POWERLED.mult1_un166_sum_cry_5 ));
    InMux I__2752 (
            .O(N__18290),
            .I(N__18287));
    LocalMux I__2751 (
            .O(N__18287),
            .I(N__18284));
    Odrv4 I__2750 (
            .O(N__18284),
            .I(\POWERLED.un85_clk_100khz_0 ));
    InMux I__2749 (
            .O(N__18281),
            .I(N__18278));
    LocalMux I__2748 (
            .O(N__18278),
            .I(N__18275));
    Odrv4 I__2747 (
            .O(N__18275),
            .I(\POWERLED.un85_clk_100khz_2 ));
    InMux I__2746 (
            .O(N__18272),
            .I(N__18269));
    LocalMux I__2745 (
            .O(N__18269),
            .I(\POWERLED.un85_clk_100khz_3 ));
    InMux I__2744 (
            .O(N__18266),
            .I(\POWERLED.mult1_un131_sum_cry_7 ));
    CascadeMux I__2743 (
            .O(N__18263),
            .I(N__18258));
    CascadeMux I__2742 (
            .O(N__18262),
            .I(N__18255));
    CascadeMux I__2741 (
            .O(N__18261),
            .I(N__18252));
    InMux I__2740 (
            .O(N__18258),
            .I(N__18249));
    InMux I__2739 (
            .O(N__18255),
            .I(N__18244));
    InMux I__2738 (
            .O(N__18252),
            .I(N__18244));
    LocalMux I__2737 (
            .O(N__18249),
            .I(\POWERLED.mult1_un124_sum_i_0_8 ));
    LocalMux I__2736 (
            .O(N__18244),
            .I(\POWERLED.mult1_un124_sum_i_0_8 ));
    InMux I__2735 (
            .O(N__18239),
            .I(\POWERLED.mult1_un145_sum_cry_2_c ));
    InMux I__2734 (
            .O(N__18236),
            .I(\POWERLED.mult1_un145_sum_cry_3_c ));
    InMux I__2733 (
            .O(N__18233),
            .I(\POWERLED.mult1_un145_sum_cry_4_c ));
    InMux I__2732 (
            .O(N__18230),
            .I(\POWERLED.mult1_un145_sum_cry_5_c ));
    InMux I__2731 (
            .O(N__18227),
            .I(\POWERLED.mult1_un145_sum_cry_6_c ));
    InMux I__2730 (
            .O(N__18224),
            .I(\POWERLED.mult1_un145_sum_cry_7 ));
    CascadeMux I__2729 (
            .O(N__18221),
            .I(\POWERLED.mult1_un145_sum_s_8_cascade_ ));
    InMux I__2728 (
            .O(N__18218),
            .I(N__18214));
    InMux I__2727 (
            .O(N__18217),
            .I(N__18211));
    LocalMux I__2726 (
            .O(N__18214),
            .I(\VPP_VDDQ.count_2Z0Z_15 ));
    LocalMux I__2725 (
            .O(N__18211),
            .I(\VPP_VDDQ.count_2Z0Z_15 ));
    InMux I__2724 (
            .O(N__18206),
            .I(N__18186));
    InMux I__2723 (
            .O(N__18205),
            .I(N__18186));
    InMux I__2722 (
            .O(N__18204),
            .I(N__18186));
    InMux I__2721 (
            .O(N__18203),
            .I(N__18179));
    InMux I__2720 (
            .O(N__18202),
            .I(N__18179));
    InMux I__2719 (
            .O(N__18201),
            .I(N__18179));
    InMux I__2718 (
            .O(N__18200),
            .I(N__18170));
    InMux I__2717 (
            .O(N__18199),
            .I(N__18170));
    InMux I__2716 (
            .O(N__18198),
            .I(N__18170));
    InMux I__2715 (
            .O(N__18197),
            .I(N__18170));
    InMux I__2714 (
            .O(N__18196),
            .I(N__18161));
    InMux I__2713 (
            .O(N__18195),
            .I(N__18161));
    InMux I__2712 (
            .O(N__18194),
            .I(N__18161));
    InMux I__2711 (
            .O(N__18193),
            .I(N__18161));
    LocalMux I__2710 (
            .O(N__18186),
            .I(N__18155));
    LocalMux I__2709 (
            .O(N__18179),
            .I(N__18155));
    LocalMux I__2708 (
            .O(N__18170),
            .I(N__18150));
    LocalMux I__2707 (
            .O(N__18161),
            .I(N__18150));
    CascadeMux I__2706 (
            .O(N__18160),
            .I(N__18146));
    Span4Mux_v I__2705 (
            .O(N__18155),
            .I(N__18142));
    Span4Mux_v I__2704 (
            .O(N__18150),
            .I(N__18139));
    InMux I__2703 (
            .O(N__18149),
            .I(N__18132));
    InMux I__2702 (
            .O(N__18146),
            .I(N__18132));
    InMux I__2701 (
            .O(N__18145),
            .I(N__18132));
    Odrv4 I__2700 (
            .O(N__18142),
            .I(\VPP_VDDQ.count_2_1_sqmuxa ));
    Odrv4 I__2699 (
            .O(N__18139),
            .I(\VPP_VDDQ.count_2_1_sqmuxa ));
    LocalMux I__2698 (
            .O(N__18132),
            .I(\VPP_VDDQ.count_2_1_sqmuxa ));
    InMux I__2697 (
            .O(N__18125),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14 ));
    InMux I__2696 (
            .O(N__18122),
            .I(N__18118));
    InMux I__2695 (
            .O(N__18121),
            .I(N__18115));
    LocalMux I__2694 (
            .O(N__18118),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ));
    LocalMux I__2693 (
            .O(N__18115),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ));
    InMux I__2692 (
            .O(N__18110),
            .I(N__18107));
    LocalMux I__2691 (
            .O(N__18107),
            .I(\VPP_VDDQ.count_2_0_15 ));
    InMux I__2690 (
            .O(N__18104),
            .I(\POWERLED.mult1_un131_sum_cry_2 ));
    InMux I__2689 (
            .O(N__18101),
            .I(N__18098));
    LocalMux I__2688 (
            .O(N__18098),
            .I(\POWERLED.mult1_un124_sum_cry_3_s ));
    InMux I__2687 (
            .O(N__18095),
            .I(\POWERLED.mult1_un131_sum_cry_3 ));
    InMux I__2686 (
            .O(N__18092),
            .I(N__18089));
    LocalMux I__2685 (
            .O(N__18089),
            .I(\POWERLED.mult1_un124_sum_cry_4_s ));
    InMux I__2684 (
            .O(N__18086),
            .I(\POWERLED.mult1_un131_sum_cry_4 ));
    InMux I__2683 (
            .O(N__18083),
            .I(N__18080));
    LocalMux I__2682 (
            .O(N__18080),
            .I(\POWERLED.mult1_un124_sum_cry_5_s ));
    InMux I__2681 (
            .O(N__18077),
            .I(\POWERLED.mult1_un131_sum_cry_5 ));
    InMux I__2680 (
            .O(N__18074),
            .I(N__18071));
    LocalMux I__2679 (
            .O(N__18071),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    InMux I__2678 (
            .O(N__18068),
            .I(\POWERLED.mult1_un131_sum_cry_6 ));
    InMux I__2677 (
            .O(N__18065),
            .I(N__18062));
    LocalMux I__2676 (
            .O(N__18062),
            .I(\POWERLED.mult1_un131_sum_axb_8 ));
    InMux I__2675 (
            .O(N__18059),
            .I(N__18056));
    LocalMux I__2674 (
            .O(N__18056),
            .I(N__18053));
    Odrv4 I__2673 (
            .O(N__18053),
            .I(\VPP_VDDQ.un1_count_2_1_axb_7 ));
    InMux I__2672 (
            .O(N__18050),
            .I(N__18044));
    InMux I__2671 (
            .O(N__18049),
            .I(N__18044));
    LocalMux I__2670 (
            .O(N__18044),
            .I(N__18040));
    InMux I__2669 (
            .O(N__18043),
            .I(N__18037));
    Odrv4 I__2668 (
            .O(N__18040),
            .I(\VPP_VDDQ.count_2_1_7 ));
    LocalMux I__2667 (
            .O(N__18037),
            .I(\VPP_VDDQ.count_2_1_7 ));
    InMux I__2666 (
            .O(N__18032),
            .I(\VPP_VDDQ.un1_count_2_1_cry_6 ));
    InMux I__2665 (
            .O(N__18029),
            .I(N__18025));
    InMux I__2664 (
            .O(N__18028),
            .I(N__18022));
    LocalMux I__2663 (
            .O(N__18025),
            .I(\VPP_VDDQ.count_2_1_8 ));
    LocalMux I__2662 (
            .O(N__18022),
            .I(\VPP_VDDQ.count_2_1_8 ));
    InMux I__2661 (
            .O(N__18017),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7 ));
    InMux I__2660 (
            .O(N__18014),
            .I(N__18011));
    LocalMux I__2659 (
            .O(N__18011),
            .I(N__18008));
    Odrv4 I__2658 (
            .O(N__18008),
            .I(\VPP_VDDQ.count_2Z0Z_9 ));
    InMux I__2657 (
            .O(N__18005),
            .I(N__17999));
    InMux I__2656 (
            .O(N__18004),
            .I(N__17999));
    LocalMux I__2655 (
            .O(N__17999),
            .I(N__17996));
    Odrv4 I__2654 (
            .O(N__17996),
            .I(\VPP_VDDQ.count_2_1_9 ));
    InMux I__2653 (
            .O(N__17993),
            .I(bfn_5_9_0_));
    InMux I__2652 (
            .O(N__17990),
            .I(N__17987));
    LocalMux I__2651 (
            .O(N__17987),
            .I(N__17983));
    InMux I__2650 (
            .O(N__17986),
            .I(N__17980));
    Odrv4 I__2649 (
            .O(N__17983),
            .I(\VPP_VDDQ.count_2Z0Z_10 ));
    LocalMux I__2648 (
            .O(N__17980),
            .I(\VPP_VDDQ.count_2Z0Z_10 ));
    InMux I__2647 (
            .O(N__17975),
            .I(N__17971));
    InMux I__2646 (
            .O(N__17974),
            .I(N__17968));
    LocalMux I__2645 (
            .O(N__17971),
            .I(N__17965));
    LocalMux I__2644 (
            .O(N__17968),
            .I(\VPP_VDDQ.count_2_1_10 ));
    Odrv4 I__2643 (
            .O(N__17965),
            .I(\VPP_VDDQ.count_2_1_10 ));
    InMux I__2642 (
            .O(N__17960),
            .I(\VPP_VDDQ.un1_count_2_1_cry_9 ));
    InMux I__2641 (
            .O(N__17957),
            .I(N__17953));
    CascadeMux I__2640 (
            .O(N__17956),
            .I(N__17950));
    LocalMux I__2639 (
            .O(N__17953),
            .I(N__17947));
    InMux I__2638 (
            .O(N__17950),
            .I(N__17944));
    Odrv4 I__2637 (
            .O(N__17947),
            .I(\VPP_VDDQ.count_2Z0Z_11 ));
    LocalMux I__2636 (
            .O(N__17944),
            .I(\VPP_VDDQ.count_2Z0Z_11 ));
    InMux I__2635 (
            .O(N__17939),
            .I(N__17933));
    InMux I__2634 (
            .O(N__17938),
            .I(N__17933));
    LocalMux I__2633 (
            .O(N__17933),
            .I(N__17930));
    Odrv4 I__2632 (
            .O(N__17930),
            .I(\VPP_VDDQ.count_2_1_11 ));
    InMux I__2631 (
            .O(N__17927),
            .I(\VPP_VDDQ.un1_count_2_1_cry_10 ));
    InMux I__2630 (
            .O(N__17924),
            .I(N__17920));
    InMux I__2629 (
            .O(N__17923),
            .I(N__17917));
    LocalMux I__2628 (
            .O(N__17920),
            .I(\VPP_VDDQ.count_2Z0Z_12 ));
    LocalMux I__2627 (
            .O(N__17917),
            .I(\VPP_VDDQ.count_2Z0Z_12 ));
    InMux I__2626 (
            .O(N__17912),
            .I(N__17906));
    InMux I__2625 (
            .O(N__17911),
            .I(N__17906));
    LocalMux I__2624 (
            .O(N__17906),
            .I(\VPP_VDDQ.count_2_1_12 ));
    InMux I__2623 (
            .O(N__17903),
            .I(\VPP_VDDQ.un1_count_2_1_cry_11 ));
    CascadeMux I__2622 (
            .O(N__17900),
            .I(N__17896));
    InMux I__2621 (
            .O(N__17899),
            .I(N__17893));
    InMux I__2620 (
            .O(N__17896),
            .I(N__17890));
    LocalMux I__2619 (
            .O(N__17893),
            .I(\VPP_VDDQ.count_2Z0Z_13 ));
    LocalMux I__2618 (
            .O(N__17890),
            .I(\VPP_VDDQ.count_2Z0Z_13 ));
    InMux I__2617 (
            .O(N__17885),
            .I(N__17879));
    InMux I__2616 (
            .O(N__17884),
            .I(N__17879));
    LocalMux I__2615 (
            .O(N__17879),
            .I(\VPP_VDDQ.count_2_1_13 ));
    InMux I__2614 (
            .O(N__17876),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12 ));
    InMux I__2613 (
            .O(N__17873),
            .I(N__17869));
    InMux I__2612 (
            .O(N__17872),
            .I(N__17866));
    LocalMux I__2611 (
            .O(N__17869),
            .I(\VPP_VDDQ.count_2Z0Z_14 ));
    LocalMux I__2610 (
            .O(N__17866),
            .I(\VPP_VDDQ.count_2Z0Z_14 ));
    InMux I__2609 (
            .O(N__17861),
            .I(N__17855));
    InMux I__2608 (
            .O(N__17860),
            .I(N__17855));
    LocalMux I__2607 (
            .O(N__17855),
            .I(\VPP_VDDQ.count_2_1_14 ));
    InMux I__2606 (
            .O(N__17852),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13 ));
    InMux I__2605 (
            .O(N__17849),
            .I(N__17846));
    LocalMux I__2604 (
            .O(N__17846),
            .I(N__17843));
    Odrv4 I__2603 (
            .O(N__17843),
            .I(\VPP_VDDQ.count_2_0_5 ));
    InMux I__2602 (
            .O(N__17840),
            .I(N__17837));
    LocalMux I__2601 (
            .O(N__17837),
            .I(N__17834));
    Odrv4 I__2600 (
            .O(N__17834),
            .I(\VPP_VDDQ.count_2_0_8 ));
    InMux I__2599 (
            .O(N__17831),
            .I(N__17828));
    LocalMux I__2598 (
            .O(N__17828),
            .I(N__17825));
    Odrv4 I__2597 (
            .O(N__17825),
            .I(\VPP_VDDQ.count_2_0_10 ));
    InMux I__2596 (
            .O(N__17822),
            .I(N__17817));
    InMux I__2595 (
            .O(N__17821),
            .I(N__17810));
    InMux I__2594 (
            .O(N__17820),
            .I(N__17810));
    LocalMux I__2593 (
            .O(N__17817),
            .I(N__17807));
    InMux I__2592 (
            .O(N__17816),
            .I(N__17802));
    InMux I__2591 (
            .O(N__17815),
            .I(N__17802));
    LocalMux I__2590 (
            .O(N__17810),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    Odrv4 I__2589 (
            .O(N__17807),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    LocalMux I__2588 (
            .O(N__17802),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    CascadeMux I__2587 (
            .O(N__17795),
            .I(N__17792));
    InMux I__2586 (
            .O(N__17792),
            .I(N__17789));
    LocalMux I__2585 (
            .O(N__17789),
            .I(N__17784));
    InMux I__2584 (
            .O(N__17788),
            .I(N__17779));
    InMux I__2583 (
            .O(N__17787),
            .I(N__17779));
    Span4Mux_v I__2582 (
            .O(N__17784),
            .I(N__17776));
    LocalMux I__2581 (
            .O(N__17779),
            .I(\VPP_VDDQ.un1_count_2_1_axb_1 ));
    Odrv4 I__2580 (
            .O(N__17776),
            .I(\VPP_VDDQ.un1_count_2_1_axb_1 ));
    InMux I__2579 (
            .O(N__17771),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1 ));
    InMux I__2578 (
            .O(N__17768),
            .I(N__17764));
    InMux I__2577 (
            .O(N__17767),
            .I(N__17761));
    LocalMux I__2576 (
            .O(N__17764),
            .I(\VPP_VDDQ.count_2_1_3 ));
    LocalMux I__2575 (
            .O(N__17761),
            .I(\VPP_VDDQ.count_2_1_3 ));
    InMux I__2574 (
            .O(N__17756),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2 ));
    InMux I__2573 (
            .O(N__17753),
            .I(\VPP_VDDQ.un1_count_2_1_cry_3 ));
    InMux I__2572 (
            .O(N__17750),
            .I(N__17746));
    InMux I__2571 (
            .O(N__17749),
            .I(N__17743));
    LocalMux I__2570 (
            .O(N__17746),
            .I(\VPP_VDDQ.count_2_1_5 ));
    LocalMux I__2569 (
            .O(N__17743),
            .I(\VPP_VDDQ.count_2_1_5 ));
    InMux I__2568 (
            .O(N__17738),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4 ));
    InMux I__2567 (
            .O(N__17735),
            .I(\VPP_VDDQ.un1_count_2_1_cry_5 ));
    CEMux I__2566 (
            .O(N__17732),
            .I(N__17729));
    LocalMux I__2565 (
            .O(N__17729),
            .I(N__17726));
    Span4Mux_h I__2564 (
            .O(N__17726),
            .I(N__17723));
    Odrv4 I__2563 (
            .O(N__17723),
            .I(\RSMRST_PWRGD.N_92_1 ));
    InMux I__2562 (
            .O(N__17720),
            .I(N__17717));
    LocalMux I__2561 (
            .O(N__17717),
            .I(N__17714));
    Odrv4 I__2560 (
            .O(N__17714),
            .I(\VPP_VDDQ.count_2_0_3 ));
    InMux I__2559 (
            .O(N__17711),
            .I(\HDA_STRAP.un1_count_1_cry_13 ));
    InMux I__2558 (
            .O(N__17708),
            .I(\HDA_STRAP.un1_count_1_cry_14 ));
    InMux I__2557 (
            .O(N__17705),
            .I(bfn_5_3_0_));
    InMux I__2556 (
            .O(N__17702),
            .I(\HDA_STRAP.un1_count_1_cry_16 ));
    InMux I__2555 (
            .O(N__17699),
            .I(\HDA_STRAP.un1_count_1_cry_4 ));
    InMux I__2554 (
            .O(N__17696),
            .I(N__17693));
    LocalMux I__2553 (
            .O(N__17693),
            .I(\HDA_STRAP.un1_count_1_cry_5_THRU_CO ));
    InMux I__2552 (
            .O(N__17690),
            .I(\HDA_STRAP.un1_count_1_cry_5 ));
    InMux I__2551 (
            .O(N__17687),
            .I(\HDA_STRAP.un1_count_1_cry_6 ));
    InMux I__2550 (
            .O(N__17684),
            .I(N__17681));
    LocalMux I__2549 (
            .O(N__17681),
            .I(\HDA_STRAP.un1_count_1_cry_7_THRU_CO ));
    InMux I__2548 (
            .O(N__17678),
            .I(bfn_5_2_0_));
    InMux I__2547 (
            .O(N__17675),
            .I(\HDA_STRAP.un1_count_1_cry_8 ));
    InMux I__2546 (
            .O(N__17672),
            .I(N__17669));
    LocalMux I__2545 (
            .O(N__17669),
            .I(\HDA_STRAP.un1_count_1_cry_9_THRU_CO ));
    InMux I__2544 (
            .O(N__17666),
            .I(\HDA_STRAP.un1_count_1_cry_9 ));
    InMux I__2543 (
            .O(N__17663),
            .I(N__17660));
    LocalMux I__2542 (
            .O(N__17660),
            .I(\HDA_STRAP.un1_count_1_cry_10_THRU_CO ));
    InMux I__2541 (
            .O(N__17657),
            .I(\HDA_STRAP.un1_count_1_cry_10 ));
    InMux I__2540 (
            .O(N__17654),
            .I(\HDA_STRAP.un1_count_1_cry_11 ));
    InMux I__2539 (
            .O(N__17651),
            .I(\HDA_STRAP.un1_count_1_cry_12 ));
    InMux I__2538 (
            .O(N__17648),
            .I(N__17645));
    LocalMux I__2537 (
            .O(N__17645),
            .I(N__17641));
    CascadeMux I__2536 (
            .O(N__17644),
            .I(N__17637));
    Span4Mux_v I__2535 (
            .O(N__17641),
            .I(N__17634));
    InMux I__2534 (
            .O(N__17640),
            .I(N__17631));
    InMux I__2533 (
            .O(N__17637),
            .I(N__17628));
    Odrv4 I__2532 (
            .O(N__17634),
            .I(\POWERLED.countZ0Z_15 ));
    LocalMux I__2531 (
            .O(N__17631),
            .I(\POWERLED.countZ0Z_15 ));
    LocalMux I__2530 (
            .O(N__17628),
            .I(\POWERLED.countZ0Z_15 ));
    CascadeMux I__2529 (
            .O(N__17621),
            .I(N__17618));
    InMux I__2528 (
            .O(N__17618),
            .I(N__17615));
    LocalMux I__2527 (
            .O(N__17615),
            .I(\POWERLED.N_5050_i ));
    InMux I__2526 (
            .O(N__17612),
            .I(bfn_4_16_0_));
    InMux I__2525 (
            .O(N__17609),
            .I(N__17604));
    InMux I__2524 (
            .O(N__17608),
            .I(N__17598));
    InMux I__2523 (
            .O(N__17607),
            .I(N__17598));
    LocalMux I__2522 (
            .O(N__17604),
            .I(N__17595));
    InMux I__2521 (
            .O(N__17603),
            .I(N__17592));
    LocalMux I__2520 (
            .O(N__17598),
            .I(N__17589));
    Span4Mux_v I__2519 (
            .O(N__17595),
            .I(N__17586));
    LocalMux I__2518 (
            .O(N__17592),
            .I(N__17583));
    Span4Mux_s3_h I__2517 (
            .O(N__17589),
            .I(N__17580));
    Odrv4 I__2516 (
            .O(N__17586),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    Odrv12 I__2515 (
            .O(N__17583),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    Odrv4 I__2514 (
            .O(N__17580),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    InMux I__2513 (
            .O(N__17573),
            .I(N__17570));
    LocalMux I__2512 (
            .O(N__17570),
            .I(\POWERLED.mult1_un89_sum_i_8 ));
    CascadeMux I__2511 (
            .O(N__17567),
            .I(N__17564));
    InMux I__2510 (
            .O(N__17564),
            .I(N__17561));
    LocalMux I__2509 (
            .O(N__17561),
            .I(\POWERLED.mult1_un68_sum_i_8 ));
    InMux I__2508 (
            .O(N__17558),
            .I(\HDA_STRAP.un1_count_1_cry_0 ));
    InMux I__2507 (
            .O(N__17555),
            .I(\HDA_STRAP.un1_count_1_cry_1 ));
    InMux I__2506 (
            .O(N__17552),
            .I(\HDA_STRAP.un1_count_1_cry_2 ));
    InMux I__2505 (
            .O(N__17549),
            .I(\HDA_STRAP.un1_count_1_cry_3 ));
    CascadeMux I__2504 (
            .O(N__17546),
            .I(N__17543));
    InMux I__2503 (
            .O(N__17543),
            .I(N__17540));
    LocalMux I__2502 (
            .O(N__17540),
            .I(N__17537));
    Odrv4 I__2501 (
            .O(N__17537),
            .I(\POWERLED.mult1_un110_sum_i_8 ));
    InMux I__2500 (
            .O(N__17534),
            .I(N__17531));
    LocalMux I__2499 (
            .O(N__17531),
            .I(N__17527));
    CascadeMux I__2498 (
            .O(N__17530),
            .I(N__17523));
    Span4Mux_v I__2497 (
            .O(N__17527),
            .I(N__17520));
    InMux I__2496 (
            .O(N__17526),
            .I(N__17517));
    InMux I__2495 (
            .O(N__17523),
            .I(N__17514));
    Odrv4 I__2494 (
            .O(N__17520),
            .I(\POWERLED.countZ0Z_8 ));
    LocalMux I__2493 (
            .O(N__17517),
            .I(\POWERLED.countZ0Z_8 ));
    LocalMux I__2492 (
            .O(N__17514),
            .I(\POWERLED.countZ0Z_8 ));
    InMux I__2491 (
            .O(N__17507),
            .I(N__17504));
    LocalMux I__2490 (
            .O(N__17504),
            .I(\POWERLED.N_5043_i ));
    InMux I__2489 (
            .O(N__17501),
            .I(N__17498));
    LocalMux I__2488 (
            .O(N__17498),
            .I(N__17494));
    CascadeMux I__2487 (
            .O(N__17497),
            .I(N__17490));
    Span4Mux_v I__2486 (
            .O(N__17494),
            .I(N__17487));
    InMux I__2485 (
            .O(N__17493),
            .I(N__17484));
    InMux I__2484 (
            .O(N__17490),
            .I(N__17481));
    Odrv4 I__2483 (
            .O(N__17487),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__2482 (
            .O(N__17484),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__2481 (
            .O(N__17481),
            .I(\POWERLED.countZ0Z_9 ));
    InMux I__2480 (
            .O(N__17474),
            .I(N__17471));
    LocalMux I__2479 (
            .O(N__17471),
            .I(\POWERLED.N_5044_i ));
    InMux I__2478 (
            .O(N__17468),
            .I(N__17465));
    LocalMux I__2477 (
            .O(N__17465),
            .I(N__17461));
    CascadeMux I__2476 (
            .O(N__17464),
            .I(N__17458));
    Span4Mux_s3_v I__2475 (
            .O(N__17461),
            .I(N__17455));
    InMux I__2474 (
            .O(N__17458),
            .I(N__17451));
    Span4Mux_v I__2473 (
            .O(N__17455),
            .I(N__17448));
    InMux I__2472 (
            .O(N__17454),
            .I(N__17445));
    LocalMux I__2471 (
            .O(N__17451),
            .I(N__17442));
    Odrv4 I__2470 (
            .O(N__17448),
            .I(\POWERLED.countZ0Z_10 ));
    LocalMux I__2469 (
            .O(N__17445),
            .I(\POWERLED.countZ0Z_10 ));
    Odrv4 I__2468 (
            .O(N__17442),
            .I(\POWERLED.countZ0Z_10 ));
    CascadeMux I__2467 (
            .O(N__17435),
            .I(N__17432));
    InMux I__2466 (
            .O(N__17432),
            .I(N__17429));
    LocalMux I__2465 (
            .O(N__17429),
            .I(N__17426));
    Span4Mux_h I__2464 (
            .O(N__17426),
            .I(N__17423));
    Odrv4 I__2463 (
            .O(N__17423),
            .I(\POWERLED.mult1_un96_sum_i_8 ));
    InMux I__2462 (
            .O(N__17420),
            .I(N__17417));
    LocalMux I__2461 (
            .O(N__17417),
            .I(\POWERLED.N_5045_i ));
    InMux I__2460 (
            .O(N__17414),
            .I(N__17411));
    LocalMux I__2459 (
            .O(N__17411),
            .I(N__17407));
    CascadeMux I__2458 (
            .O(N__17410),
            .I(N__17404));
    Span4Mux_v I__2457 (
            .O(N__17407),
            .I(N__17400));
    InMux I__2456 (
            .O(N__17404),
            .I(N__17397));
    InMux I__2455 (
            .O(N__17403),
            .I(N__17394));
    Span4Mux_h I__2454 (
            .O(N__17400),
            .I(N__17389));
    LocalMux I__2453 (
            .O(N__17397),
            .I(N__17389));
    LocalMux I__2452 (
            .O(N__17394),
            .I(\POWERLED.countZ0Z_11 ));
    Odrv4 I__2451 (
            .O(N__17389),
            .I(\POWERLED.countZ0Z_11 ));
    CascadeMux I__2450 (
            .O(N__17384),
            .I(N__17381));
    InMux I__2449 (
            .O(N__17381),
            .I(N__17378));
    LocalMux I__2448 (
            .O(N__17378),
            .I(\POWERLED.N_5046_i ));
    InMux I__2447 (
            .O(N__17375),
            .I(N__17372));
    LocalMux I__2446 (
            .O(N__17372),
            .I(N__17368));
    CascadeMux I__2445 (
            .O(N__17371),
            .I(N__17365));
    Span4Mux_v I__2444 (
            .O(N__17368),
            .I(N__17361));
    InMux I__2443 (
            .O(N__17365),
            .I(N__17358));
    InMux I__2442 (
            .O(N__17364),
            .I(N__17355));
    Span4Mux_h I__2441 (
            .O(N__17361),
            .I(N__17350));
    LocalMux I__2440 (
            .O(N__17358),
            .I(N__17350));
    LocalMux I__2439 (
            .O(N__17355),
            .I(\POWERLED.countZ0Z_12 ));
    Odrv4 I__2438 (
            .O(N__17350),
            .I(\POWERLED.countZ0Z_12 ));
    CascadeMux I__2437 (
            .O(N__17345),
            .I(N__17342));
    InMux I__2436 (
            .O(N__17342),
            .I(N__17339));
    LocalMux I__2435 (
            .O(N__17339),
            .I(N__17336));
    Odrv4 I__2434 (
            .O(N__17336),
            .I(\POWERLED.N_5047_i ));
    InMux I__2433 (
            .O(N__17333),
            .I(N__17330));
    LocalMux I__2432 (
            .O(N__17330),
            .I(N__17325));
    InMux I__2431 (
            .O(N__17329),
            .I(N__17322));
    CascadeMux I__2430 (
            .O(N__17328),
            .I(N__17319));
    Span4Mux_v I__2429 (
            .O(N__17325),
            .I(N__17316));
    LocalMux I__2428 (
            .O(N__17322),
            .I(N__17313));
    InMux I__2427 (
            .O(N__17319),
            .I(N__17310));
    Odrv4 I__2426 (
            .O(N__17316),
            .I(\POWERLED.countZ0Z_13 ));
    Odrv4 I__2425 (
            .O(N__17313),
            .I(\POWERLED.countZ0Z_13 ));
    LocalMux I__2424 (
            .O(N__17310),
            .I(\POWERLED.countZ0Z_13 ));
    InMux I__2423 (
            .O(N__17303),
            .I(N__17300));
    LocalMux I__2422 (
            .O(N__17300),
            .I(\POWERLED.N_5048_i ));
    InMux I__2421 (
            .O(N__17297),
            .I(N__17294));
    LocalMux I__2420 (
            .O(N__17294),
            .I(N__17289));
    InMux I__2419 (
            .O(N__17293),
            .I(N__17286));
    CascadeMux I__2418 (
            .O(N__17292),
            .I(N__17283));
    Span4Mux_h I__2417 (
            .O(N__17289),
            .I(N__17280));
    LocalMux I__2416 (
            .O(N__17286),
            .I(N__17277));
    InMux I__2415 (
            .O(N__17283),
            .I(N__17274));
    Odrv4 I__2414 (
            .O(N__17280),
            .I(\POWERLED.countZ0Z_14 ));
    Odrv4 I__2413 (
            .O(N__17277),
            .I(\POWERLED.countZ0Z_14 ));
    LocalMux I__2412 (
            .O(N__17274),
            .I(\POWERLED.countZ0Z_14 ));
    InMux I__2411 (
            .O(N__17267),
            .I(N__17264));
    LocalMux I__2410 (
            .O(N__17264),
            .I(\POWERLED.N_5049_i ));
    InMux I__2409 (
            .O(N__17261),
            .I(N__17258));
    LocalMux I__2408 (
            .O(N__17258),
            .I(N__17255));
    Span4Mux_v I__2407 (
            .O(N__17255),
            .I(N__17248));
    InMux I__2406 (
            .O(N__17254),
            .I(N__17241));
    InMux I__2405 (
            .O(N__17253),
            .I(N__17241));
    InMux I__2404 (
            .O(N__17252),
            .I(N__17241));
    InMux I__2403 (
            .O(N__17251),
            .I(N__17238));
    Odrv4 I__2402 (
            .O(N__17248),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__2401 (
            .O(N__17241),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__2400 (
            .O(N__17238),
            .I(\POWERLED.countZ0Z_0 ));
    CascadeMux I__2399 (
            .O(N__17231),
            .I(N__17228));
    InMux I__2398 (
            .O(N__17228),
            .I(N__17225));
    LocalMux I__2397 (
            .O(N__17225),
            .I(\POWERLED.un1_count_cry_0_i ));
    InMux I__2396 (
            .O(N__17222),
            .I(N__17219));
    LocalMux I__2395 (
            .O(N__17219),
            .I(N__17215));
    CascadeMux I__2394 (
            .O(N__17218),
            .I(N__17211));
    Span12Mux_s6_v I__2393 (
            .O(N__17215),
            .I(N__17208));
    InMux I__2392 (
            .O(N__17214),
            .I(N__17205));
    InMux I__2391 (
            .O(N__17211),
            .I(N__17202));
    Odrv12 I__2390 (
            .O(N__17208),
            .I(\POWERLED.countZ0Z_1 ));
    LocalMux I__2389 (
            .O(N__17205),
            .I(\POWERLED.countZ0Z_1 ));
    LocalMux I__2388 (
            .O(N__17202),
            .I(\POWERLED.countZ0Z_1 ));
    CascadeMux I__2387 (
            .O(N__17195),
            .I(N__17192));
    InMux I__2386 (
            .O(N__17192),
            .I(N__17189));
    LocalMux I__2385 (
            .O(N__17189),
            .I(N__17186));
    Odrv4 I__2384 (
            .O(N__17186),
            .I(\POWERLED.N_5036_i ));
    InMux I__2383 (
            .O(N__17183),
            .I(N__17180));
    LocalMux I__2382 (
            .O(N__17180),
            .I(N__17176));
    CascadeMux I__2381 (
            .O(N__17179),
            .I(N__17173));
    Span4Mux_s3_v I__2380 (
            .O(N__17176),
            .I(N__17170));
    InMux I__2379 (
            .O(N__17173),
            .I(N__17166));
    Span4Mux_v I__2378 (
            .O(N__17170),
            .I(N__17163));
    InMux I__2377 (
            .O(N__17169),
            .I(N__17160));
    LocalMux I__2376 (
            .O(N__17166),
            .I(N__17157));
    Odrv4 I__2375 (
            .O(N__17163),
            .I(\POWERLED.countZ0Z_2 ));
    LocalMux I__2374 (
            .O(N__17160),
            .I(\POWERLED.countZ0Z_2 ));
    Odrv4 I__2373 (
            .O(N__17157),
            .I(\POWERLED.countZ0Z_2 ));
    CascadeMux I__2372 (
            .O(N__17150),
            .I(N__17147));
    InMux I__2371 (
            .O(N__17147),
            .I(N__17144));
    LocalMux I__2370 (
            .O(N__17144),
            .I(\POWERLED.N_5037_i ));
    InMux I__2369 (
            .O(N__17141),
            .I(N__17137));
    CascadeMux I__2368 (
            .O(N__17140),
            .I(N__17134));
    LocalMux I__2367 (
            .O(N__17137),
            .I(N__17131));
    InMux I__2366 (
            .O(N__17134),
            .I(N__17127));
    Span12Mux_s7_v I__2365 (
            .O(N__17131),
            .I(N__17124));
    InMux I__2364 (
            .O(N__17130),
            .I(N__17121));
    LocalMux I__2363 (
            .O(N__17127),
            .I(N__17118));
    Odrv12 I__2362 (
            .O(N__17124),
            .I(\POWERLED.countZ0Z_3 ));
    LocalMux I__2361 (
            .O(N__17121),
            .I(\POWERLED.countZ0Z_3 ));
    Odrv4 I__2360 (
            .O(N__17118),
            .I(\POWERLED.countZ0Z_3 ));
    CascadeMux I__2359 (
            .O(N__17111),
            .I(N__17108));
    InMux I__2358 (
            .O(N__17108),
            .I(N__17105));
    LocalMux I__2357 (
            .O(N__17105),
            .I(\POWERLED.N_5038_i ));
    InMux I__2356 (
            .O(N__17102),
            .I(N__17099));
    LocalMux I__2355 (
            .O(N__17099),
            .I(N__17095));
    CascadeMux I__2354 (
            .O(N__17098),
            .I(N__17091));
    Span4Mux_v I__2353 (
            .O(N__17095),
            .I(N__17088));
    InMux I__2352 (
            .O(N__17094),
            .I(N__17085));
    InMux I__2351 (
            .O(N__17091),
            .I(N__17082));
    Odrv4 I__2350 (
            .O(N__17088),
            .I(\POWERLED.countZ0Z_4 ));
    LocalMux I__2349 (
            .O(N__17085),
            .I(\POWERLED.countZ0Z_4 ));
    LocalMux I__2348 (
            .O(N__17082),
            .I(\POWERLED.countZ0Z_4 ));
    CascadeMux I__2347 (
            .O(N__17075),
            .I(N__17072));
    InMux I__2346 (
            .O(N__17072),
            .I(N__17069));
    LocalMux I__2345 (
            .O(N__17069),
            .I(\POWERLED.N_5039_i ));
    InMux I__2344 (
            .O(N__17066),
            .I(N__17063));
    LocalMux I__2343 (
            .O(N__17063),
            .I(N__17060));
    Span4Mux_v I__2342 (
            .O(N__17060),
            .I(N__17055));
    InMux I__2341 (
            .O(N__17059),
            .I(N__17052));
    CascadeMux I__2340 (
            .O(N__17058),
            .I(N__17049));
    Span4Mux_h I__2339 (
            .O(N__17055),
            .I(N__17046));
    LocalMux I__2338 (
            .O(N__17052),
            .I(N__17043));
    InMux I__2337 (
            .O(N__17049),
            .I(N__17040));
    Odrv4 I__2336 (
            .O(N__17046),
            .I(\POWERLED.countZ0Z_5 ));
    Odrv4 I__2335 (
            .O(N__17043),
            .I(\POWERLED.countZ0Z_5 ));
    LocalMux I__2334 (
            .O(N__17040),
            .I(\POWERLED.countZ0Z_5 ));
    CascadeMux I__2333 (
            .O(N__17033),
            .I(N__17030));
    InMux I__2332 (
            .O(N__17030),
            .I(N__17027));
    LocalMux I__2331 (
            .O(N__17027),
            .I(\POWERLED.N_5040_i ));
    InMux I__2330 (
            .O(N__17024),
            .I(N__17021));
    LocalMux I__2329 (
            .O(N__17021),
            .I(N__17016));
    InMux I__2328 (
            .O(N__17020),
            .I(N__17013));
    CascadeMux I__2327 (
            .O(N__17019),
            .I(N__17010));
    Span4Mux_v I__2326 (
            .O(N__17016),
            .I(N__17007));
    LocalMux I__2325 (
            .O(N__17013),
            .I(N__17004));
    InMux I__2324 (
            .O(N__17010),
            .I(N__17001));
    Odrv4 I__2323 (
            .O(N__17007),
            .I(\POWERLED.countZ0Z_6 ));
    Odrv4 I__2322 (
            .O(N__17004),
            .I(\POWERLED.countZ0Z_6 ));
    LocalMux I__2321 (
            .O(N__17001),
            .I(\POWERLED.countZ0Z_6 ));
    CascadeMux I__2320 (
            .O(N__16994),
            .I(N__16991));
    InMux I__2319 (
            .O(N__16991),
            .I(N__16988));
    LocalMux I__2318 (
            .O(N__16988),
            .I(N__16985));
    Odrv4 I__2317 (
            .O(N__16985),
            .I(\POWERLED.N_5041_i ));
    InMux I__2316 (
            .O(N__16982),
            .I(N__16979));
    LocalMux I__2315 (
            .O(N__16979),
            .I(N__16976));
    Span4Mux_v I__2314 (
            .O(N__16976),
            .I(N__16971));
    InMux I__2313 (
            .O(N__16975),
            .I(N__16968));
    InMux I__2312 (
            .O(N__16974),
            .I(N__16965));
    Odrv4 I__2311 (
            .O(N__16971),
            .I(\POWERLED.countZ0Z_7 ));
    LocalMux I__2310 (
            .O(N__16968),
            .I(\POWERLED.countZ0Z_7 ));
    LocalMux I__2309 (
            .O(N__16965),
            .I(\POWERLED.countZ0Z_7 ));
    InMux I__2308 (
            .O(N__16958),
            .I(N__16955));
    LocalMux I__2307 (
            .O(N__16955),
            .I(N__16952));
    Odrv12 I__2306 (
            .O(N__16952),
            .I(\POWERLED.mult1_un117_sum_i_8 ));
    CascadeMux I__2305 (
            .O(N__16949),
            .I(N__16946));
    InMux I__2304 (
            .O(N__16946),
            .I(N__16943));
    LocalMux I__2303 (
            .O(N__16943),
            .I(\POWERLED.N_5042_i ));
    CascadeMux I__2302 (
            .O(N__16940),
            .I(\POWERLED.mult1_un110_sum_s_8_cascade_ ));
    CascadeMux I__2301 (
            .O(N__16937),
            .I(N__16934));
    InMux I__2300 (
            .O(N__16934),
            .I(N__16931));
    LocalMux I__2299 (
            .O(N__16931),
            .I(\POWERLED.mult1_un103_sum_cry_3_s ));
    InMux I__2298 (
            .O(N__16928),
            .I(\POWERLED.mult1_un103_sum_cry_2 ));
    InMux I__2297 (
            .O(N__16925),
            .I(N__16922));
    LocalMux I__2296 (
            .O(N__16922),
            .I(\POWERLED.mult1_un103_sum_cry_4_s ));
    InMux I__2295 (
            .O(N__16919),
            .I(\POWERLED.mult1_un103_sum_cry_3 ));
    CascadeMux I__2294 (
            .O(N__16916),
            .I(N__16913));
    InMux I__2293 (
            .O(N__16913),
            .I(N__16910));
    LocalMux I__2292 (
            .O(N__16910),
            .I(\POWERLED.mult1_un103_sum_cry_5_s ));
    InMux I__2291 (
            .O(N__16907),
            .I(\POWERLED.mult1_un103_sum_cry_4 ));
    InMux I__2290 (
            .O(N__16904),
            .I(N__16901));
    LocalMux I__2289 (
            .O(N__16901),
            .I(\POWERLED.mult1_un103_sum_cry_6_s ));
    InMux I__2288 (
            .O(N__16898),
            .I(\POWERLED.mult1_un103_sum_cry_5 ));
    CascadeMux I__2287 (
            .O(N__16895),
            .I(N__16892));
    InMux I__2286 (
            .O(N__16892),
            .I(N__16889));
    LocalMux I__2285 (
            .O(N__16889),
            .I(\POWERLED.mult1_un110_sum_axb_8 ));
    InMux I__2284 (
            .O(N__16886),
            .I(\POWERLED.mult1_un103_sum_cry_6 ));
    InMux I__2283 (
            .O(N__16883),
            .I(\POWERLED.mult1_un103_sum_cry_7 ));
    CascadeMux I__2282 (
            .O(N__16880),
            .I(\POWERLED.mult1_un103_sum_s_8_cascade_ ));
    CascadeMux I__2281 (
            .O(N__16877),
            .I(N__16873));
    CascadeMux I__2280 (
            .O(N__16876),
            .I(N__16869));
    InMux I__2279 (
            .O(N__16873),
            .I(N__16862));
    InMux I__2278 (
            .O(N__16872),
            .I(N__16862));
    InMux I__2277 (
            .O(N__16869),
            .I(N__16862));
    LocalMux I__2276 (
            .O(N__16862),
            .I(\POWERLED.mult1_un103_sum_i_0_8 ));
    CascadeMux I__2275 (
            .O(N__16859),
            .I(N__16855));
    CascadeMux I__2274 (
            .O(N__16858),
            .I(N__16851));
    InMux I__2273 (
            .O(N__16855),
            .I(N__16844));
    InMux I__2272 (
            .O(N__16854),
            .I(N__16844));
    InMux I__2271 (
            .O(N__16851),
            .I(N__16844));
    LocalMux I__2270 (
            .O(N__16844),
            .I(\POWERLED.mult1_un110_sum_i_0_8 ));
    CascadeMux I__2269 (
            .O(N__16841),
            .I(N__16838));
    InMux I__2268 (
            .O(N__16838),
            .I(N__16835));
    LocalMux I__2267 (
            .O(N__16835),
            .I(\POWERLED.mult1_un110_sum_cry_3_s ));
    InMux I__2266 (
            .O(N__16832),
            .I(\POWERLED.mult1_un110_sum_cry_2 ));
    InMux I__2265 (
            .O(N__16829),
            .I(N__16826));
    LocalMux I__2264 (
            .O(N__16826),
            .I(\POWERLED.mult1_un110_sum_cry_4_s ));
    InMux I__2263 (
            .O(N__16823),
            .I(\POWERLED.mult1_un110_sum_cry_3 ));
    InMux I__2262 (
            .O(N__16820),
            .I(N__16817));
    LocalMux I__2261 (
            .O(N__16817),
            .I(\POWERLED.mult1_un110_sum_cry_5_s ));
    InMux I__2260 (
            .O(N__16814),
            .I(\POWERLED.mult1_un110_sum_cry_4 ));
    InMux I__2259 (
            .O(N__16811),
            .I(N__16808));
    LocalMux I__2258 (
            .O(N__16808),
            .I(\POWERLED.mult1_un110_sum_cry_6_s ));
    InMux I__2257 (
            .O(N__16805),
            .I(\POWERLED.mult1_un110_sum_cry_5 ));
    InMux I__2256 (
            .O(N__16802),
            .I(N__16799));
    LocalMux I__2255 (
            .O(N__16799),
            .I(\POWERLED.mult1_un117_sum_axb_8 ));
    InMux I__2254 (
            .O(N__16796),
            .I(\POWERLED.mult1_un110_sum_cry_6 ));
    InMux I__2253 (
            .O(N__16793),
            .I(\POWERLED.mult1_un110_sum_cry_7 ));
    CascadeMux I__2252 (
            .O(N__16790),
            .I(N__16786));
    CascadeMux I__2251 (
            .O(N__16789),
            .I(N__16783));
    InMux I__2250 (
            .O(N__16786),
            .I(N__16778));
    InMux I__2249 (
            .O(N__16783),
            .I(N__16773));
    InMux I__2248 (
            .O(N__16782),
            .I(N__16773));
    InMux I__2247 (
            .O(N__16781),
            .I(N__16770));
    LocalMux I__2246 (
            .O(N__16778),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__2245 (
            .O(N__16773),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__2244 (
            .O(N__16770),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    InMux I__2243 (
            .O(N__16763),
            .I(\POWERLED.mult1_un124_sum_cry_7 ));
    InMux I__2242 (
            .O(N__16760),
            .I(N__16757));
    LocalMux I__2241 (
            .O(N__16757),
            .I(\POWERLED.mult1_un124_sum_axb_7_l_fx ));
    InMux I__2240 (
            .O(N__16754),
            .I(N__16751));
    LocalMux I__2239 (
            .O(N__16751),
            .I(N__16747));
    InMux I__2238 (
            .O(N__16750),
            .I(N__16744));
    Odrv4 I__2237 (
            .O(N__16747),
            .I(\POWERLED.mult1_un117_sum_cry_3_s ));
    LocalMux I__2236 (
            .O(N__16744),
            .I(\POWERLED.mult1_un117_sum_cry_3_s ));
    InMux I__2235 (
            .O(N__16739),
            .I(\POWERLED.mult1_un117_sum_cry_2 ));
    CascadeMux I__2234 (
            .O(N__16736),
            .I(N__16733));
    InMux I__2233 (
            .O(N__16733),
            .I(N__16730));
    LocalMux I__2232 (
            .O(N__16730),
            .I(\POWERLED.mult1_un117_sum_cry_4_s ));
    InMux I__2231 (
            .O(N__16727),
            .I(\POWERLED.mult1_un117_sum_cry_3 ));
    InMux I__2230 (
            .O(N__16724),
            .I(N__16721));
    LocalMux I__2229 (
            .O(N__16721),
            .I(\POWERLED.mult1_un117_sum_cry_5_s ));
    InMux I__2228 (
            .O(N__16718),
            .I(\POWERLED.mult1_un117_sum_cry_4 ));
    CascadeMux I__2227 (
            .O(N__16715),
            .I(N__16712));
    InMux I__2226 (
            .O(N__16712),
            .I(N__16706));
    InMux I__2225 (
            .O(N__16711),
            .I(N__16706));
    LocalMux I__2224 (
            .O(N__16706),
            .I(\POWERLED.mult1_un117_sum_cry_6_s ));
    InMux I__2223 (
            .O(N__16703),
            .I(\POWERLED.mult1_un117_sum_cry_5 ));
    InMux I__2222 (
            .O(N__16700),
            .I(N__16697));
    LocalMux I__2221 (
            .O(N__16697),
            .I(\POWERLED.mult1_un124_sum_axb_8 ));
    InMux I__2220 (
            .O(N__16694),
            .I(\POWERLED.mult1_un117_sum_cry_6 ));
    InMux I__2219 (
            .O(N__16691),
            .I(\POWERLED.mult1_un117_sum_cry_7 ));
    InMux I__2218 (
            .O(N__16688),
            .I(N__16685));
    LocalMux I__2217 (
            .O(N__16685),
            .I(N__16679));
    InMux I__2216 (
            .O(N__16684),
            .I(N__16674));
    InMux I__2215 (
            .O(N__16683),
            .I(N__16674));
    CascadeMux I__2214 (
            .O(N__16682),
            .I(N__16671));
    Span12Mux_s4_v I__2213 (
            .O(N__16679),
            .I(N__16665));
    LocalMux I__2212 (
            .O(N__16674),
            .I(N__16662));
    InMux I__2211 (
            .O(N__16671),
            .I(N__16655));
    InMux I__2210 (
            .O(N__16670),
            .I(N__16655));
    InMux I__2209 (
            .O(N__16669),
            .I(N__16655));
    InMux I__2208 (
            .O(N__16668),
            .I(N__16652));
    Odrv12 I__2207 (
            .O(N__16665),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    Odrv4 I__2206 (
            .O(N__16662),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__2205 (
            .O(N__16655),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__2204 (
            .O(N__16652),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    InMux I__2203 (
            .O(N__16643),
            .I(N__16640));
    LocalMux I__2202 (
            .O(N__16640),
            .I(N__16637));
    Span4Mux_v I__2201 (
            .O(N__16637),
            .I(N__16634));
    Odrv4 I__2200 (
            .O(N__16634),
            .I(\POWERLED.mult1_un117_sum_i ));
    CascadeMux I__2199 (
            .O(N__16631),
            .I(N__16628));
    InMux I__2198 (
            .O(N__16628),
            .I(N__16625));
    LocalMux I__2197 (
            .O(N__16625),
            .I(N__16622));
    Odrv12 I__2196 (
            .O(N__16622),
            .I(\POWERLED.mult1_un117_sum_i_0_8 ));
    InMux I__2195 (
            .O(N__16619),
            .I(\POWERLED.mult1_un124_sum_cry_2 ));
    CascadeMux I__2194 (
            .O(N__16616),
            .I(N__16613));
    InMux I__2193 (
            .O(N__16613),
            .I(N__16610));
    LocalMux I__2192 (
            .O(N__16610),
            .I(N__16607));
    Odrv4 I__2191 (
            .O(N__16607),
            .I(\POWERLED.mult1_un124_sum_axb_4_l_fx ));
    InMux I__2190 (
            .O(N__16604),
            .I(\POWERLED.mult1_un124_sum_cry_3 ));
    InMux I__2189 (
            .O(N__16601),
            .I(\POWERLED.mult1_un124_sum_cry_4 ));
    InMux I__2188 (
            .O(N__16598),
            .I(\POWERLED.mult1_un124_sum_cry_5 ));
    InMux I__2187 (
            .O(N__16595),
            .I(\POWERLED.mult1_un124_sum_cry_6 ));
    InMux I__2186 (
            .O(N__16592),
            .I(N__16589));
    LocalMux I__2185 (
            .O(N__16589),
            .I(\VPP_VDDQ.count_2_0_12 ));
    InMux I__2184 (
            .O(N__16586),
            .I(N__16583));
    LocalMux I__2183 (
            .O(N__16583),
            .I(\VPP_VDDQ.count_2_0_13 ));
    InMux I__2182 (
            .O(N__16580),
            .I(N__16577));
    LocalMux I__2181 (
            .O(N__16577),
            .I(\VPP_VDDQ.count_2_0_14 ));
    InMux I__2180 (
            .O(N__16574),
            .I(N__16571));
    LocalMux I__2179 (
            .O(N__16571),
            .I(N__16561));
    InMux I__2178 (
            .O(N__16570),
            .I(N__16556));
    InMux I__2177 (
            .O(N__16569),
            .I(N__16556));
    InMux I__2176 (
            .O(N__16568),
            .I(N__16551));
    InMux I__2175 (
            .O(N__16567),
            .I(N__16551));
    InMux I__2174 (
            .O(N__16566),
            .I(N__16544));
    InMux I__2173 (
            .O(N__16565),
            .I(N__16544));
    InMux I__2172 (
            .O(N__16564),
            .I(N__16544));
    Span4Mux_h I__2171 (
            .O(N__16561),
            .I(N__16539));
    LocalMux I__2170 (
            .O(N__16556),
            .I(N__16539));
    LocalMux I__2169 (
            .O(N__16551),
            .I(\POWERLED.N_2305_i ));
    LocalMux I__2168 (
            .O(N__16544),
            .I(\POWERLED.N_2305_i ));
    Odrv4 I__2167 (
            .O(N__16539),
            .I(\POWERLED.N_2305_i ));
    InMux I__2166 (
            .O(N__16532),
            .I(N__16529));
    LocalMux I__2165 (
            .O(N__16529),
            .I(N__16526));
    Span4Mux_h I__2164 (
            .O(N__16526),
            .I(N__16522));
    InMux I__2163 (
            .O(N__16525),
            .I(N__16519));
    Span4Mux_v I__2162 (
            .O(N__16522),
            .I(N__16516));
    LocalMux I__2161 (
            .O(N__16519),
            .I(\POWERLED.N_660 ));
    Odrv4 I__2160 (
            .O(N__16516),
            .I(\POWERLED.N_660 ));
    InMux I__2159 (
            .O(N__16511),
            .I(N__16508));
    LocalMux I__2158 (
            .O(N__16508),
            .I(N__16505));
    Span4Mux_v I__2157 (
            .O(N__16505),
            .I(N__16502));
    Odrv4 I__2156 (
            .O(N__16502),
            .I(\POWERLED.curr_state_1_0 ));
    CascadeMux I__2155 (
            .O(N__16499),
            .I(N__16496));
    InMux I__2154 (
            .O(N__16496),
            .I(N__16488));
    InMux I__2153 (
            .O(N__16495),
            .I(N__16485));
    InMux I__2152 (
            .O(N__16494),
            .I(N__16482));
    InMux I__2151 (
            .O(N__16493),
            .I(N__16479));
    InMux I__2150 (
            .O(N__16492),
            .I(N__16476));
    InMux I__2149 (
            .O(N__16491),
            .I(N__16473));
    LocalMux I__2148 (
            .O(N__16488),
            .I(N__16470));
    LocalMux I__2147 (
            .O(N__16485),
            .I(N__16458));
    LocalMux I__2146 (
            .O(N__16482),
            .I(N__16455));
    LocalMux I__2145 (
            .O(N__16479),
            .I(N__16452));
    LocalMux I__2144 (
            .O(N__16476),
            .I(N__16449));
    LocalMux I__2143 (
            .O(N__16473),
            .I(N__16446));
    Glb2LocalMux I__2142 (
            .O(N__16470),
            .I(N__16415));
    CEMux I__2141 (
            .O(N__16469),
            .I(N__16415));
    CEMux I__2140 (
            .O(N__16468),
            .I(N__16415));
    CEMux I__2139 (
            .O(N__16467),
            .I(N__16415));
    CEMux I__2138 (
            .O(N__16466),
            .I(N__16415));
    CEMux I__2137 (
            .O(N__16465),
            .I(N__16415));
    CEMux I__2136 (
            .O(N__16464),
            .I(N__16415));
    CEMux I__2135 (
            .O(N__16463),
            .I(N__16415));
    CEMux I__2134 (
            .O(N__16462),
            .I(N__16415));
    CEMux I__2133 (
            .O(N__16461),
            .I(N__16415));
    Glb2LocalMux I__2132 (
            .O(N__16458),
            .I(N__16415));
    Glb2LocalMux I__2131 (
            .O(N__16455),
            .I(N__16415));
    Glb2LocalMux I__2130 (
            .O(N__16452),
            .I(N__16415));
    Glb2LocalMux I__2129 (
            .O(N__16449),
            .I(N__16415));
    Glb2LocalMux I__2128 (
            .O(N__16446),
            .I(N__16415));
    GlobalMux I__2127 (
            .O(N__16415),
            .I(N__16412));
    gio2CtrlBuf I__2126 (
            .O(N__16412),
            .I(N_557_g));
    InMux I__2125 (
            .O(N__16409),
            .I(N__16406));
    LocalMux I__2124 (
            .O(N__16406),
            .I(N__16403));
    Span4Mux_v I__2123 (
            .O(N__16403),
            .I(N__16397));
    InMux I__2122 (
            .O(N__16402),
            .I(N__16390));
    InMux I__2121 (
            .O(N__16401),
            .I(N__16390));
    InMux I__2120 (
            .O(N__16400),
            .I(N__16390));
    Odrv4 I__2119 (
            .O(N__16397),
            .I(N_639));
    LocalMux I__2118 (
            .O(N__16390),
            .I(N_639));
    InMux I__2117 (
            .O(N__16385),
            .I(N__16381));
    InMux I__2116 (
            .O(N__16384),
            .I(N__16377));
    LocalMux I__2115 (
            .O(N__16381),
            .I(N__16374));
    CascadeMux I__2114 (
            .O(N__16380),
            .I(N__16371));
    LocalMux I__2113 (
            .O(N__16377),
            .I(N__16364));
    Span4Mux_v I__2112 (
            .O(N__16374),
            .I(N__16361));
    InMux I__2111 (
            .O(N__16371),
            .I(N__16350));
    InMux I__2110 (
            .O(N__16370),
            .I(N__16350));
    InMux I__2109 (
            .O(N__16369),
            .I(N__16350));
    InMux I__2108 (
            .O(N__16368),
            .I(N__16350));
    InMux I__2107 (
            .O(N__16367),
            .I(N__16350));
    Span4Mux_h I__2106 (
            .O(N__16364),
            .I(N__16347));
    Odrv4 I__2105 (
            .O(N__16361),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__2104 (
            .O(N__16350),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    Odrv4 I__2103 (
            .O(N__16347),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    CascadeMux I__2102 (
            .O(N__16340),
            .I(N__16337));
    InMux I__2101 (
            .O(N__16337),
            .I(N__16334));
    LocalMux I__2100 (
            .O(N__16334),
            .I(N__16331));
    Span4Mux_v I__2099 (
            .O(N__16331),
            .I(N__16326));
    InMux I__2098 (
            .O(N__16330),
            .I(N__16321));
    InMux I__2097 (
            .O(N__16329),
            .I(N__16321));
    Odrv4 I__2096 (
            .O(N__16326),
            .I(\VPP_VDDQ.curr_state_2_RNIZ0Z_1 ));
    LocalMux I__2095 (
            .O(N__16321),
            .I(\VPP_VDDQ.curr_state_2_RNIZ0Z_1 ));
    CascadeMux I__2094 (
            .O(N__16316),
            .I(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0_cascade_ ));
    InMux I__2093 (
            .O(N__16313),
            .I(N__16310));
    LocalMux I__2092 (
            .O(N__16310),
            .I(\VPP_VDDQ.count_2_0_9 ));
    CascadeMux I__2091 (
            .O(N__16307),
            .I(\VPP_VDDQ.count_2Z0Z_9_cascade_ ));
    InMux I__2090 (
            .O(N__16304),
            .I(N__16301));
    LocalMux I__2089 (
            .O(N__16301),
            .I(\VPP_VDDQ.un9_clk_100khz_7 ));
    InMux I__2088 (
            .O(N__16298),
            .I(N__16292));
    InMux I__2087 (
            .O(N__16297),
            .I(N__16292));
    LocalMux I__2086 (
            .O(N__16292),
            .I(\VPP_VDDQ.count_2Z0Z_7 ));
    InMux I__2085 (
            .O(N__16289),
            .I(N__16286));
    LocalMux I__2084 (
            .O(N__16286),
            .I(\VPP_VDDQ.count_2_0_11 ));
    InMux I__2083 (
            .O(N__16283),
            .I(N__16280));
    LocalMux I__2082 (
            .O(N__16280),
            .I(N__16277));
    Odrv4 I__2081 (
            .O(N__16277),
            .I(\VPP_VDDQ.un9_clk_100khz_10 ));
    CascadeMux I__2080 (
            .O(N__16274),
            .I(\VPP_VDDQ.count_2_1_1_cascade_ ));
    InMux I__2079 (
            .O(N__16271),
            .I(N__16268));
    LocalMux I__2078 (
            .O(N__16268),
            .I(N__16264));
    InMux I__2077 (
            .O(N__16267),
            .I(N__16261));
    Span4Mux_v I__2076 (
            .O(N__16264),
            .I(N__16258));
    LocalMux I__2075 (
            .O(N__16261),
            .I(N__16255));
    Span4Mux_v I__2074 (
            .O(N__16258),
            .I(N__16252));
    IoSpan4Mux I__2073 (
            .O(N__16255),
            .I(N__16249));
    Span4Mux_h I__2072 (
            .O(N__16252),
            .I(N__16246));
    IoSpan4Mux I__2071 (
            .O(N__16249),
            .I(N__16243));
    Odrv4 I__2070 (
            .O(N__16246),
            .I(slp_susn));
    Odrv4 I__2069 (
            .O(N__16243),
            .I(slp_susn));
    InMux I__2068 (
            .O(N__16238),
            .I(N__16235));
    LocalMux I__2067 (
            .O(N__16235),
            .I(N__16232));
    Span4Mux_v I__2066 (
            .O(N__16232),
            .I(N__16229));
    Odrv4 I__2065 (
            .O(N__16229),
            .I(v5a_ok));
    IoInMux I__2064 (
            .O(N__16226),
            .I(N__16222));
    IoInMux I__2063 (
            .O(N__16225),
            .I(N__16218));
    LocalMux I__2062 (
            .O(N__16222),
            .I(N__16215));
    CascadeMux I__2061 (
            .O(N__16221),
            .I(N__16212));
    LocalMux I__2060 (
            .O(N__16218),
            .I(N__16209));
    Span4Mux_s3_h I__2059 (
            .O(N__16215),
            .I(N__16206));
    InMux I__2058 (
            .O(N__16212),
            .I(N__16203));
    IoSpan4Mux I__2057 (
            .O(N__16209),
            .I(N__16200));
    Sp12to4 I__2056 (
            .O(N__16206),
            .I(N__16195));
    LocalMux I__2055 (
            .O(N__16203),
            .I(N__16195));
    IoSpan4Mux I__2054 (
            .O(N__16200),
            .I(N__16192));
    Span12Mux_v I__2053 (
            .O(N__16195),
            .I(N__16189));
    IoSpan4Mux I__2052 (
            .O(N__16192),
            .I(N__16186));
    Odrv12 I__2051 (
            .O(N__16189),
            .I(v33a_ok));
    Odrv4 I__2050 (
            .O(N__16186),
            .I(v33a_ok));
    IoInMux I__2049 (
            .O(N__16181),
            .I(N__16178));
    LocalMux I__2048 (
            .O(N__16178),
            .I(N__16174));
    InMux I__2047 (
            .O(N__16177),
            .I(N__16171));
    Span4Mux_s2_h I__2046 (
            .O(N__16174),
            .I(N__16168));
    LocalMux I__2045 (
            .O(N__16171),
            .I(N__16165));
    Sp12to4 I__2044 (
            .O(N__16168),
            .I(N__16162));
    Span4Mux_v I__2043 (
            .O(N__16165),
            .I(N__16159));
    Span12Mux_s11_v I__2042 (
            .O(N__16162),
            .I(N__16156));
    Span4Mux_v I__2041 (
            .O(N__16159),
            .I(N__16153));
    Odrv12 I__2040 (
            .O(N__16156),
            .I(v1p8a_ok));
    Odrv4 I__2039 (
            .O(N__16153),
            .I(v1p8a_ok));
    CascadeMux I__2038 (
            .O(N__16148),
            .I(rsmrst_pwrgd_signal_cascade_));
    CascadeMux I__2037 (
            .O(N__16145),
            .I(\RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_ ));
    CascadeMux I__2036 (
            .O(N__16142),
            .I(N__16138));
    InMux I__2035 (
            .O(N__16141),
            .I(N__16135));
    InMux I__2034 (
            .O(N__16138),
            .I(N__16132));
    LocalMux I__2033 (
            .O(N__16135),
            .I(N__16127));
    LocalMux I__2032 (
            .O(N__16132),
            .I(N__16127));
    Span4Mux_h I__2031 (
            .O(N__16127),
            .I(N__16124));
    Span4Mux_v I__2030 (
            .O(N__16124),
            .I(N__16121));
    Odrv4 I__2029 (
            .O(N__16121),
            .I(\RSMRST_PWRGD.N_264_i ));
    InMux I__2028 (
            .O(N__16118),
            .I(N__16115));
    LocalMux I__2027 (
            .O(N__16115),
            .I(\VPP_VDDQ.un9_clk_100khz_1 ));
    CascadeMux I__2026 (
            .O(N__16112),
            .I(\VPP_VDDQ.un9_clk_100khz_13_cascade_ ));
    InMux I__2025 (
            .O(N__16109),
            .I(N__16103));
    InMux I__2024 (
            .O(N__16108),
            .I(N__16103));
    LocalMux I__2023 (
            .O(N__16103),
            .I(N__16099));
    InMux I__2022 (
            .O(N__16102),
            .I(N__16096));
    Span4Mux_s3_h I__2021 (
            .O(N__16099),
            .I(N__16093));
    LocalMux I__2020 (
            .O(N__16096),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv4 I__2019 (
            .O(N__16093),
            .I(\VPP_VDDQ.N_1_i ));
    InMux I__2018 (
            .O(N__16088),
            .I(N__16084));
    InMux I__2017 (
            .O(N__16087),
            .I(N__16080));
    LocalMux I__2016 (
            .O(N__16084),
            .I(N__16077));
    CascadeMux I__2015 (
            .O(N__16083),
            .I(N__16074));
    LocalMux I__2014 (
            .O(N__16080),
            .I(N__16070));
    Span4Mux_v I__2013 (
            .O(N__16077),
            .I(N__16067));
    InMux I__2012 (
            .O(N__16074),
            .I(N__16064));
    InMux I__2011 (
            .O(N__16073),
            .I(N__16061));
    Span4Mux_h I__2010 (
            .O(N__16070),
            .I(N__16058));
    Odrv4 I__2009 (
            .O(N__16067),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    LocalMux I__2008 (
            .O(N__16064),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    LocalMux I__2007 (
            .O(N__16061),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    Odrv4 I__2006 (
            .O(N__16058),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    CascadeMux I__2005 (
            .O(N__16049),
            .I(\VPP_VDDQ.N_1_i_cascade_ ));
    InMux I__2004 (
            .O(N__16046),
            .I(N__16040));
    InMux I__2003 (
            .O(N__16045),
            .I(N__16040));
    LocalMux I__2002 (
            .O(N__16040),
            .I(N__16037));
    Span4Mux_s3_h I__2001 (
            .O(N__16037),
            .I(N__16034));
    Odrv4 I__2000 (
            .O(N__16034),
            .I(\VPP_VDDQ.N_664 ));
    CascadeMux I__1999 (
            .O(N__16031),
            .I(\VPP_VDDQ.count_2_1_sqmuxa_cascade_ ));
    CascadeMux I__1998 (
            .O(N__16028),
            .I(\VPP_VDDQ.count_2_1_0_cascade_ ));
    CascadeMux I__1997 (
            .O(N__16025),
            .I(\VPP_VDDQ.count_2Z0Z_0_cascade_ ));
    InMux I__1996 (
            .O(N__16022),
            .I(N__16019));
    LocalMux I__1995 (
            .O(N__16019),
            .I(\VPP_VDDQ.count_2_0_0 ));
    InMux I__1994 (
            .O(N__16016),
            .I(N__16013));
    LocalMux I__1993 (
            .O(N__16013),
            .I(\VPP_VDDQ.count_2_1_1 ));
    InMux I__1992 (
            .O(N__16010),
            .I(N__16004));
    InMux I__1991 (
            .O(N__16009),
            .I(N__16004));
    LocalMux I__1990 (
            .O(N__16004),
            .I(\VPP_VDDQ.count_2Z0Z_1 ));
    InMux I__1989 (
            .O(N__16001),
            .I(N__15998));
    LocalMux I__1988 (
            .O(N__15998),
            .I(N__15995));
    Span4Mux_v I__1987 (
            .O(N__15995),
            .I(N__15992));
    Span4Mux_h I__1986 (
            .O(N__15992),
            .I(N__15989));
    Odrv4 I__1985 (
            .O(N__15989),
            .I(gpio_fpga_soc_1));
    CascadeMux I__1984 (
            .O(N__15986),
            .I(\HDA_STRAP.m14_i_0_cascade_ ));
    InMux I__1983 (
            .O(N__15983),
            .I(N__15977));
    InMux I__1982 (
            .O(N__15982),
            .I(N__15977));
    LocalMux I__1981 (
            .O(N__15977),
            .I(N__15974));
    Span4Mux_v I__1980 (
            .O(N__15974),
            .I(N__15971));
    Span4Mux_v I__1979 (
            .O(N__15971),
            .I(N__15966));
    InMux I__1978 (
            .O(N__15970),
            .I(N__15963));
    InMux I__1977 (
            .O(N__15969),
            .I(N__15960));
    Odrv4 I__1976 (
            .O(N__15966),
            .I(N_428));
    LocalMux I__1975 (
            .O(N__15963),
            .I(N_428));
    LocalMux I__1974 (
            .O(N__15960),
            .I(N_428));
    InMux I__1973 (
            .O(N__15953),
            .I(N__15938));
    InMux I__1972 (
            .O(N__15952),
            .I(N__15938));
    InMux I__1971 (
            .O(N__15951),
            .I(N__15938));
    InMux I__1970 (
            .O(N__15950),
            .I(N__15938));
    InMux I__1969 (
            .O(N__15949),
            .I(N__15938));
    LocalMux I__1968 (
            .O(N__15938),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    InMux I__1967 (
            .O(N__15935),
            .I(N__15927));
    InMux I__1966 (
            .O(N__15934),
            .I(N__15927));
    CascadeMux I__1965 (
            .O(N__15933),
            .I(N__15924));
    CascadeMux I__1964 (
            .O(N__15932),
            .I(N__15921));
    LocalMux I__1963 (
            .O(N__15927),
            .I(N__15917));
    InMux I__1962 (
            .O(N__15924),
            .I(N__15910));
    InMux I__1961 (
            .O(N__15921),
            .I(N__15910));
    InMux I__1960 (
            .O(N__15920),
            .I(N__15910));
    Odrv4 I__1959 (
            .O(N__15917),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__1958 (
            .O(N__15910),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    InMux I__1957 (
            .O(N__15905),
            .I(N__15901));
    InMux I__1956 (
            .O(N__15904),
            .I(N__15898));
    LocalMux I__1955 (
            .O(N__15901),
            .I(\HDA_STRAP.curr_stateZ0Z_2 ));
    LocalMux I__1954 (
            .O(N__15898),
            .I(\HDA_STRAP.curr_stateZ0Z_2 ));
    InMux I__1953 (
            .O(N__15893),
            .I(N__15890));
    LocalMux I__1952 (
            .O(N__15890),
            .I(\HDA_STRAP.HDA_SDO_ATP_3_0 ));
    CascadeMux I__1951 (
            .O(N__15887),
            .I(\HDA_STRAP.HDA_SDO_ATP_3_0_cascade_ ));
    IoInMux I__1950 (
            .O(N__15884),
            .I(N__15881));
    LocalMux I__1949 (
            .O(N__15881),
            .I(N__15878));
    Span4Mux_s3_h I__1948 (
            .O(N__15878),
            .I(N__15875));
    Span4Mux_v I__1947 (
            .O(N__15875),
            .I(N__15872));
    Odrv4 I__1946 (
            .O(N__15872),
            .I(hda_sdo_atp));
    InMux I__1945 (
            .O(N__15869),
            .I(N__15866));
    LocalMux I__1944 (
            .O(N__15866),
            .I(N__15863));
    Span4Mux_v I__1943 (
            .O(N__15863),
            .I(N__15859));
    CascadeMux I__1942 (
            .O(N__15862),
            .I(N__15856));
    Span4Mux_h I__1941 (
            .O(N__15859),
            .I(N__15853));
    InMux I__1940 (
            .O(N__15856),
            .I(N__15850));
    Odrv4 I__1939 (
            .O(N__15853),
            .I(\PCH_PWRGD.N_670 ));
    LocalMux I__1938 (
            .O(N__15850),
            .I(\PCH_PWRGD.N_670 ));
    InMux I__1937 (
            .O(N__15845),
            .I(N__15842));
    LocalMux I__1936 (
            .O(N__15842),
            .I(N__15836));
    InMux I__1935 (
            .O(N__15841),
            .I(N__15828));
    InMux I__1934 (
            .O(N__15840),
            .I(N__15828));
    InMux I__1933 (
            .O(N__15839),
            .I(N__15828));
    Span4Mux_h I__1932 (
            .O(N__15836),
            .I(N__15825));
    InMux I__1931 (
            .O(N__15835),
            .I(N__15822));
    LocalMux I__1930 (
            .O(N__15828),
            .I(\PCH_PWRGD.N_2266_i ));
    Odrv4 I__1929 (
            .O(N__15825),
            .I(\PCH_PWRGD.N_2266_i ));
    LocalMux I__1928 (
            .O(N__15822),
            .I(\PCH_PWRGD.N_2266_i ));
    CascadeMux I__1927 (
            .O(N__15815),
            .I(N__15812));
    InMux I__1926 (
            .O(N__15812),
            .I(N__15809));
    LocalMux I__1925 (
            .O(N__15809),
            .I(\PCH_PWRGD.N_38_f0 ));
    InMux I__1924 (
            .O(N__15806),
            .I(N__15802));
    InMux I__1923 (
            .O(N__15805),
            .I(N__15799));
    LocalMux I__1922 (
            .O(N__15802),
            .I(N__15793));
    LocalMux I__1921 (
            .O(N__15799),
            .I(N__15793));
    InMux I__1920 (
            .O(N__15798),
            .I(N__15790));
    Span12Mux_s6_v I__1919 (
            .O(N__15793),
            .I(N__15787));
    LocalMux I__1918 (
            .O(N__15790),
            .I(\PCH_PWRGD.curr_state_0_sqmuxa ));
    Odrv12 I__1917 (
            .O(N__15787),
            .I(\PCH_PWRGD.curr_state_0_sqmuxa ));
    CascadeMux I__1916 (
            .O(N__15782),
            .I(\PCH_PWRGD.N_38_f0_cascade_ ));
    InMux I__1915 (
            .O(N__15779),
            .I(N__15775));
    InMux I__1914 (
            .O(N__15778),
            .I(N__15772));
    LocalMux I__1913 (
            .O(N__15775),
            .I(\PCH_PWRGD.delayed_vccin_ok_0 ));
    LocalMux I__1912 (
            .O(N__15772),
            .I(\PCH_PWRGD.delayed_vccin_ok_0 ));
    CascadeMux I__1911 (
            .O(N__15767),
            .I(\VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_ ));
    CascadeMux I__1910 (
            .O(N__15764),
            .I(\HDA_STRAP.N_16_cascade_ ));
    CascadeMux I__1909 (
            .O(N__15761),
            .I(\PCH_PWRGD.delayed_vccin_okZ0_cascade_ ));
    CascadeMux I__1908 (
            .O(N__15758),
            .I(N_428_cascade_));
    InMux I__1907 (
            .O(N__15755),
            .I(N__15749));
    InMux I__1906 (
            .O(N__15754),
            .I(N__15749));
    LocalMux I__1905 (
            .O(N__15749),
            .I(\POWERLED.count_1_5 ));
    InMux I__1904 (
            .O(N__15746),
            .I(N__15743));
    LocalMux I__1903 (
            .O(N__15743),
            .I(\POWERLED.count_0_5 ));
    CascadeMux I__1902 (
            .O(N__15740),
            .I(N__15737));
    InMux I__1901 (
            .O(N__15737),
            .I(N__15731));
    InMux I__1900 (
            .O(N__15736),
            .I(N__15731));
    LocalMux I__1899 (
            .O(N__15731),
            .I(\POWERLED.count_1_14 ));
    InMux I__1898 (
            .O(N__15728),
            .I(N__15725));
    LocalMux I__1897 (
            .O(N__15725),
            .I(\POWERLED.count_0_14 ));
    InMux I__1896 (
            .O(N__15722),
            .I(N__15716));
    InMux I__1895 (
            .O(N__15721),
            .I(N__15716));
    LocalMux I__1894 (
            .O(N__15716),
            .I(\POWERLED.count_1_6 ));
    InMux I__1893 (
            .O(N__15713),
            .I(N__15710));
    LocalMux I__1892 (
            .O(N__15710),
            .I(\POWERLED.count_0_6 ));
    InMux I__1891 (
            .O(N__15707),
            .I(N__15703));
    InMux I__1890 (
            .O(N__15706),
            .I(N__15700));
    LocalMux I__1889 (
            .O(N__15703),
            .I(N__15697));
    LocalMux I__1888 (
            .O(N__15700),
            .I(\POWERLED.count_1_10 ));
    Odrv4 I__1887 (
            .O(N__15697),
            .I(\POWERLED.count_1_10 ));
    InMux I__1886 (
            .O(N__15692),
            .I(N__15689));
    LocalMux I__1885 (
            .O(N__15689),
            .I(N__15686));
    Span4Mux_s2_h I__1884 (
            .O(N__15686),
            .I(N__15683));
    Odrv4 I__1883 (
            .O(N__15683),
            .I(\POWERLED.count_0_10 ));
    IoInMux I__1882 (
            .O(N__15680),
            .I(N__15677));
    LocalMux I__1881 (
            .O(N__15677),
            .I(N__15674));
    Span4Mux_s1_h I__1880 (
            .O(N__15674),
            .I(N__15671));
    Odrv4 I__1879 (
            .O(N__15671),
            .I(v33a_enn));
    CascadeMux I__1878 (
            .O(N__15668),
            .I(N__15665));
    InMux I__1877 (
            .O(N__15665),
            .I(N__15659));
    InMux I__1876 (
            .O(N__15664),
            .I(N__15659));
    LocalMux I__1875 (
            .O(N__15659),
            .I(\POWERLED.un1_count_cry_14_c_RNIDQ1DZ0 ));
    InMux I__1874 (
            .O(N__15656),
            .I(N__15653));
    LocalMux I__1873 (
            .O(N__15653),
            .I(\POWERLED.count_0_15 ));
    InMux I__1872 (
            .O(N__15650),
            .I(N__15644));
    InMux I__1871 (
            .O(N__15649),
            .I(N__15644));
    LocalMux I__1870 (
            .O(N__15644),
            .I(\POWERLED.count_1_7 ));
    InMux I__1869 (
            .O(N__15641),
            .I(N__15638));
    LocalMux I__1868 (
            .O(N__15638),
            .I(\POWERLED.count_0_7 ));
    InMux I__1867 (
            .O(N__15635),
            .I(N__15629));
    InMux I__1866 (
            .O(N__15634),
            .I(N__15629));
    LocalMux I__1865 (
            .O(N__15629),
            .I(\POWERLED.count_1_8 ));
    InMux I__1864 (
            .O(N__15626),
            .I(N__15623));
    LocalMux I__1863 (
            .O(N__15623),
            .I(\POWERLED.count_0_8 ));
    InMux I__1862 (
            .O(N__15620),
            .I(N__15614));
    InMux I__1861 (
            .O(N__15619),
            .I(N__15614));
    LocalMux I__1860 (
            .O(N__15614),
            .I(\POWERLED.count_1_9 ));
    InMux I__1859 (
            .O(N__15611),
            .I(N__15608));
    LocalMux I__1858 (
            .O(N__15608),
            .I(\POWERLED.count_0_9 ));
    CascadeMux I__1857 (
            .O(N__15605),
            .I(N__15602));
    InMux I__1856 (
            .O(N__15602),
            .I(N__15596));
    InMux I__1855 (
            .O(N__15601),
            .I(N__15596));
    LocalMux I__1854 (
            .O(N__15596),
            .I(\POWERLED.count_1_13 ));
    InMux I__1853 (
            .O(N__15593),
            .I(N__15590));
    LocalMux I__1852 (
            .O(N__15590),
            .I(\POWERLED.count_0_13 ));
    SRMux I__1851 (
            .O(N__15587),
            .I(N__15584));
    LocalMux I__1850 (
            .O(N__15584),
            .I(N__15581));
    Span4Mux_v I__1849 (
            .O(N__15581),
            .I(N__15578));
    Odrv4 I__1848 (
            .O(N__15578),
            .I(\POWERLED.pwm_out_1_sqmuxa ));
    InMux I__1847 (
            .O(N__15575),
            .I(N__15572));
    LocalMux I__1846 (
            .O(N__15572),
            .I(\POWERLED.un79_clk_100khzlt6 ));
    CascadeMux I__1845 (
            .O(N__15569),
            .I(\POWERLED.un79_clk_100khzlto15_5_cascade_ ));
    InMux I__1844 (
            .O(N__15566),
            .I(N__15563));
    LocalMux I__1843 (
            .O(N__15563),
            .I(\POWERLED.un79_clk_100khzlto15_4 ));
    CascadeMux I__1842 (
            .O(N__15560),
            .I(\POWERLED.un79_clk_100khzlto15_7_cascade_ ));
    InMux I__1841 (
            .O(N__15557),
            .I(N__15554));
    LocalMux I__1840 (
            .O(N__15554),
            .I(N__15549));
    InMux I__1839 (
            .O(N__15553),
            .I(N__15546));
    InMux I__1838 (
            .O(N__15552),
            .I(N__15543));
    Span4Mux_s1_h I__1837 (
            .O(N__15549),
            .I(N__15538));
    LocalMux I__1836 (
            .O(N__15546),
            .I(N__15538));
    LocalMux I__1835 (
            .O(N__15543),
            .I(\POWERLED.un79_clk_100khz ));
    Odrv4 I__1834 (
            .O(N__15538),
            .I(\POWERLED.un79_clk_100khz ));
    CascadeMux I__1833 (
            .O(N__15533),
            .I(\POWERLED.un79_clk_100khz_cascade_ ));
    CascadeMux I__1832 (
            .O(N__15530),
            .I(N__15527));
    InMux I__1831 (
            .O(N__15527),
            .I(N__15524));
    LocalMux I__1830 (
            .O(N__15524),
            .I(N__15521));
    Odrv4 I__1829 (
            .O(N__15521),
            .I(\POWERLED.g0_2_1 ));
    CascadeMux I__1828 (
            .O(N__15518),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ));
    CascadeMux I__1827 (
            .O(N__15515),
            .I(\VPP_VDDQ.N_60_cascade_ ));
    SRMux I__1826 (
            .O(N__15512),
            .I(N__15509));
    LocalMux I__1825 (
            .O(N__15509),
            .I(N__15506));
    Span4Mux_s2_h I__1824 (
            .O(N__15506),
            .I(N__15503));
    Odrv4 I__1823 (
            .O(N__15503),
            .I(\VPP_VDDQ.N_60_i ));
    InMux I__1822 (
            .O(N__15500),
            .I(N__15493));
    InMux I__1821 (
            .O(N__15499),
            .I(N__15493));
    InMux I__1820 (
            .O(N__15498),
            .I(N__15490));
    LocalMux I__1819 (
            .O(N__15493),
            .I(\VPP_VDDQ.N_60 ));
    LocalMux I__1818 (
            .O(N__15490),
            .I(\VPP_VDDQ.N_60 ));
    CascadeMux I__1817 (
            .O(N__15485),
            .I(N__15481));
    InMux I__1816 (
            .O(N__15484),
            .I(N__15476));
    InMux I__1815 (
            .O(N__15481),
            .I(N__15476));
    LocalMux I__1814 (
            .O(N__15476),
            .I(\VPP_VDDQ.delayed_vddq_okZ0 ));
    InMux I__1813 (
            .O(N__15473),
            .I(N__15467));
    InMux I__1812 (
            .O(N__15472),
            .I(N__15467));
    LocalMux I__1811 (
            .O(N__15467),
            .I(\VPP_VDDQ.delayed_vddq_ok_en ));
    CascadeMux I__1810 (
            .O(N__15464),
            .I(VPP_VDDQ_delayed_vddq_ok_cascade_));
    IoInMux I__1809 (
            .O(N__15461),
            .I(N__15458));
    LocalMux I__1808 (
            .O(N__15458),
            .I(N__15455));
    Span4Mux_s0_v I__1807 (
            .O(N__15455),
            .I(N__15452));
    Span4Mux_v I__1806 (
            .O(N__15452),
            .I(N__15449));
    Span4Mux_v I__1805 (
            .O(N__15449),
            .I(N__15446));
    Odrv4 I__1804 (
            .O(N__15446),
            .I(vccst_pwrgd));
    CascadeMux I__1803 (
            .O(N__15443),
            .I(\VPP_VDDQ.curr_state_2_RNIZ0Z_1_cascade_ ));
    IoInMux I__1802 (
            .O(N__15440),
            .I(N__15436));
    IoInMux I__1801 (
            .O(N__15439),
            .I(N__15433));
    LocalMux I__1800 (
            .O(N__15436),
            .I(N__15430));
    LocalMux I__1799 (
            .O(N__15433),
            .I(N__15427));
    Span4Mux_s1_h I__1798 (
            .O(N__15430),
            .I(N__15424));
    Span12Mux_s10_h I__1797 (
            .O(N__15427),
            .I(N__15421));
    Span4Mux_v I__1796 (
            .O(N__15424),
            .I(N__15418));
    Odrv12 I__1795 (
            .O(N__15421),
            .I(pch_pwrok));
    Odrv4 I__1794 (
            .O(N__15418),
            .I(pch_pwrok));
    InMux I__1793 (
            .O(N__15413),
            .I(N__15410));
    LocalMux I__1792 (
            .O(N__15410),
            .I(\PCH_PWRGD.curr_state_7_0 ));
    InMux I__1791 (
            .O(N__15407),
            .I(N__15403));
    InMux I__1790 (
            .O(N__15406),
            .I(N__15400));
    LocalMux I__1789 (
            .O(N__15403),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__1788 (
            .O(N__15400),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    CascadeMux I__1787 (
            .O(N__15395),
            .I(\PCH_PWRGD.curr_stateZ0Z_0_cascade_ ));
    InMux I__1786 (
            .O(N__15392),
            .I(N__15383));
    InMux I__1785 (
            .O(N__15391),
            .I(N__15383));
    InMux I__1784 (
            .O(N__15390),
            .I(N__15383));
    LocalMux I__1783 (
            .O(N__15383),
            .I(\PCH_PWRGD.N_655 ));
    CascadeMux I__1782 (
            .O(N__15380),
            .I(N__15376));
    InMux I__1781 (
            .O(N__15379),
            .I(N__15370));
    InMux I__1780 (
            .O(N__15376),
            .I(N__15361));
    InMux I__1779 (
            .O(N__15375),
            .I(N__15361));
    InMux I__1778 (
            .O(N__15374),
            .I(N__15361));
    InMux I__1777 (
            .O(N__15373),
            .I(N__15361));
    LocalMux I__1776 (
            .O(N__15370),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__1775 (
            .O(N__15361),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    InMux I__1774 (
            .O(N__15356),
            .I(N__15340));
    InMux I__1773 (
            .O(N__15355),
            .I(N__15340));
    InMux I__1772 (
            .O(N__15354),
            .I(N__15340));
    InMux I__1771 (
            .O(N__15353),
            .I(N__15340));
    CascadeMux I__1770 (
            .O(N__15352),
            .I(N__15337));
    InMux I__1769 (
            .O(N__15351),
            .I(N__15331));
    CascadeMux I__1768 (
            .O(N__15350),
            .I(N__15325));
    CascadeMux I__1767 (
            .O(N__15349),
            .I(N__15320));
    LocalMux I__1766 (
            .O(N__15340),
            .I(N__15316));
    InMux I__1765 (
            .O(N__15337),
            .I(N__15307));
    InMux I__1764 (
            .O(N__15336),
            .I(N__15307));
    InMux I__1763 (
            .O(N__15335),
            .I(N__15307));
    InMux I__1762 (
            .O(N__15334),
            .I(N__15307));
    LocalMux I__1761 (
            .O(N__15331),
            .I(N__15304));
    InMux I__1760 (
            .O(N__15330),
            .I(N__15299));
    InMux I__1759 (
            .O(N__15329),
            .I(N__15299));
    InMux I__1758 (
            .O(N__15328),
            .I(N__15296));
    InMux I__1757 (
            .O(N__15325),
            .I(N__15285));
    InMux I__1756 (
            .O(N__15324),
            .I(N__15285));
    InMux I__1755 (
            .O(N__15323),
            .I(N__15285));
    InMux I__1754 (
            .O(N__15320),
            .I(N__15285));
    InMux I__1753 (
            .O(N__15319),
            .I(N__15285));
    Span4Mux_s1_h I__1752 (
            .O(N__15316),
            .I(N__15280));
    LocalMux I__1751 (
            .O(N__15307),
            .I(N__15280));
    Odrv4 I__1750 (
            .O(N__15304),
            .I(\PCH_PWRGD.N_386 ));
    LocalMux I__1749 (
            .O(N__15299),
            .I(\PCH_PWRGD.N_386 ));
    LocalMux I__1748 (
            .O(N__15296),
            .I(\PCH_PWRGD.N_386 ));
    LocalMux I__1747 (
            .O(N__15285),
            .I(\PCH_PWRGD.N_386 ));
    Odrv4 I__1746 (
            .O(N__15280),
            .I(\PCH_PWRGD.N_386 ));
    CascadeMux I__1745 (
            .O(N__15269),
            .I(\PCH_PWRGD.curr_state_0_sqmuxa_cascade_ ));
    InMux I__1744 (
            .O(N__15266),
            .I(N__15263));
    LocalMux I__1743 (
            .O(N__15263),
            .I(\PCH_PWRGD.curr_state_0_0 ));
    CascadeMux I__1742 (
            .O(N__15260),
            .I(\VPP_VDDQ.N_53_cascade_ ));
    CascadeMux I__1741 (
            .O(N__15257),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ));
    InMux I__1740 (
            .O(N__15254),
            .I(N__15251));
    LocalMux I__1739 (
            .O(N__15251),
            .I(\VPP_VDDQ.curr_state_2_0_1 ));
    InMux I__1738 (
            .O(N__15248),
            .I(N__15245));
    LocalMux I__1737 (
            .O(N__15245),
            .I(\VPP_VDDQ.curr_state_2_0_0 ));
    CascadeMux I__1736 (
            .O(N__15242),
            .I(\VPP_VDDQ.m4_0_0_cascade_ ));
    InMux I__1735 (
            .O(N__15239),
            .I(N__15236));
    LocalMux I__1734 (
            .O(N__15236),
            .I(\PCH_PWRGD.count_1_i_a2_2_0 ));
    InMux I__1733 (
            .O(N__15233),
            .I(N__15230));
    LocalMux I__1732 (
            .O(N__15230),
            .I(N__15225));
    InMux I__1731 (
            .O(N__15229),
            .I(N__15220));
    InMux I__1730 (
            .O(N__15228),
            .I(N__15220));
    Odrv4 I__1729 (
            .O(N__15225),
            .I(\PCH_PWRGD.count_1_i_a2_11_0 ));
    LocalMux I__1728 (
            .O(N__15220),
            .I(\PCH_PWRGD.count_1_i_a2_11_0 ));
    InMux I__1727 (
            .O(N__15215),
            .I(N__15209));
    InMux I__1726 (
            .O(N__15214),
            .I(N__15209));
    LocalMux I__1725 (
            .O(N__15209),
            .I(\PCH_PWRGD.count_rst ));
    InMux I__1724 (
            .O(N__15206),
            .I(N__15203));
    LocalMux I__1723 (
            .O(N__15203),
            .I(\PCH_PWRGD.count_0_15 ));
    InMux I__1722 (
            .O(N__15200),
            .I(N__15191));
    InMux I__1721 (
            .O(N__15199),
            .I(N__15191));
    InMux I__1720 (
            .O(N__15198),
            .I(N__15191));
    LocalMux I__1719 (
            .O(N__15191),
            .I(\PCH_PWRGD.count_rst_1 ));
    InMux I__1718 (
            .O(N__15188),
            .I(N__15182));
    InMux I__1717 (
            .O(N__15187),
            .I(N__15182));
    LocalMux I__1716 (
            .O(N__15182),
            .I(\PCH_PWRGD.count_0_13 ));
    CascadeMux I__1715 (
            .O(N__15179),
            .I(N__15175));
    InMux I__1714 (
            .O(N__15178),
            .I(N__15171));
    InMux I__1713 (
            .O(N__15175),
            .I(N__15168));
    InMux I__1712 (
            .O(N__15174),
            .I(N__15165));
    LocalMux I__1711 (
            .O(N__15171),
            .I(N__15162));
    LocalMux I__1710 (
            .O(N__15168),
            .I(\PCH_PWRGD.count_rst_4 ));
    LocalMux I__1709 (
            .O(N__15165),
            .I(\PCH_PWRGD.count_rst_4 ));
    Odrv4 I__1708 (
            .O(N__15162),
            .I(\PCH_PWRGD.count_rst_4 ));
    InMux I__1707 (
            .O(N__15155),
            .I(N__15152));
    LocalMux I__1706 (
            .O(N__15152),
            .I(N__15148));
    InMux I__1705 (
            .O(N__15151),
            .I(N__15145));
    Odrv12 I__1704 (
            .O(N__15148),
            .I(\PCH_PWRGD.count_0_10 ));
    LocalMux I__1703 (
            .O(N__15145),
            .I(\PCH_PWRGD.count_0_10 ));
    CEMux I__1702 (
            .O(N__15140),
            .I(N__15133));
    CEMux I__1701 (
            .O(N__15139),
            .I(N__15127));
    CEMux I__1700 (
            .O(N__15138),
            .I(N__15124));
    InMux I__1699 (
            .O(N__15137),
            .I(N__15119));
    CEMux I__1698 (
            .O(N__15136),
            .I(N__15119));
    LocalMux I__1697 (
            .O(N__15133),
            .I(N__15116));
    CEMux I__1696 (
            .O(N__15132),
            .I(N__15113));
    InMux I__1695 (
            .O(N__15131),
            .I(N__15108));
    CEMux I__1694 (
            .O(N__15130),
            .I(N__15108));
    LocalMux I__1693 (
            .O(N__15127),
            .I(N__15103));
    LocalMux I__1692 (
            .O(N__15124),
            .I(N__15103));
    LocalMux I__1691 (
            .O(N__15119),
            .I(N__15095));
    Span4Mux_v I__1690 (
            .O(N__15116),
            .I(N__15090));
    LocalMux I__1689 (
            .O(N__15113),
            .I(N__15090));
    LocalMux I__1688 (
            .O(N__15108),
            .I(N__15085));
    Span4Mux_s3_v I__1687 (
            .O(N__15103),
            .I(N__15082));
    InMux I__1686 (
            .O(N__15102),
            .I(N__15073));
    InMux I__1685 (
            .O(N__15101),
            .I(N__15073));
    InMux I__1684 (
            .O(N__15100),
            .I(N__15073));
    InMux I__1683 (
            .O(N__15099),
            .I(N__15073));
    CascadeMux I__1682 (
            .O(N__15098),
            .I(N__15061));
    Span4Mux_h I__1681 (
            .O(N__15095),
            .I(N__15056));
    Span4Mux_v I__1680 (
            .O(N__15090),
            .I(N__15056));
    InMux I__1679 (
            .O(N__15089),
            .I(N__15048));
    InMux I__1678 (
            .O(N__15088),
            .I(N__15048));
    Span4Mux_v I__1677 (
            .O(N__15085),
            .I(N__15041));
    Span4Mux_s1_h I__1676 (
            .O(N__15082),
            .I(N__15041));
    LocalMux I__1675 (
            .O(N__15073),
            .I(N__15041));
    InMux I__1674 (
            .O(N__15072),
            .I(N__15036));
    CEMux I__1673 (
            .O(N__15071),
            .I(N__15036));
    CEMux I__1672 (
            .O(N__15070),
            .I(N__15033));
    InMux I__1671 (
            .O(N__15069),
            .I(N__15026));
    InMux I__1670 (
            .O(N__15068),
            .I(N__15026));
    InMux I__1669 (
            .O(N__15067),
            .I(N__15026));
    InMux I__1668 (
            .O(N__15066),
            .I(N__15019));
    InMux I__1667 (
            .O(N__15065),
            .I(N__15019));
    InMux I__1666 (
            .O(N__15064),
            .I(N__15019));
    InMux I__1665 (
            .O(N__15061),
            .I(N__15013));
    Span4Mux_s0_h I__1664 (
            .O(N__15056),
            .I(N__15010));
    InMux I__1663 (
            .O(N__15055),
            .I(N__15003));
    InMux I__1662 (
            .O(N__15054),
            .I(N__15003));
    InMux I__1661 (
            .O(N__15053),
            .I(N__15003));
    LocalMux I__1660 (
            .O(N__15048),
            .I(N__14998));
    Span4Mux_h I__1659 (
            .O(N__15041),
            .I(N__14998));
    LocalMux I__1658 (
            .O(N__15036),
            .I(N__14989));
    LocalMux I__1657 (
            .O(N__15033),
            .I(N__14989));
    LocalMux I__1656 (
            .O(N__15026),
            .I(N__14989));
    LocalMux I__1655 (
            .O(N__15019),
            .I(N__14989));
    InMux I__1654 (
            .O(N__15018),
            .I(N__14984));
    InMux I__1653 (
            .O(N__15017),
            .I(N__14984));
    InMux I__1652 (
            .O(N__15016),
            .I(N__14981));
    LocalMux I__1651 (
            .O(N__15013),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    Odrv4 I__1650 (
            .O(N__15010),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    LocalMux I__1649 (
            .O(N__15003),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    Odrv4 I__1648 (
            .O(N__14998),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    Odrv12 I__1647 (
            .O(N__14989),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    LocalMux I__1646 (
            .O(N__14984),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    LocalMux I__1645 (
            .O(N__14981),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ));
    SRMux I__1644 (
            .O(N__14966),
            .I(N__14962));
    SRMux I__1643 (
            .O(N__14965),
            .I(N__14954));
    LocalMux I__1642 (
            .O(N__14962),
            .I(N__14951));
    SRMux I__1641 (
            .O(N__14961),
            .I(N__14948));
    InMux I__1640 (
            .O(N__14960),
            .I(N__14945));
    SRMux I__1639 (
            .O(N__14959),
            .I(N__14942));
    InMux I__1638 (
            .O(N__14958),
            .I(N__14918));
    InMux I__1637 (
            .O(N__14957),
            .I(N__14918));
    LocalMux I__1636 (
            .O(N__14954),
            .I(N__14913));
    Span4Mux_v I__1635 (
            .O(N__14951),
            .I(N__14908));
    LocalMux I__1634 (
            .O(N__14948),
            .I(N__14908));
    LocalMux I__1633 (
            .O(N__14945),
            .I(N__14903));
    LocalMux I__1632 (
            .O(N__14942),
            .I(N__14903));
    SRMux I__1631 (
            .O(N__14941),
            .I(N__14900));
    InMux I__1630 (
            .O(N__14940),
            .I(N__14897));
    InMux I__1629 (
            .O(N__14939),
            .I(N__14894));
    InMux I__1628 (
            .O(N__14938),
            .I(N__14885));
    InMux I__1627 (
            .O(N__14937),
            .I(N__14885));
    InMux I__1626 (
            .O(N__14936),
            .I(N__14885));
    InMux I__1625 (
            .O(N__14935),
            .I(N__14885));
    InMux I__1624 (
            .O(N__14934),
            .I(N__14876));
    InMux I__1623 (
            .O(N__14933),
            .I(N__14876));
    InMux I__1622 (
            .O(N__14932),
            .I(N__14876));
    InMux I__1621 (
            .O(N__14931),
            .I(N__14876));
    InMux I__1620 (
            .O(N__14930),
            .I(N__14871));
    SRMux I__1619 (
            .O(N__14929),
            .I(N__14871));
    InMux I__1618 (
            .O(N__14928),
            .I(N__14864));
    InMux I__1617 (
            .O(N__14927),
            .I(N__14864));
    InMux I__1616 (
            .O(N__14926),
            .I(N__14864));
    InMux I__1615 (
            .O(N__14925),
            .I(N__14857));
    InMux I__1614 (
            .O(N__14924),
            .I(N__14857));
    InMux I__1613 (
            .O(N__14923),
            .I(N__14857));
    LocalMux I__1612 (
            .O(N__14918),
            .I(N__14854));
    InMux I__1611 (
            .O(N__14917),
            .I(N__14851));
    SRMux I__1610 (
            .O(N__14916),
            .I(N__14841));
    Span4Mux_v I__1609 (
            .O(N__14913),
            .I(N__14836));
    Span4Mux_h I__1608 (
            .O(N__14908),
            .I(N__14836));
    Span4Mux_h I__1607 (
            .O(N__14903),
            .I(N__14833));
    LocalMux I__1606 (
            .O(N__14900),
            .I(N__14822));
    LocalMux I__1605 (
            .O(N__14897),
            .I(N__14822));
    LocalMux I__1604 (
            .O(N__14894),
            .I(N__14822));
    LocalMux I__1603 (
            .O(N__14885),
            .I(N__14822));
    LocalMux I__1602 (
            .O(N__14876),
            .I(N__14822));
    LocalMux I__1601 (
            .O(N__14871),
            .I(N__14811));
    LocalMux I__1600 (
            .O(N__14864),
            .I(N__14811));
    LocalMux I__1599 (
            .O(N__14857),
            .I(N__14811));
    Span4Mux_h I__1598 (
            .O(N__14854),
            .I(N__14811));
    LocalMux I__1597 (
            .O(N__14851),
            .I(N__14811));
    InMux I__1596 (
            .O(N__14850),
            .I(N__14800));
    InMux I__1595 (
            .O(N__14849),
            .I(N__14800));
    InMux I__1594 (
            .O(N__14848),
            .I(N__14800));
    InMux I__1593 (
            .O(N__14847),
            .I(N__14800));
    InMux I__1592 (
            .O(N__14846),
            .I(N__14800));
    SRMux I__1591 (
            .O(N__14845),
            .I(N__14795));
    InMux I__1590 (
            .O(N__14844),
            .I(N__14795));
    LocalMux I__1589 (
            .O(N__14841),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__1588 (
            .O(N__14836),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__1587 (
            .O(N__14833),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv12 I__1586 (
            .O(N__14822),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__1585 (
            .O(N__14811),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    LocalMux I__1584 (
            .O(N__14800),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    LocalMux I__1583 (
            .O(N__14795),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    CascadeMux I__1582 (
            .O(N__14780),
            .I(\PCH_PWRGD.N_2266_i_cascade_ ));
    InMux I__1581 (
            .O(N__14777),
            .I(N__14774));
    LocalMux I__1580 (
            .O(N__14774),
            .I(\PCH_PWRGD.curr_state_0_1 ));
    CascadeMux I__1579 (
            .O(N__14771),
            .I(\PCH_PWRGD.m6_i_i_a2_cascade_ ));
    CascadeMux I__1578 (
            .O(N__14768),
            .I(\PCH_PWRGD.count_rst_14_cascade_ ));
    InMux I__1577 (
            .O(N__14765),
            .I(N__14762));
    LocalMux I__1576 (
            .O(N__14762),
            .I(\PCH_PWRGD.count_rst_7 ));
    InMux I__1575 (
            .O(N__14759),
            .I(N__14753));
    InMux I__1574 (
            .O(N__14758),
            .I(N__14753));
    LocalMux I__1573 (
            .O(N__14753),
            .I(\PCH_PWRGD.count_0_7 ));
    CascadeMux I__1572 (
            .O(N__14750),
            .I(N__14745));
    CascadeMux I__1571 (
            .O(N__14749),
            .I(N__14742));
    InMux I__1570 (
            .O(N__14748),
            .I(N__14739));
    InMux I__1569 (
            .O(N__14745),
            .I(N__14735));
    InMux I__1568 (
            .O(N__14742),
            .I(N__14732));
    LocalMux I__1567 (
            .O(N__14739),
            .I(N__14729));
    InMux I__1566 (
            .O(N__14738),
            .I(N__14726));
    LocalMux I__1565 (
            .O(N__14735),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    LocalMux I__1564 (
            .O(N__14732),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    Odrv12 I__1563 (
            .O(N__14729),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    LocalMux I__1562 (
            .O(N__14726),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    InMux I__1561 (
            .O(N__14717),
            .I(N__14714));
    LocalMux I__1560 (
            .O(N__14714),
            .I(\PCH_PWRGD.count_1_i_a2_6_0 ));
    InMux I__1559 (
            .O(N__14711),
            .I(N__14708));
    LocalMux I__1558 (
            .O(N__14708),
            .I(N__14705));
    Odrv4 I__1557 (
            .O(N__14705),
            .I(\PCH_PWRGD.count_1_i_a2_4_0 ));
    CascadeMux I__1556 (
            .O(N__14702),
            .I(\PCH_PWRGD.count_1_i_a2_5_0_cascade_ ));
    InMux I__1555 (
            .O(N__14699),
            .I(N__14696));
    LocalMux I__1554 (
            .O(N__14696),
            .I(N__14693));
    Span4Mux_h I__1553 (
            .O(N__14693),
            .I(N__14690));
    Odrv4 I__1552 (
            .O(N__14690),
            .I(\PCH_PWRGD.count_1_i_a2_3_0 ));
    InMux I__1551 (
            .O(N__14687),
            .I(N__14683));
    InMux I__1550 (
            .O(N__14686),
            .I(N__14680));
    LocalMux I__1549 (
            .O(N__14683),
            .I(\PCH_PWRGD.count_1_i_a2_12_0 ));
    LocalMux I__1548 (
            .O(N__14680),
            .I(\PCH_PWRGD.count_1_i_a2_12_0 ));
    CascadeMux I__1547 (
            .O(N__14675),
            .I(N__14671));
    CascadeMux I__1546 (
            .O(N__14674),
            .I(N__14664));
    InMux I__1545 (
            .O(N__14671),
            .I(N__14661));
    InMux I__1544 (
            .O(N__14670),
            .I(N__14658));
    InMux I__1543 (
            .O(N__14669),
            .I(N__14653));
    InMux I__1542 (
            .O(N__14668),
            .I(N__14653));
    InMux I__1541 (
            .O(N__14667),
            .I(N__14650));
    InMux I__1540 (
            .O(N__14664),
            .I(N__14647));
    LocalMux I__1539 (
            .O(N__14661),
            .I(N__14640));
    LocalMux I__1538 (
            .O(N__14658),
            .I(N__14640));
    LocalMux I__1537 (
            .O(N__14653),
            .I(N__14640));
    LocalMux I__1536 (
            .O(N__14650),
            .I(N__14637));
    LocalMux I__1535 (
            .O(N__14647),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    Odrv4 I__1534 (
            .O(N__14640),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    Odrv4 I__1533 (
            .O(N__14637),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    CascadeMux I__1532 (
            .O(N__14630),
            .I(\PCH_PWRGD.count_1_i_a2_12_0_cascade_ ));
    InMux I__1531 (
            .O(N__14627),
            .I(N__14624));
    LocalMux I__1530 (
            .O(N__14624),
            .I(\PCH_PWRGD.count_0_0 ));
    InMux I__1529 (
            .O(N__14621),
            .I(N__14618));
    LocalMux I__1528 (
            .O(N__14618),
            .I(N__14615));
    Odrv4 I__1527 (
            .O(N__14615),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    CascadeMux I__1526 (
            .O(N__14612),
            .I(\PCH_PWRGD.countZ0Z_15_cascade_ ));
    InMux I__1525 (
            .O(N__14609),
            .I(N__14606));
    LocalMux I__1524 (
            .O(N__14606),
            .I(\PCH_PWRGD.un2_count_1_axb_13 ));
    CascadeMux I__1523 (
            .O(N__14603),
            .I(N__14600));
    InMux I__1522 (
            .O(N__14600),
            .I(N__14597));
    LocalMux I__1521 (
            .O(N__14597),
            .I(N__14593));
    InMux I__1520 (
            .O(N__14596),
            .I(N__14590));
    Odrv4 I__1519 (
            .O(N__14593),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    LocalMux I__1518 (
            .O(N__14590),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    InMux I__1517 (
            .O(N__14585),
            .I(N__14581));
    InMux I__1516 (
            .O(N__14584),
            .I(N__14578));
    LocalMux I__1515 (
            .O(N__14581),
            .I(N__14573));
    LocalMux I__1514 (
            .O(N__14578),
            .I(N__14573));
    Odrv4 I__1513 (
            .O(N__14573),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    InMux I__1512 (
            .O(N__14570),
            .I(N__14567));
    LocalMux I__1511 (
            .O(N__14567),
            .I(\PCH_PWRGD.count_1_i_a2_1_0 ));
    CascadeMux I__1510 (
            .O(N__14564),
            .I(\PCH_PWRGD.count_1_i_a2_0_0_cascade_ ));
    InMux I__1509 (
            .O(N__14561),
            .I(N__14558));
    LocalMux I__1508 (
            .O(N__14558),
            .I(\PCH_PWRGD.count_0_5 ));
    CascadeMux I__1507 (
            .O(N__14555),
            .I(\PCH_PWRGD.count_rst_9_cascade_ ));
    CascadeMux I__1506 (
            .O(N__14552),
            .I(N__14549));
    InMux I__1505 (
            .O(N__14549),
            .I(N__14546));
    LocalMux I__1504 (
            .O(N__14546),
            .I(N__14543));
    Odrv4 I__1503 (
            .O(N__14543),
            .I(\PCH_PWRGD.un2_count_1_axb_10 ));
    InMux I__1502 (
            .O(N__14540),
            .I(N__14536));
    InMux I__1501 (
            .O(N__14539),
            .I(N__14533));
    LocalMux I__1500 (
            .O(N__14536),
            .I(N__14530));
    LocalMux I__1499 (
            .O(N__14533),
            .I(N__14527));
    Odrv4 I__1498 (
            .O(N__14530),
            .I(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ));
    Odrv4 I__1497 (
            .O(N__14527),
            .I(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ));
    CascadeMux I__1496 (
            .O(N__14522),
            .I(\PCH_PWRGD.N_386_cascade_ ));
    InMux I__1495 (
            .O(N__14519),
            .I(N__14516));
    LocalMux I__1494 (
            .O(N__14516),
            .I(\PCH_PWRGD.count_0_11 ));
    CascadeMux I__1493 (
            .O(N__14513),
            .I(\PCH_PWRGD.count_rst_3_cascade_ ));
    InMux I__1492 (
            .O(N__14510),
            .I(N__14504));
    InMux I__1491 (
            .O(N__14509),
            .I(N__14501));
    CascadeMux I__1490 (
            .O(N__14508),
            .I(N__14498));
    InMux I__1489 (
            .O(N__14507),
            .I(N__14495));
    LocalMux I__1488 (
            .O(N__14504),
            .I(N__14490));
    LocalMux I__1487 (
            .O(N__14501),
            .I(N__14490));
    InMux I__1486 (
            .O(N__14498),
            .I(N__14487));
    LocalMux I__1485 (
            .O(N__14495),
            .I(N__14482));
    Span4Mux_v I__1484 (
            .O(N__14490),
            .I(N__14482));
    LocalMux I__1483 (
            .O(N__14487),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    Odrv4 I__1482 (
            .O(N__14482),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    CascadeMux I__1481 (
            .O(N__14477),
            .I(\PCH_PWRGD.count_rst_7_cascade_ ));
    InMux I__1480 (
            .O(N__14474),
            .I(N__14470));
    InMux I__1479 (
            .O(N__14473),
            .I(N__14467));
    LocalMux I__1478 (
            .O(N__14470),
            .I(\PCH_PWRGD.un2_count_1_axb_7 ));
    LocalMux I__1477 (
            .O(N__14467),
            .I(\PCH_PWRGD.un2_count_1_axb_7 ));
    CascadeMux I__1476 (
            .O(N__14462),
            .I(N__14458));
    InMux I__1475 (
            .O(N__14461),
            .I(N__14455));
    InMux I__1474 (
            .O(N__14458),
            .I(N__14452));
    LocalMux I__1473 (
            .O(N__14455),
            .I(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ));
    LocalMux I__1472 (
            .O(N__14452),
            .I(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ));
    CascadeMux I__1471 (
            .O(N__14447),
            .I(\PCH_PWRGD.un2_count_1_axb_7_cascade_ ));
    InMux I__1470 (
            .O(N__14444),
            .I(N__14440));
    InMux I__1469 (
            .O(N__14443),
            .I(N__14437));
    LocalMux I__1468 (
            .O(N__14440),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    LocalMux I__1467 (
            .O(N__14437),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    InMux I__1466 (
            .O(N__14432),
            .I(\RSMRST_PWRGD.un1_count_1_cry_11 ));
    InMux I__1465 (
            .O(N__14429),
            .I(N__14425));
    InMux I__1464 (
            .O(N__14428),
            .I(N__14422));
    LocalMux I__1463 (
            .O(N__14425),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    LocalMux I__1462 (
            .O(N__14422),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    InMux I__1461 (
            .O(N__14417),
            .I(\RSMRST_PWRGD.un1_count_1_cry_12 ));
    InMux I__1460 (
            .O(N__14414),
            .I(N__14410));
    InMux I__1459 (
            .O(N__14413),
            .I(N__14407));
    LocalMux I__1458 (
            .O(N__14410),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    LocalMux I__1457 (
            .O(N__14407),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    InMux I__1456 (
            .O(N__14402),
            .I(\RSMRST_PWRGD.un1_count_1_cry_13 ));
    InMux I__1455 (
            .O(N__14399),
            .I(bfn_2_3_0_));
    CascadeMux I__1454 (
            .O(N__14396),
            .I(N__14393));
    InMux I__1453 (
            .O(N__14393),
            .I(N__14389));
    InMux I__1452 (
            .O(N__14392),
            .I(N__14386));
    LocalMux I__1451 (
            .O(N__14389),
            .I(N__14383));
    LocalMux I__1450 (
            .O(N__14386),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    Odrv4 I__1449 (
            .O(N__14383),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    InMux I__1448 (
            .O(N__14378),
            .I(N__14375));
    LocalMux I__1447 (
            .O(N__14375),
            .I(\PCH_PWRGD.count_0_12 ));
    InMux I__1446 (
            .O(N__14372),
            .I(N__14366));
    InMux I__1445 (
            .O(N__14371),
            .I(N__14366));
    LocalMux I__1444 (
            .O(N__14366),
            .I(N__14363));
    Odrv4 I__1443 (
            .O(N__14363),
            .I(\PCH_PWRGD.count_rst_2 ));
    InMux I__1442 (
            .O(N__14360),
            .I(N__14356));
    InMux I__1441 (
            .O(N__14359),
            .I(N__14353));
    LocalMux I__1440 (
            .O(N__14356),
            .I(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ));
    LocalMux I__1439 (
            .O(N__14353),
            .I(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ));
    InMux I__1438 (
            .O(N__14348),
            .I(N__14344));
    InMux I__1437 (
            .O(N__14347),
            .I(N__14341));
    LocalMux I__1436 (
            .O(N__14344),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    LocalMux I__1435 (
            .O(N__14341),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    InMux I__1434 (
            .O(N__14336),
            .I(\RSMRST_PWRGD.un1_count_1_cry_2 ));
    InMux I__1433 (
            .O(N__14333),
            .I(N__14329));
    InMux I__1432 (
            .O(N__14332),
            .I(N__14326));
    LocalMux I__1431 (
            .O(N__14329),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    LocalMux I__1430 (
            .O(N__14326),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    InMux I__1429 (
            .O(N__14321),
            .I(\RSMRST_PWRGD.un1_count_1_cry_3 ));
    CascadeMux I__1428 (
            .O(N__14318),
            .I(N__14315));
    InMux I__1427 (
            .O(N__14315),
            .I(N__14311));
    InMux I__1426 (
            .O(N__14314),
            .I(N__14308));
    LocalMux I__1425 (
            .O(N__14311),
            .I(N__14305));
    LocalMux I__1424 (
            .O(N__14308),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    Odrv4 I__1423 (
            .O(N__14305),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    InMux I__1422 (
            .O(N__14300),
            .I(\RSMRST_PWRGD.un1_count_1_cry_4 ));
    InMux I__1421 (
            .O(N__14297),
            .I(N__14293));
    InMux I__1420 (
            .O(N__14296),
            .I(N__14290));
    LocalMux I__1419 (
            .O(N__14293),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    LocalMux I__1418 (
            .O(N__14290),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    InMux I__1417 (
            .O(N__14285),
            .I(\RSMRST_PWRGD.un1_count_1_cry_5 ));
    InMux I__1416 (
            .O(N__14282),
            .I(N__14278));
    InMux I__1415 (
            .O(N__14281),
            .I(N__14275));
    LocalMux I__1414 (
            .O(N__14278),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    LocalMux I__1413 (
            .O(N__14275),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    InMux I__1412 (
            .O(N__14270),
            .I(\RSMRST_PWRGD.un1_count_1_cry_6 ));
    InMux I__1411 (
            .O(N__14267),
            .I(N__14263));
    InMux I__1410 (
            .O(N__14266),
            .I(N__14260));
    LocalMux I__1409 (
            .O(N__14263),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    LocalMux I__1408 (
            .O(N__14260),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    InMux I__1407 (
            .O(N__14255),
            .I(bfn_2_2_0_));
    InMux I__1406 (
            .O(N__14252),
            .I(N__14248));
    InMux I__1405 (
            .O(N__14251),
            .I(N__14245));
    LocalMux I__1404 (
            .O(N__14248),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    LocalMux I__1403 (
            .O(N__14245),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    InMux I__1402 (
            .O(N__14240),
            .I(\RSMRST_PWRGD.un1_count_1_cry_8 ));
    InMux I__1401 (
            .O(N__14237),
            .I(N__14233));
    InMux I__1400 (
            .O(N__14236),
            .I(N__14230));
    LocalMux I__1399 (
            .O(N__14233),
            .I(N__14227));
    LocalMux I__1398 (
            .O(N__14230),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    Odrv4 I__1397 (
            .O(N__14227),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    InMux I__1396 (
            .O(N__14222),
            .I(\RSMRST_PWRGD.un1_count_1_cry_9 ));
    InMux I__1395 (
            .O(N__14219),
            .I(N__14215));
    InMux I__1394 (
            .O(N__14218),
            .I(N__14212));
    LocalMux I__1393 (
            .O(N__14215),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    LocalMux I__1392 (
            .O(N__14212),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    InMux I__1391 (
            .O(N__14207),
            .I(\RSMRST_PWRGD.un1_count_1_cry_10 ));
    CascadeMux I__1390 (
            .O(N__14204),
            .I(\POWERLED.N_660_cascade_ ));
    InMux I__1389 (
            .O(N__14201),
            .I(N__14177));
    InMux I__1388 (
            .O(N__14200),
            .I(N__14177));
    InMux I__1387 (
            .O(N__14199),
            .I(N__14177));
    InMux I__1386 (
            .O(N__14198),
            .I(N__14168));
    InMux I__1385 (
            .O(N__14197),
            .I(N__14168));
    InMux I__1384 (
            .O(N__14196),
            .I(N__14168));
    InMux I__1383 (
            .O(N__14195),
            .I(N__14168));
    InMux I__1382 (
            .O(N__14194),
            .I(N__14159));
    InMux I__1381 (
            .O(N__14193),
            .I(N__14159));
    InMux I__1380 (
            .O(N__14192),
            .I(N__14159));
    InMux I__1379 (
            .O(N__14191),
            .I(N__14159));
    InMux I__1378 (
            .O(N__14190),
            .I(N__14150));
    InMux I__1377 (
            .O(N__14189),
            .I(N__14150));
    InMux I__1376 (
            .O(N__14188),
            .I(N__14150));
    InMux I__1375 (
            .O(N__14187),
            .I(N__14150));
    InMux I__1374 (
            .O(N__14186),
            .I(N__14143));
    InMux I__1373 (
            .O(N__14185),
            .I(N__14143));
    InMux I__1372 (
            .O(N__14184),
            .I(N__14143));
    LocalMux I__1371 (
            .O(N__14177),
            .I(N__14140));
    LocalMux I__1370 (
            .O(N__14168),
            .I(N__14137));
    LocalMux I__1369 (
            .O(N__14159),
            .I(N__14134));
    LocalMux I__1368 (
            .O(N__14150),
            .I(\POWERLED.count_0_sqmuxa_i ));
    LocalMux I__1367 (
            .O(N__14143),
            .I(\POWERLED.count_0_sqmuxa_i ));
    Odrv4 I__1366 (
            .O(N__14140),
            .I(\POWERLED.count_0_sqmuxa_i ));
    Odrv4 I__1365 (
            .O(N__14137),
            .I(\POWERLED.count_0_sqmuxa_i ));
    Odrv12 I__1364 (
            .O(N__14134),
            .I(\POWERLED.count_0_sqmuxa_i ));
    InMux I__1363 (
            .O(N__14123),
            .I(N__14120));
    LocalMux I__1362 (
            .O(N__14120),
            .I(\POWERLED.pwm_out_1_sqmuxa_0 ));
    CascadeMux I__1361 (
            .O(N__14117),
            .I(\POWERLED.pwm_out_en_cascade_ ));
    InMux I__1360 (
            .O(N__14114),
            .I(N__14110));
    InMux I__1359 (
            .O(N__14113),
            .I(N__14107));
    LocalMux I__1358 (
            .O(N__14110),
            .I(\POWERLED.pwm_outZ0 ));
    LocalMux I__1357 (
            .O(N__14107),
            .I(\POWERLED.pwm_outZ0 ));
    IoInMux I__1356 (
            .O(N__14102),
            .I(N__14099));
    LocalMux I__1355 (
            .O(N__14099),
            .I(N__14096));
    Odrv4 I__1354 (
            .O(N__14096),
            .I(pwrbtn_led));
    InMux I__1353 (
            .O(N__14093),
            .I(N__14090));
    LocalMux I__1352 (
            .O(N__14090),
            .I(N__14087));
    Span4Mux_s3_v I__1351 (
            .O(N__14087),
            .I(N__14084));
    Odrv4 I__1350 (
            .O(N__14084),
            .I(vpp_ok));
    IoInMux I__1349 (
            .O(N__14081),
            .I(N__14078));
    LocalMux I__1348 (
            .O(N__14078),
            .I(N__14075));
    Odrv4 I__1347 (
            .O(N__14075),
            .I(vddq_en));
    InMux I__1346 (
            .O(N__14072),
            .I(N__14068));
    InMux I__1345 (
            .O(N__14071),
            .I(N__14065));
    LocalMux I__1344 (
            .O(N__14068),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    LocalMux I__1343 (
            .O(N__14065),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    InMux I__1342 (
            .O(N__14060),
            .I(N__14056));
    InMux I__1341 (
            .O(N__14059),
            .I(N__14053));
    LocalMux I__1340 (
            .O(N__14056),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    LocalMux I__1339 (
            .O(N__14053),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    InMux I__1338 (
            .O(N__14048),
            .I(\RSMRST_PWRGD.un1_count_1_cry_0 ));
    CascadeMux I__1337 (
            .O(N__14045),
            .I(N__14041));
    InMux I__1336 (
            .O(N__14044),
            .I(N__14038));
    InMux I__1335 (
            .O(N__14041),
            .I(N__14035));
    LocalMux I__1334 (
            .O(N__14038),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    LocalMux I__1333 (
            .O(N__14035),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    InMux I__1332 (
            .O(N__14030),
            .I(\RSMRST_PWRGD.un1_count_1_cry_1 ));
    InMux I__1331 (
            .O(N__14027),
            .I(\POWERLED.un1_count_cry_11 ));
    InMux I__1330 (
            .O(N__14024),
            .I(\POWERLED.un1_count_cry_12 ));
    InMux I__1329 (
            .O(N__14021),
            .I(\POWERLED.un1_count_cry_13 ));
    InMux I__1328 (
            .O(N__14018),
            .I(\POWERLED.un1_count_cry_14 ));
    InMux I__1327 (
            .O(N__14015),
            .I(N__14011));
    InMux I__1326 (
            .O(N__14014),
            .I(N__14008));
    LocalMux I__1325 (
            .O(N__14011),
            .I(N__14005));
    LocalMux I__1324 (
            .O(N__14008),
            .I(\POWERLED.count_1_12 ));
    Odrv4 I__1323 (
            .O(N__14005),
            .I(\POWERLED.count_1_12 ));
    InMux I__1322 (
            .O(N__14000),
            .I(N__13997));
    LocalMux I__1321 (
            .O(N__13997),
            .I(N__13994));
    Odrv12 I__1320 (
            .O(N__13994),
            .I(\POWERLED.count_0_12 ));
    CascadeMux I__1319 (
            .O(N__13991),
            .I(\POWERLED.N_437_cascade_ ));
    CascadeMux I__1318 (
            .O(N__13988),
            .I(\POWERLED.N_2305_i_cascade_ ));
    InMux I__1317 (
            .O(N__13985),
            .I(N__13979));
    InMux I__1316 (
            .O(N__13984),
            .I(N__13979));
    LocalMux I__1315 (
            .O(N__13979),
            .I(N__13976));
    Odrv4 I__1314 (
            .O(N__13976),
            .I(\POWERLED.count_1_3 ));
    InMux I__1313 (
            .O(N__13973),
            .I(\POWERLED.un1_count_cry_2_cZ0 ));
    InMux I__1312 (
            .O(N__13970),
            .I(N__13964));
    InMux I__1311 (
            .O(N__13969),
            .I(N__13964));
    LocalMux I__1310 (
            .O(N__13964),
            .I(\POWERLED.count_1_4 ));
    InMux I__1309 (
            .O(N__13961),
            .I(\POWERLED.un1_count_cry_3_cZ0 ));
    InMux I__1308 (
            .O(N__13958),
            .I(\POWERLED.un1_count_cry_4_cZ0 ));
    InMux I__1307 (
            .O(N__13955),
            .I(\POWERLED.un1_count_cry_5 ));
    InMux I__1306 (
            .O(N__13952),
            .I(\POWERLED.un1_count_cry_6 ));
    InMux I__1305 (
            .O(N__13949),
            .I(\POWERLED.un1_count_cry_7 ));
    InMux I__1304 (
            .O(N__13946),
            .I(bfn_1_12_0_));
    InMux I__1303 (
            .O(N__13943),
            .I(\POWERLED.un1_count_cry_9 ));
    CascadeMux I__1302 (
            .O(N__13940),
            .I(N__13937));
    InMux I__1301 (
            .O(N__13937),
            .I(N__13931));
    InMux I__1300 (
            .O(N__13936),
            .I(N__13931));
    LocalMux I__1299 (
            .O(N__13931),
            .I(N__13928));
    Odrv4 I__1298 (
            .O(N__13928),
            .I(\POWERLED.count_1_11 ));
    InMux I__1297 (
            .O(N__13925),
            .I(\POWERLED.un1_count_cry_10 ));
    InMux I__1296 (
            .O(N__13922),
            .I(N__13919));
    LocalMux I__1295 (
            .O(N__13919),
            .I(\POWERLED.count_0_0 ));
    CascadeMux I__1294 (
            .O(N__13916),
            .I(\POWERLED.count_1_0_cascade_ ));
    CascadeMux I__1293 (
            .O(N__13913),
            .I(\POWERLED.countZ0Z_0_cascade_ ));
    CascadeMux I__1292 (
            .O(N__13910),
            .I(\POWERLED.count_1_1_cascade_ ));
    CascadeMux I__1291 (
            .O(N__13907),
            .I(\POWERLED.countZ0Z_1_cascade_ ));
    InMux I__1290 (
            .O(N__13904),
            .I(N__13901));
    LocalMux I__1289 (
            .O(N__13901),
            .I(\POWERLED.count_0_1 ));
    InMux I__1288 (
            .O(N__13898),
            .I(N__13895));
    LocalMux I__1287 (
            .O(N__13895),
            .I(\POWERLED.count_0_4 ));
    InMux I__1286 (
            .O(N__13892),
            .I(N__13886));
    InMux I__1285 (
            .O(N__13891),
            .I(N__13886));
    LocalMux I__1284 (
            .O(N__13886),
            .I(N__13883));
    Odrv4 I__1283 (
            .O(N__13883),
            .I(\POWERLED.count_1_2 ));
    InMux I__1282 (
            .O(N__13880),
            .I(\POWERLED.un1_count_cry_1 ));
    InMux I__1281 (
            .O(N__13877),
            .I(N__13874));
    LocalMux I__1280 (
            .O(N__13874),
            .I(\POWERLED.count_0_2 ));
    IoInMux I__1279 (
            .O(N__13871),
            .I(N__13868));
    LocalMux I__1278 (
            .O(N__13868),
            .I(G_12));
    InMux I__1277 (
            .O(N__13865),
            .I(N__13862));
    LocalMux I__1276 (
            .O(N__13862),
            .I(\POWERLED.count_0_11 ));
    InMux I__1275 (
            .O(N__13859),
            .I(N__13856));
    LocalMux I__1274 (
            .O(N__13856),
            .I(\POWERLED.count_0_3 ));
    InMux I__1273 (
            .O(N__13853),
            .I(N__13850));
    LocalMux I__1272 (
            .O(N__13850),
            .I(\PCH_PWRGD.count_0_6 ));
    CascadeMux I__1271 (
            .O(N__13847),
            .I(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0_cascade_ ));
    InMux I__1270 (
            .O(N__13844),
            .I(N__13838));
    InMux I__1269 (
            .O(N__13843),
            .I(N__13838));
    LocalMux I__1268 (
            .O(N__13838),
            .I(N__13835));
    Odrv4 I__1267 (
            .O(N__13835),
            .I(\PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0 ));
    CascadeMux I__1266 (
            .O(N__13832),
            .I(\PCH_PWRGD.un2_count_1_axb_1_cascade_ ));
    CascadeMux I__1265 (
            .O(N__13829),
            .I(\PCH_PWRGD.N_2284_i_cascade_ ));
    CascadeMux I__1264 (
            .O(N__13826),
            .I(\PCH_PWRGD.N_655_cascade_ ));
    CascadeMux I__1263 (
            .O(N__13823),
            .I(\PCH_PWRGD.count_0_sqmuxa_cascade_ ));
    InMux I__1262 (
            .O(N__13820),
            .I(N__13816));
    InMux I__1261 (
            .O(N__13819),
            .I(N__13813));
    LocalMux I__1260 (
            .O(N__13816),
            .I(N__13810));
    LocalMux I__1259 (
            .O(N__13813),
            .I(\PCH_PWRGD.un2_count_1_axb_1 ));
    Odrv4 I__1258 (
            .O(N__13810),
            .I(\PCH_PWRGD.un2_count_1_axb_1 ));
    InMux I__1257 (
            .O(N__13805),
            .I(N__13799));
    InMux I__1256 (
            .O(N__13804),
            .I(N__13799));
    LocalMux I__1255 (
            .O(N__13799),
            .I(\PCH_PWRGD.count_0_1 ));
    CascadeMux I__1254 (
            .O(N__13796),
            .I(N__13793));
    InMux I__1253 (
            .O(N__13793),
            .I(N__13787));
    InMux I__1252 (
            .O(N__13792),
            .I(N__13787));
    LocalMux I__1251 (
            .O(N__13787),
            .I(\PCH_PWRGD.count_rst_13 ));
    InMux I__1250 (
            .O(N__13784),
            .I(N__13780));
    InMux I__1249 (
            .O(N__13783),
            .I(N__13777));
    LocalMux I__1248 (
            .O(N__13780),
            .I(vr_ready_vccin));
    LocalMux I__1247 (
            .O(N__13777),
            .I(vr_ready_vccin));
    InMux I__1246 (
            .O(N__13772),
            .I(N__13769));
    LocalMux I__1245 (
            .O(N__13769),
            .I(\PCH_PWRGD.N_2284_i ));
    InMux I__1244 (
            .O(N__13766),
            .I(\PCH_PWRGD.un2_count_1_cry_13 ));
    InMux I__1243 (
            .O(N__13763),
            .I(\PCH_PWRGD.un2_count_1_cry_14 ));
    InMux I__1242 (
            .O(N__13760),
            .I(N__13757));
    LocalMux I__1241 (
            .O(N__13757),
            .I(N__13754));
    Odrv4 I__1240 (
            .O(N__13754),
            .I(\PCH_PWRGD.un2_count_1_axb_2 ));
    InMux I__1239 (
            .O(N__13751),
            .I(N__13744));
    InMux I__1238 (
            .O(N__13750),
            .I(N__13744));
    InMux I__1237 (
            .O(N__13749),
            .I(N__13741));
    LocalMux I__1236 (
            .O(N__13744),
            .I(N__13738));
    LocalMux I__1235 (
            .O(N__13741),
            .I(\PCH_PWRGD.count_rst_12 ));
    Odrv4 I__1234 (
            .O(N__13738),
            .I(\PCH_PWRGD.count_rst_12 ));
    InMux I__1233 (
            .O(N__13733),
            .I(N__13729));
    InMux I__1232 (
            .O(N__13732),
            .I(N__13726));
    LocalMux I__1231 (
            .O(N__13729),
            .I(\PCH_PWRGD.count_0_2 ));
    LocalMux I__1230 (
            .O(N__13726),
            .I(\PCH_PWRGD.count_0_2 ));
    InMux I__1229 (
            .O(N__13721),
            .I(N__13718));
    LocalMux I__1228 (
            .O(N__13718),
            .I(\PCH_PWRGD.count_0_14 ));
    CascadeMux I__1227 (
            .O(N__13715),
            .I(N__13711));
    InMux I__1226 (
            .O(N__13714),
            .I(N__13706));
    InMux I__1225 (
            .O(N__13711),
            .I(N__13706));
    LocalMux I__1224 (
            .O(N__13706),
            .I(\PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7 ));
    InMux I__1223 (
            .O(N__13703),
            .I(N__13697));
    InMux I__1222 (
            .O(N__13702),
            .I(N__13697));
    LocalMux I__1221 (
            .O(N__13697),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    InMux I__1220 (
            .O(N__13694),
            .I(\PCH_PWRGD.un2_count_1_cry_4 ));
    InMux I__1219 (
            .O(N__13691),
            .I(\PCH_PWRGD.un2_count_1_cry_5 ));
    InMux I__1218 (
            .O(N__13688),
            .I(\PCH_PWRGD.un2_count_1_cry_6 ));
    InMux I__1217 (
            .O(N__13685),
            .I(N__13680));
    InMux I__1216 (
            .O(N__13684),
            .I(N__13677));
    InMux I__1215 (
            .O(N__13683),
            .I(N__13674));
    LocalMux I__1214 (
            .O(N__13680),
            .I(N__13671));
    LocalMux I__1213 (
            .O(N__13677),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    LocalMux I__1212 (
            .O(N__13674),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    Odrv4 I__1211 (
            .O(N__13671),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    CascadeMux I__1210 (
            .O(N__13664),
            .I(N__13660));
    CascadeMux I__1209 (
            .O(N__13663),
            .I(N__13657));
    InMux I__1208 (
            .O(N__13660),
            .I(N__13654));
    InMux I__1207 (
            .O(N__13657),
            .I(N__13651));
    LocalMux I__1206 (
            .O(N__13654),
            .I(N__13646));
    LocalMux I__1205 (
            .O(N__13651),
            .I(N__13646));
    Span4Mux_s2_v I__1204 (
            .O(N__13646),
            .I(N__13643));
    Odrv4 I__1203 (
            .O(N__13643),
            .I(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ));
    InMux I__1202 (
            .O(N__13640),
            .I(\PCH_PWRGD.un2_count_1_cry_7 ));
    CascadeMux I__1201 (
            .O(N__13637),
            .I(N__13634));
    InMux I__1200 (
            .O(N__13634),
            .I(N__13630));
    InMux I__1199 (
            .O(N__13633),
            .I(N__13627));
    LocalMux I__1198 (
            .O(N__13630),
            .I(N__13624));
    LocalMux I__1197 (
            .O(N__13627),
            .I(N__13621));
    Odrv4 I__1196 (
            .O(N__13624),
            .I(\PCH_PWRGD.un2_count_1_axb_9 ));
    Odrv4 I__1195 (
            .O(N__13621),
            .I(\PCH_PWRGD.un2_count_1_axb_9 ));
    InMux I__1194 (
            .O(N__13616),
            .I(N__13610));
    InMux I__1193 (
            .O(N__13615),
            .I(N__13610));
    LocalMux I__1192 (
            .O(N__13610),
            .I(N__13607));
    Odrv4 I__1191 (
            .O(N__13607),
            .I(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ));
    InMux I__1190 (
            .O(N__13604),
            .I(bfn_1_6_0_));
    InMux I__1189 (
            .O(N__13601),
            .I(\PCH_PWRGD.un2_count_1_cry_9 ));
    InMux I__1188 (
            .O(N__13598),
            .I(\PCH_PWRGD.un2_count_1_cry_10 ));
    InMux I__1187 (
            .O(N__13595),
            .I(\PCH_PWRGD.un2_count_1_cry_11 ));
    InMux I__1186 (
            .O(N__13592),
            .I(\PCH_PWRGD.un2_count_1_cry_12 ));
    CascadeMux I__1185 (
            .O(N__13589),
            .I(\PCH_PWRGD.un2_count_1_axb_4_cascade_ ));
    InMux I__1184 (
            .O(N__13586),
            .I(N__13583));
    LocalMux I__1183 (
            .O(N__13583),
            .I(\PCH_PWRGD.count_0_3 ));
    InMux I__1182 (
            .O(N__13580),
            .I(N__13577));
    LocalMux I__1181 (
            .O(N__13577),
            .I(\PCH_PWRGD.count_rst_10 ));
    InMux I__1180 (
            .O(N__13574),
            .I(N__13568));
    InMux I__1179 (
            .O(N__13573),
            .I(N__13568));
    LocalMux I__1178 (
            .O(N__13568),
            .I(N__13565));
    Odrv4 I__1177 (
            .O(N__13565),
            .I(\PCH_PWRGD.count_0_4 ));
    CascadeMux I__1176 (
            .O(N__13562),
            .I(\PCH_PWRGD.count_rst_10_cascade_ ));
    InMux I__1175 (
            .O(N__13559),
            .I(\PCH_PWRGD.un2_count_1_cry_1 ));
    InMux I__1174 (
            .O(N__13556),
            .I(N__13548));
    InMux I__1173 (
            .O(N__13555),
            .I(N__13548));
    InMux I__1172 (
            .O(N__13554),
            .I(N__13545));
    InMux I__1171 (
            .O(N__13553),
            .I(N__13542));
    LocalMux I__1170 (
            .O(N__13548),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    LocalMux I__1169 (
            .O(N__13545),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    LocalMux I__1168 (
            .O(N__13542),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    CascadeMux I__1167 (
            .O(N__13535),
            .I(N__13531));
    CascadeMux I__1166 (
            .O(N__13534),
            .I(N__13528));
    InMux I__1165 (
            .O(N__13531),
            .I(N__13523));
    InMux I__1164 (
            .O(N__13528),
            .I(N__13523));
    LocalMux I__1163 (
            .O(N__13523),
            .I(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ));
    InMux I__1162 (
            .O(N__13520),
            .I(\PCH_PWRGD.un2_count_1_cry_2 ));
    InMux I__1161 (
            .O(N__13517),
            .I(N__13513));
    InMux I__1160 (
            .O(N__13516),
            .I(N__13510));
    LocalMux I__1159 (
            .O(N__13513),
            .I(\PCH_PWRGD.un2_count_1_axb_4 ));
    LocalMux I__1158 (
            .O(N__13510),
            .I(\PCH_PWRGD.un2_count_1_axb_4 ));
    InMux I__1157 (
            .O(N__13505),
            .I(N__13499));
    InMux I__1156 (
            .O(N__13504),
            .I(N__13499));
    LocalMux I__1155 (
            .O(N__13499),
            .I(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ));
    InMux I__1154 (
            .O(N__13496),
            .I(\PCH_PWRGD.un2_count_1_cry_3 ));
    CascadeMux I__1153 (
            .O(N__13493),
            .I(\PCH_PWRGD.count_rst_5_cascade_ ));
    CascadeMux I__1152 (
            .O(N__13490),
            .I(\PCH_PWRGD.un2_count_1_axb_9_cascade_ ));
    InMux I__1151 (
            .O(N__13487),
            .I(N__13484));
    LocalMux I__1150 (
            .O(N__13484),
            .I(\PCH_PWRGD.count_0_8 ));
    CascadeMux I__1149 (
            .O(N__13481),
            .I(\PCH_PWRGD.count_rst_6_cascade_ ));
    InMux I__1148 (
            .O(N__13478),
            .I(N__13472));
    InMux I__1147 (
            .O(N__13477),
            .I(N__13472));
    LocalMux I__1146 (
            .O(N__13472),
            .I(\PCH_PWRGD.count_0_9 ));
    CascadeMux I__1145 (
            .O(N__13469),
            .I(\PCH_PWRGD.countZ0Z_8_cascade_ ));
    InMux I__1144 (
            .O(N__13466),
            .I(N__13463));
    LocalMux I__1143 (
            .O(N__13463),
            .I(\PCH_PWRGD.count_rst_5 ));
    CascadeMux I__1142 (
            .O(N__13460),
            .I(\PCH_PWRGD.count_rst_11_cascade_ ));
    CascadeMux I__1141 (
            .O(N__13457),
            .I(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_10_cascade_ ));
    InMux I__1140 (
            .O(N__13454),
            .I(N__13451));
    LocalMux I__1139 (
            .O(N__13451),
            .I(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_11 ));
    CascadeMux I__1138 (
            .O(N__13448),
            .I(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_0_cascade_ ));
    InMux I__1137 (
            .O(N__13445),
            .I(N__13442));
    LocalMux I__1136 (
            .O(N__13442),
            .I(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_12 ));
    InMux I__1135 (
            .O(N__13439),
            .I(N__13436));
    LocalMux I__1134 (
            .O(N__13436),
            .I(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_9 ));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_7_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_3_0_));
    defparam IN_MUX_bfv_7_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_4_0_ (
            .carryinitin(\POWERLED.un3_count_off_1_cry_8 ),
            .carryinitout(bfn_7_4_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_6_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_16_0_));
    defparam IN_MUX_bfv_6_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_15_0_));
    defparam IN_MUX_bfv_6_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_14_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_6_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_12_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_4_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_10_0_));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_11_0_));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\POWERLED.un1_count_cry_8 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_12_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_5_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_1_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_5_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(\PCH_PWRGD.un2_count_1_cry_8 ),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_5_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_1_0_));
    defparam IN_MUX_bfv_5_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_2_0_ (
            .carryinitin(\HDA_STRAP.un1_count_1_cry_7 ),
            .carryinitout(bfn_5_2_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(\HDA_STRAP.un1_count_1_cry_15 ),
            .carryinitout(bfn_5_3_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(COUNTER_un4_counter_7),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(\COUNTER.counter_1_cry_8 ),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(\COUNTER.counter_1_cry_16 ),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(\COUNTER.counter_1_cry_24 ),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_11_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_2_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_7 ),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_11_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_4_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_11_4_0_));
    defparam IN_MUX_bfv_2_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_1_0_));
    defparam IN_MUX_bfv_2_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_2_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_2_2_0_));
    defparam IN_MUX_bfv_2_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_3_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_2_3_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_4_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_15_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_7 ),
            .carryinitout(bfn_4_15_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_94_cry_7_cZ0 ),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_7 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_15 ),
            .carryinitout(bfn_7_15_0_));
    ICE_GB N_92_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__13871),
            .GLOBALBUFFEROUTPUT(N_92_g));
    ICE_GB N_557_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__32674),
            .GLOBALBUFFEROUTPUT(N_557_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI4MLK1_1_LC_1_1_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI4MLK1_1_LC_1_1_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI4MLK1_1_LC_1_1_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.count_RNI4MLK1_1_LC_1_1_0  (
            .in0(N__14251),
            .in1(N__14332),
            .in2(N__14045),
            .in3(N__14059),
            .lcout(),
            .ltout(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIST215_10_LC_1_1_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIST215_10_LC_1_1_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIST215_10_LC_1_1_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIST215_10_LC_1_1_1  (
            .in0(N__13454),
            .in1(N__13439),
            .in2(N__13457),
            .in3(N__13445),
            .lcout(N_662),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIMVQE1_3_LC_1_1_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIMVQE1_3_LC_1_1_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIMVQE1_3_LC_1_1_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIMVQE1_3_LC_1_1_2  (
            .in0(N__21173),
            .in1(N__14347),
            .in2(N__14318),
            .in3(N__14296),
            .lcout(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIVSS4_11_LC_1_1_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIVSS4_11_LC_1_1_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIVSS4_11_LC_1_1_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIVSS4_11_LC_1_1_3  (
            .in0(_gnd_net_),
            .in1(N__14443),
            .in2(_gnd_net_),
            .in3(N__14218),
            .lcout(),
            .ltout(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI6CM11_10_LC_1_1_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI6CM11_10_LC_1_1_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI6CM11_10_LC_1_1_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNI6CM11_10_LC_1_1_4  (
            .in0(N__14237),
            .in1(N__14266),
            .in2(N__13448),
            .in3(N__14281),
            .lcout(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_RNISRRR_15_LC_1_1_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_RNISRRR_15_LC_1_1_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_esr_RNISRRR_15_LC_1_1_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \RSMRST_PWRGD.count_esr_RNISRRR_15_LC_1_1_5  (
            .in0(N__14428),
            .in1(N__14413),
            .in2(N__14396),
            .in3(N__14071),
            .lcout(\RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_8_LC_1_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_8_LC_1_2_2 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_8_LC_1_2_2 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \PCH_PWRGD.count_8_LC_1_2_2  (
            .in0(N__15351),
            .in1(N__14940),
            .in2(N__13664),
            .in3(N__13683),
            .lcout(\PCH_PWRGD.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32317),
            .ce(N__15138),
            .sr(N__14941));
    defparam \PCH_PWRGD.count_11_LC_1_3_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_11_LC_1_3_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_11_LC_1_3_0 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \PCH_PWRGD.count_11_LC_1_3_0  (
            .in0(N__14937),
            .in1(N__15355),
            .in2(N__14508),
            .in3(N__14539),
            .lcout(\PCH_PWRGD.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32355),
            .ce(N__15132),
            .sr(N__14965));
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIQKDU1_LC_1_3_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIQKDU1_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIQKDU1_LC_1_3_2 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_c_RNIQKDU1_LC_1_3_2  (
            .in0(N__14936),
            .in1(N__13615),
            .in2(N__13637),
            .in3(N__15354),
            .lcout(\PCH_PWRGD.count_rst_5 ),
            .ltout(\PCH_PWRGD.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI27DA2_9_LC_1_3_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI27DA2_9_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI27DA2_9_LC_1_3_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNI27DA2_9_LC_1_3_3  (
            .in0(N__15068),
            .in1(_gnd_net_),
            .in2(N__13493),
            .in3(N__13477),
            .lcout(\PCH_PWRGD.un2_count_1_axb_9 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_9_LC_1_3_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_9_LC_1_3_4 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_9_LC_1_3_4 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \PCH_PWRGD.count_9_LC_1_3_4  (
            .in0(N__14938),
            .in1(N__15356),
            .in2(N__13490),
            .in3(N__13616),
            .lcout(\PCH_PWRGD.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32355),
            .ce(N__15132),
            .sr(N__14965));
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIPICU1_LC_1_3_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIPICU1_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIPICU1_LC_1_3_5 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_c_RNIPICU1_LC_1_3_5  (
            .in0(N__15353),
            .in1(N__14935),
            .in2(N__13663),
            .in3(N__13684),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIQOP84_8_LC_1_3_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQOP84_8_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQOP84_8_LC_1_3_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.count_RNIQOP84_8_LC_1_3_6  (
            .in0(_gnd_net_),
            .in1(N__13487),
            .in2(N__13481),
            .in3(N__15067),
            .lcout(\PCH_PWRGD.countZ0Z_8 ),
            .ltout(\PCH_PWRGD.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI27DA2_0_9_LC_1_3_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI27DA2_0_9_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI27DA2_0_9_LC_1_3_7 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \PCH_PWRGD.count_RNI27DA2_0_9_LC_1_3_7  (
            .in0(N__15069),
            .in1(N__13478),
            .in2(N__13469),
            .in3(N__13466),
            .lcout(\PCH_PWRGD.count_1_i_a2_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNIK87U1_LC_1_4_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNIK87U1_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNIK87U1_LC_1_4_0 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_c_RNIK87U1_LC_1_4_0  (
            .in0(N__13556),
            .in1(N__15319),
            .in2(N__13534),
            .in3(N__14931),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIG9K84_3_LC_1_4_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIG9K84_3_LC_1_4_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIG9K84_3_LC_1_4_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNIG9K84_3_LC_1_4_1  (
            .in0(N__15064),
            .in1(_gnd_net_),
            .in2(N__13460),
            .in3(N__13586),
            .lcout(\PCH_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIT1DA2_4_LC_1_4_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIT1DA2_4_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIT1DA2_4_LC_1_4_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \PCH_PWRGD.count_RNIT1DA2_4_LC_1_4_2  (
            .in0(N__13573),
            .in1(N__15065),
            .in2(_gnd_net_),
            .in3(N__13580),
            .lcout(\PCH_PWRGD.un2_count_1_axb_4 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_4_LC_1_4_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_4_LC_1_4_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_4_LC_1_4_3 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \PCH_PWRGD.count_4_LC_1_4_3  (
            .in0(N__15324),
            .in1(N__14960),
            .in2(N__13589),
            .in3(N__13505),
            .lcout(\PCH_PWRGD.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32335),
            .ce(N__15070),
            .sr(N__14966));
    defparam \PCH_PWRGD.count_3_LC_1_4_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_3_LC_1_4_4 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_3_LC_1_4_4 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \PCH_PWRGD.count_3_LC_1_4_4  (
            .in0(N__13555),
            .in1(N__15323),
            .in2(N__13535),
            .in3(N__14934),
            .lcout(\PCH_PWRGD.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32335),
            .ce(N__15070),
            .sr(N__14966));
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNILA8U1_LC_1_4_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNILA8U1_LC_1_4_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNILA8U1_LC_1_4_5 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_c_RNILA8U1_LC_1_4_5  (
            .in0(N__14932),
            .in1(N__13517),
            .in2(N__15349),
            .in3(N__13504),
            .lcout(\PCH_PWRGD.count_rst_10 ),
            .ltout(\PCH_PWRGD.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIT1DA2_0_4_LC_1_4_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIT1DA2_0_4_LC_1_4_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIT1DA2_0_4_LC_1_4_6 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \PCH_PWRGD.count_RNIT1DA2_0_4_LC_1_4_6  (
            .in0(N__13574),
            .in1(N__15066),
            .in2(N__13562),
            .in3(N__13554),
            .lcout(\PCH_PWRGD.count_1_i_a2_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_5_LC_1_4_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_5_LC_1_4_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_5_LC_1_4_7 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \PCH_PWRGD.count_5_LC_1_4_7  (
            .in0(N__14933),
            .in1(N__14748),
            .in2(N__15350),
            .in3(N__14360),
            .lcout(\PCH_PWRGD.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32335),
            .ce(N__15070),
            .sr(N__14966));
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_5_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(N__13820),
            .in2(N__14674),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_5_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNIJ66U1_LC_1_5_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNIJ66U1_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNIJ66U1_LC_1_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_1_c_RNIJ66U1_LC_1_5_1  (
            .in0(N__14917),
            .in1(N__13760),
            .in2(_gnd_net_),
            .in3(N__13559),
            .lcout(\PCH_PWRGD.count_rst_12 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_1 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_5_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_5_2  (
            .in0(_gnd_net_),
            .in1(N__13553),
            .in2(_gnd_net_),
            .in3(N__13520),
            .lcout(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_2 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_5_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_5_3  (
            .in0(_gnd_net_),
            .in1(N__13516),
            .in2(_gnd_net_),
            .in3(N__13496),
            .lcout(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_3 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_5_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(N__14738),
            .in2(_gnd_net_),
            .in3(N__13694),
            .lcout(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_4 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_1_5_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_1_5_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14603),
            .in3(N__13691),
            .lcout(\PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_5 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_5_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_5_6  (
            .in0(_gnd_net_),
            .in1(N__14473),
            .in2(_gnd_net_),
            .in3(N__13688),
            .lcout(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_6 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_5_7 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_5_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(N__13685),
            .in2(_gnd_net_),
            .in3(N__13640),
            .lcout(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_7 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_6_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__13633),
            .in2(_gnd_net_),
            .in3(N__13604),
            .lcout(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIRMEU1_LC_1_6_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIRMEU1_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIRMEU1_LC_1_6_1 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_9_c_RNIRMEU1_LC_1_6_1  (
            .in0(N__14926),
            .in1(_gnd_net_),
            .in2(N__14552),
            .in3(N__13601),
            .lcout(\PCH_PWRGD.count_rst_4 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_9 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_6_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(N__14510),
            .in2(_gnd_net_),
            .in3(N__13598),
            .lcout(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_10 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNI402P1_LC_1_6_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNI402P1_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNI402P1_LC_1_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_11_c_RNI402P1_LC_1_6_3  (
            .in0(N__14927),
            .in1(N__14584),
            .in2(_gnd_net_),
            .in3(N__13595),
            .lcout(\PCH_PWRGD.count_rst_2 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_11 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNI523P1_LC_1_6_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNI523P1_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNI523P1_LC_1_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_12_c_RNI523P1_LC_1_6_4  (
            .in0(N__14939),
            .in1(N__14609),
            .in2(_gnd_net_),
            .in3(N__13592),
            .lcout(\PCH_PWRGD.count_rst_1 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_12 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_1_6_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_1_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(N__13702),
            .in2(_gnd_net_),
            .in3(N__13766),
            .lcout(\PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_13 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNI765P1_LC_1_6_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNI765P1_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNI765P1_LC_1_6_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_14_c_RNI765P1_LC_1_6_6  (
            .in0(N__14621),
            .in1(N__14928),
            .in2(_gnd_net_),
            .in3(N__13763),
            .lcout(\PCH_PWRGD.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIE6J84_0_2_LC_1_6_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIE6J84_0_2_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIE6J84_0_2_LC_1_6_7 .LUT_INIT=16'b0000000001010011;
    LogicCell40 \PCH_PWRGD.count_RNIE6J84_0_2_LC_1_6_7  (
            .in0(N__13749),
            .in1(N__13733),
            .in2(N__15098),
            .in3(N__13703),
            .lcout(\PCH_PWRGD.count_1_i_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_6_LC_1_7_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_6_LC_1_7_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_6_LC_1_7_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \PCH_PWRGD.count_6_LC_1_7_0  (
            .in0(N__13843),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14849),
            .lcout(\PCH_PWRGD.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32401),
            .ce(N__15140),
            .sr(N__14916));
    defparam \PCH_PWRGD.count_RNIE6J84_2_LC_1_7_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIE6J84_2_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIE6J84_2_LC_1_7_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \PCH_PWRGD.count_RNIE6J84_2_LC_1_7_1  (
            .in0(N__13732),
            .in1(N__15017),
            .in2(_gnd_net_),
            .in3(N__13750),
            .lcout(\PCH_PWRGD.un2_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_2_LC_1_7_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_2_LC_1_7_2 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_2_LC_1_7_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_2_LC_1_7_2  (
            .in0(N__13751),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32401),
            .ce(N__15140),
            .sr(N__14916));
    defparam \PCH_PWRGD.count_14_LC_1_7_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_14_LC_1_7_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_14_LC_1_7_3 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \PCH_PWRGD.count_14_LC_1_7_3  (
            .in0(N__14848),
            .in1(N__13714),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32401),
            .ce(N__15140),
            .sr(N__14916));
    defparam \PCH_PWRGD.count_RNIKP0C4_14_LC_1_7_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIKP0C4_14_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIKP0C4_14_LC_1_7_4 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \PCH_PWRGD.count_RNIKP0C4_14_LC_1_7_4  (
            .in0(N__15018),
            .in1(N__13721),
            .in2(N__13715),
            .in3(N__14847),
            .lcout(\PCH_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNISDK72_0_LC_1_7_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNISDK72_0_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNISDK72_0_LC_1_7_6 .LUT_INIT=16'b1100110100000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNISDK72_0_LC_1_7_6  (
            .in0(N__15407),
            .in1(N__14846),
            .in2(N__15862),
            .in3(N__32675),
            .lcout(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0 ),
            .ltout(\PCH_PWRGD.curr_state_RNISDK72Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIMIN84_6_LC_1_7_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIMIN84_6_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIMIN84_6_LC_1_7_7 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \PCH_PWRGD.count_RNIMIN84_6_LC_1_7_7  (
            .in0(N__14850),
            .in1(N__13853),
            .in2(N__13847),
            .in3(N__13844),
            .lcout(\PCH_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIQUCA2_1_LC_1_8_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQUCA2_1_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQUCA2_1_LC_1_8_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \PCH_PWRGD.count_RNIQUCA2_1_LC_1_8_0  (
            .in0(N__13792),
            .in1(N__15016),
            .in2(_gnd_net_),
            .in3(N__13805),
            .lcout(\PCH_PWRGD.un2_count_1_axb_1 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIRP9H1_1_LC_1_8_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIRP9H1_1_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIRP9H1_1_LC_1_8_1 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \PCH_PWRGD.count_RNIRP9H1_1_LC_1_8_1  (
            .in0(_gnd_net_),
            .in1(N__14668),
            .in2(N__13832),
            .in3(N__14844),
            .lcout(\PCH_PWRGD.count_rst_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_1_8_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_1_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_1_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15379),
            .lcout(\PCH_PWRGD.N_2284_i ),
            .ltout(\PCH_PWRGD.N_2284_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIDKSB1_0_1_LC_1_8_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIDKSB1_0_1_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIDKSB1_0_1_LC_1_8_3 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNIDKSB1_0_1_LC_1_8_3  (
            .in0(_gnd_net_),
            .in1(N__13783),
            .in2(N__13829),
            .in3(N__29609),
            .lcout(\PCH_PWRGD.N_655 ),
            .ltout(\PCH_PWRGD.N_655_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIRP9H1_0_LC_1_8_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIRP9H1_0_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIRP9H1_0_LC_1_8_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNIRP9H1_0_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(N__15835),
            .in2(N__13826),
            .in3(N__25739),
            .lcout(\PCH_PWRGD.count_0_sqmuxa ),
            .ltout(\PCH_PWRGD.count_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_1_LC_1_8_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_1_LC_1_8_5 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_1_LC_1_8_5 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \PCH_PWRGD.count_1_LC_1_8_5  (
            .in0(_gnd_net_),
            .in1(N__14669),
            .in2(N__13823),
            .in3(N__13819),
            .lcout(\PCH_PWRGD.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32431),
            .ce(N__15071),
            .sr(N__14845));
    defparam \PCH_PWRGD.count_RNIQUCA2_0_1_LC_1_8_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQUCA2_0_1_LC_1_8_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQUCA2_0_1_LC_1_8_6 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \PCH_PWRGD.count_RNIQUCA2_0_1_LC_1_8_6  (
            .in0(N__15072),
            .in1(N__13804),
            .in2(N__13796),
            .in3(N__14509),
            .lcout(\PCH_PWRGD.count_1_i_a2_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIDKSB1_1_LC_1_8_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIDKSB1_1_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIDKSB1_1_LC_1_8_7 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \PCH_PWRGD.curr_state_RNIDKSB1_1_LC_1_8_7  (
            .in0(N__13784),
            .in1(N__13772),
            .in2(_gnd_net_),
            .in3(N__29610),
            .lcout(\PCH_PWRGD.N_670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIAKSS_2_LC_1_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNIAKSS_2_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIAKSS_2_LC_1_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNIAKSS_2_LC_1_9_0  (
            .in0(N__25734),
            .in1(N__13877),
            .in2(_gnd_net_),
            .in3(N__13891),
            .lcout(\POWERLED.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_2_LC_1_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_2_LC_1_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_2_LC_1_9_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_2_LC_1_9_1  (
            .in0(N__13892),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32436),
            .ce(N__16464),
            .sr(_gnd_net_));
    defparam \POWERLED.G_12_LC_1_9_2 .C_ON=1'b0;
    defparam \POWERLED.G_12_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_12_LC_1_9_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.G_12_LC_1_9_2  (
            .in0(N__25738),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22549),
            .lcout(G_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIALHT_11_LC_1_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_RNIALHT_11_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIALHT_11_LC_1_9_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIALHT_11_LC_1_9_3  (
            .in0(N__13865),
            .in1(N__25736),
            .in2(_gnd_net_),
            .in3(N__13936),
            .lcout(\POWERLED.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_11_LC_1_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_11_LC_1_9_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_11_LC_1_9_4 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_11_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13940),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32436),
            .ce(N__16464),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNICNTS_3_LC_1_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNICNTS_3_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNICNTS_3_LC_1_9_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNICNTS_3_LC_1_9_5  (
            .in0(N__13859),
            .in1(N__25735),
            .in2(_gnd_net_),
            .in3(N__13984),
            .lcout(\POWERLED.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_3_LC_1_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_3_LC_1_9_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_3_LC_1_9_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_3_LC_1_9_6  (
            .in0(N__13985),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32436),
            .ce(N__16464),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNICOIT_12_LC_1_9_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNICOIT_12_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNICOIT_12_LC_1_9_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNICOIT_12_LC_1_9_7  (
            .in0(N__14000),
            .in1(N__25737),
            .in2(_gnd_net_),
            .in3(N__14015),
            .lcout(\POWERLED.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIEQUS_4_LC_1_10_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNIEQUS_4_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIEQUS_4_LC_1_10_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNIEQUS_4_LC_1_10_0  (
            .in0(N__25747),
            .in1(N__13898),
            .in2(_gnd_net_),
            .in3(N__13969),
            .lcout(\POWERLED.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_0_LC_1_10_1 .C_ON=1'b0;
    defparam \POWERLED.count_0_LC_1_10_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_0_LC_1_10_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.count_0_LC_1_10_1  (
            .in0(N__14193),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17252),
            .lcout(\POWERLED.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32460),
            .ce(N__16463),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIE5D5_0_LC_1_10_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNIE5D5_0_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIE5D5_0_LC_1_10_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.count_RNIE5D5_0_LC_1_10_2  (
            .in0(N__17254),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14191),
            .lcout(),
            .ltout(\POWERLED.count_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNITFSJ_0_LC_1_10_3 .C_ON=1'b0;
    defparam \POWERLED.count_RNITFSJ_0_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNITFSJ_0_LC_1_10_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_RNITFSJ_0_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__13922),
            .in2(N__13916),
            .in3(N__25745),
            .lcout(\POWERLED.countZ0Z_0 ),
            .ltout(\POWERLED.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIE5D5_1_LC_1_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNIE5D5_1_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIE5D5_1_LC_1_10_4 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \POWERLED.count_RNIE5D5_1_LC_1_10_4  (
            .in0(N__17214),
            .in1(_gnd_net_),
            .in2(N__13913),
            .in3(N__14192),
            .lcout(),
            .ltout(\POWERLED.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIUGSJ_1_LC_1_10_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNIUGSJ_1_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIUGSJ_1_LC_1_10_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_RNIUGSJ_1_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__13904),
            .in2(N__13910),
            .in3(N__25746),
            .lcout(\POWERLED.countZ0Z_1 ),
            .ltout(\POWERLED.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_1_LC_1_10_6 .C_ON=1'b0;
    defparam \POWERLED.count_1_LC_1_10_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_1_LC_1_10_6 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \POWERLED.count_1_LC_1_10_6  (
            .in0(N__17253),
            .in1(_gnd_net_),
            .in2(N__13907),
            .in3(N__14194),
            .lcout(\POWERLED.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32460),
            .ce(N__16463),
            .sr(_gnd_net_));
    defparam \POWERLED.count_4_LC_1_10_7 .C_ON=1'b0;
    defparam \POWERLED.count_4_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_4_LC_1_10_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_4_LC_1_10_7  (
            .in0(N__13970),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32460),
            .ce(N__16463),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_LC_1_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__17251),
            .in2(N__17218),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\POWERLED.un1_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_RNIP7DE_LC_1_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_RNIP7DE_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_RNIP7DE_LC_1_11_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_RNIP7DE_LC_1_11_1  (
            .in0(N__14195),
            .in1(_gnd_net_),
            .in2(N__17179),
            .in3(N__13880),
            .lcout(\POWERLED.count_1_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_1 ),
            .carryout(\POWERLED.un1_count_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_2_c_RNIQ9EE_LC_1_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_2_c_RNIQ9EE_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_2_c_RNIQ9EE_LC_1_11_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_2_c_RNIQ9EE_LC_1_11_2  (
            .in0(N__14199),
            .in1(_gnd_net_),
            .in2(N__17140),
            .in3(N__13973),
            .lcout(\POWERLED.count_1_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_2_cZ0 ),
            .carryout(\POWERLED.un1_count_cry_3_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_3_c_RNIRBFE_LC_1_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_3_c_RNIRBFE_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_3_c_RNIRBFE_LC_1_11_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_3_c_RNIRBFE_LC_1_11_3  (
            .in0(N__14196),
            .in1(_gnd_net_),
            .in2(N__17098),
            .in3(N__13961),
            .lcout(\POWERLED.count_1_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_3_cZ0 ),
            .carryout(\POWERLED.un1_count_cry_4_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_4_c_RNISDGE_LC_1_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_4_c_RNISDGE_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_4_c_RNISDGE_LC_1_11_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_4_c_RNISDGE_LC_1_11_4  (
            .in0(N__14200),
            .in1(_gnd_net_),
            .in2(N__17058),
            .in3(N__13958),
            .lcout(\POWERLED.count_1_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_4_cZ0 ),
            .carryout(\POWERLED.un1_count_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_5_c_RNITFHE_LC_1_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_5_c_RNITFHE_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_5_c_RNITFHE_LC_1_11_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_5_c_RNITFHE_LC_1_11_5  (
            .in0(N__14197),
            .in1(_gnd_net_),
            .in2(N__17019),
            .in3(N__13955),
            .lcout(\POWERLED.count_1_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_5 ),
            .carryout(\POWERLED.un1_count_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_6_c_RNIUHIE_LC_1_11_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_6_c_RNIUHIE_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_6_c_RNIUHIE_LC_1_11_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_6_c_RNIUHIE_LC_1_11_6  (
            .in0(N__14201),
            .in1(N__16974),
            .in2(_gnd_net_),
            .in3(N__13952),
            .lcout(\POWERLED.count_1_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_6 ),
            .carryout(\POWERLED.un1_count_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_7_c_RNIVJJE_LC_1_11_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_7_c_RNIVJJE_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_7_c_RNIVJJE_LC_1_11_7 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_7_c_RNIVJJE_LC_1_11_7  (
            .in0(N__14198),
            .in1(_gnd_net_),
            .in2(N__17530),
            .in3(N__13949),
            .lcout(\POWERLED.count_1_8 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_7 ),
            .carryout(\POWERLED.un1_count_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_8_c_RNI0MKE_LC_1_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_8_c_RNI0MKE_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_8_c_RNI0MKE_LC_1_12_0 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_8_c_RNI0MKE_LC_1_12_0  (
            .in0(N__14184),
            .in1(_gnd_net_),
            .in2(N__17497),
            .in3(N__13946),
            .lcout(\POWERLED.count_1_9 ),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\POWERLED.un1_count_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_9_c_RNI1OLE_LC_1_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_9_c_RNI1OLE_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_9_c_RNI1OLE_LC_1_12_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_9_c_RNI1OLE_LC_1_12_1  (
            .in0(N__14187),
            .in1(_gnd_net_),
            .in2(N__17464),
            .in3(N__13943),
            .lcout(\POWERLED.count_1_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_9 ),
            .carryout(\POWERLED.un1_count_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_10_c_RNI9ITC_LC_1_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_10_c_RNI9ITC_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_10_c_RNI9ITC_LC_1_12_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_10_c_RNI9ITC_LC_1_12_2  (
            .in0(N__14185),
            .in1(_gnd_net_),
            .in2(N__17410),
            .in3(N__13925),
            .lcout(\POWERLED.count_1_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_10 ),
            .carryout(\POWERLED.un1_count_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_11_c_RNIAKUC_LC_1_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_11_c_RNIAKUC_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_11_c_RNIAKUC_LC_1_12_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_11_c_RNIAKUC_LC_1_12_3  (
            .in0(N__14188),
            .in1(_gnd_net_),
            .in2(N__17371),
            .in3(N__14027),
            .lcout(\POWERLED.count_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_11 ),
            .carryout(\POWERLED.un1_count_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_12_c_RNIBMVC_LC_1_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_12_c_RNIBMVC_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_12_c_RNIBMVC_LC_1_12_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_12_c_RNIBMVC_LC_1_12_4  (
            .in0(N__14186),
            .in1(_gnd_net_),
            .in2(N__17328),
            .in3(N__14024),
            .lcout(\POWERLED.count_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_12 ),
            .carryout(\POWERLED.un1_count_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_13_c_RNICO0D_LC_1_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_13_c_RNICO0D_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_13_c_RNICO0D_LC_1_12_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_13_c_RNICO0D_LC_1_12_5  (
            .in0(N__14189),
            .in1(_gnd_net_),
            .in2(N__17292),
            .in3(N__14021),
            .lcout(\POWERLED.count_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_13 ),
            .carryout(\POWERLED.un1_count_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_14_c_RNIDQ1D_LC_1_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_cry_14_c_RNIDQ1D_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_14_c_RNIDQ1D_LC_1_12_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un1_count_cry_14_c_RNIDQ1D_LC_1_12_6  (
            .in0(N__17640),
            .in1(N__14190),
            .in2(_gnd_net_),
            .in3(N__14018),
            .lcout(\POWERLED.un1_count_cry_14_c_RNIDQ1DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_12_LC_1_12_7 .C_ON=1'b0;
    defparam \POWERLED.count_12_LC_1_12_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_12_LC_1_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_12_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14014),
            .lcout(\POWERLED.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32469),
            .ce(N__16469),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNIE5D5_0_LC_1_13_2 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNIE5D5_0_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNIE5D5_0_LC_1_13_2 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \POWERLED.curr_state_RNIE5D5_0_LC_1_13_2  (
            .in0(N__16565),
            .in1(_gnd_net_),
            .in2(N__25744),
            .in3(N__15557),
            .lcout(\POWERLED.pwm_out_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_LC_1_13_3 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_LC_1_13_3 .SEQ_MODE=4'b1010;
    defparam \POWERLED.pwm_out_LC_1_13_3 .LUT_INIT=16'b1100111011000000;
    LogicCell40 \POWERLED.pwm_out_LC_1_13_3  (
            .in0(N__17608),
            .in1(N__14113),
            .in2(N__15530),
            .in3(N__16564),
            .lcout(\POWERLED.pwm_outZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32470),
            .ce(),
            .sr(N__15587));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNIAVUE_LC_1_13_4 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNIAVUE_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNIAVUE_LC_1_13_4 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_RNIAVUE_LC_1_13_4  (
            .in0(N__16566),
            .in1(N__16525),
            .in2(_gnd_net_),
            .in3(N__17607),
            .lcout(),
            .ltout(\POWERLED.N_437_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNICO541_0_LC_1_13_5 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNICO541_0_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNICO541_0_LC_1_13_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.curr_state_RNICO541_0_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__16511),
            .in2(N__13991),
            .in3(N__25697),
            .lcout(\POWERLED.N_2305_i ),
            .ltout(\POWERLED.N_2305_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNI_0_LC_1_13_6 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI_0_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI_0_LC_1_13_6 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \POWERLED.curr_state_RNI_0_LC_1_13_6  (
            .in0(N__15553),
            .in1(_gnd_net_),
            .in2(N__13988),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_660 ),
            .ltout(\POWERLED.N_660_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNIE5D5_0_0_LC_1_13_7 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNIE5D5_0_0_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNIE5D5_0_0_LC_1_13_7 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \POWERLED.curr_state_RNIE5D5_0_0_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14204),
            .in3(N__25698),
            .lcout(\POWERLED.count_0_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNIPOMA1_LC_1_14_1 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNIPOMA1_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNIPOMA1_LC_1_14_1 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_RNIPOMA1_LC_1_14_1  (
            .in0(N__17609),
            .in1(N__14123),
            .in2(N__16499),
            .in3(N__16568),
            .lcout(),
            .ltout(\POWERLED.pwm_out_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNIKIDQ1_LC_1_14_2 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNIKIDQ1_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNIKIDQ1_LC_1_14_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \POWERLED.pwm_out_RNIKIDQ1_LC_1_14_2  (
            .in0(N__16567),
            .in1(_gnd_net_),
            .in2(N__14117),
            .in3(N__14114),
            .lcout(pwrbtn_led),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_1_14_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_14_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_14_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_15_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_15_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \VPP_VDDQ.un1_vddq_en_LC_1_15_5  (
            .in0(N__33131),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14093),
            .lcout(vddq_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_0_LC_2_1_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_0_LC_2_1_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_0_LC_2_1_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_0_LC_2_1_0  (
            .in0(N__25426),
            .in1(N__14072),
            .in2(N__16142),
            .in3(N__16141),
            .lcout(\RSMRST_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_2_1_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .clk(N__32235),
            .ce(),
            .sr(N__20960));
    defparam \RSMRST_PWRGD.count_1_LC_2_1_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_1_LC_2_1_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_1_LC_2_1_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_1_LC_2_1_1  (
            .in0(N__25411),
            .in1(N__14060),
            .in2(_gnd_net_),
            .in3(N__14048),
            .lcout(\RSMRST_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .clk(N__32235),
            .ce(),
            .sr(N__20960));
    defparam \RSMRST_PWRGD.count_2_LC_2_1_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_2_LC_2_1_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_2_LC_2_1_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_2_LC_2_1_2  (
            .in0(N__25427),
            .in1(N__14044),
            .in2(_gnd_net_),
            .in3(N__14030),
            .lcout(\RSMRST_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .clk(N__32235),
            .ce(),
            .sr(N__20960));
    defparam \RSMRST_PWRGD.count_3_LC_2_1_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_3_LC_2_1_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_3_LC_2_1_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_3_LC_2_1_3  (
            .in0(N__25412),
            .in1(N__14348),
            .in2(_gnd_net_),
            .in3(N__14336),
            .lcout(\RSMRST_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .clk(N__32235),
            .ce(),
            .sr(N__20960));
    defparam \RSMRST_PWRGD.count_4_LC_2_1_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_4_LC_2_1_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_4_LC_2_1_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_4_LC_2_1_4  (
            .in0(N__25428),
            .in1(N__14333),
            .in2(_gnd_net_),
            .in3(N__14321),
            .lcout(\RSMRST_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .clk(N__32235),
            .ce(),
            .sr(N__20960));
    defparam \RSMRST_PWRGD.count_5_LC_2_1_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_5_LC_2_1_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_5_LC_2_1_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_5_LC_2_1_5  (
            .in0(N__25413),
            .in1(N__14314),
            .in2(_gnd_net_),
            .in3(N__14300),
            .lcout(\RSMRST_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .clk(N__32235),
            .ce(),
            .sr(N__20960));
    defparam \RSMRST_PWRGD.count_6_LC_2_1_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_6_LC_2_1_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_6_LC_2_1_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_6_LC_2_1_6  (
            .in0(N__25429),
            .in1(N__14297),
            .in2(_gnd_net_),
            .in3(N__14285),
            .lcout(\RSMRST_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .clk(N__32235),
            .ce(),
            .sr(N__20960));
    defparam \RSMRST_PWRGD.count_7_LC_2_1_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_7_LC_2_1_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_7_LC_2_1_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_7_LC_2_1_7  (
            .in0(N__25414),
            .in1(N__14282),
            .in2(_gnd_net_),
            .in3(N__14270),
            .lcout(\RSMRST_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .clk(N__32235),
            .ce(),
            .sr(N__20960));
    defparam \RSMRST_PWRGD.count_8_LC_2_2_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_8_LC_2_2_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_8_LC_2_2_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_8_LC_2_2_0  (
            .in0(N__25425),
            .in1(N__14267),
            .in2(_gnd_net_),
            .in3(N__14255),
            .lcout(\RSMRST_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_2_2_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .clk(N__32316),
            .ce(),
            .sr(N__20955));
    defparam \RSMRST_PWRGD.count_9_LC_2_2_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_9_LC_2_2_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_9_LC_2_2_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_9_LC_2_2_1  (
            .in0(N__25410),
            .in1(N__14252),
            .in2(_gnd_net_),
            .in3(N__14240),
            .lcout(\RSMRST_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .clk(N__32316),
            .ce(),
            .sr(N__20955));
    defparam \RSMRST_PWRGD.count_10_LC_2_2_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_10_LC_2_2_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_10_LC_2_2_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_10_LC_2_2_2  (
            .in0(N__25422),
            .in1(N__14236),
            .in2(_gnd_net_),
            .in3(N__14222),
            .lcout(\RSMRST_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .clk(N__32316),
            .ce(),
            .sr(N__20955));
    defparam \RSMRST_PWRGD.count_11_LC_2_2_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_11_LC_2_2_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_11_LC_2_2_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_11_LC_2_2_3  (
            .in0(N__25408),
            .in1(N__14219),
            .in2(_gnd_net_),
            .in3(N__14207),
            .lcout(\RSMRST_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .clk(N__32316),
            .ce(),
            .sr(N__20955));
    defparam \RSMRST_PWRGD.count_12_LC_2_2_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_12_LC_2_2_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_12_LC_2_2_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_12_LC_2_2_4  (
            .in0(N__25423),
            .in1(N__14444),
            .in2(_gnd_net_),
            .in3(N__14432),
            .lcout(\RSMRST_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .clk(N__32316),
            .ce(),
            .sr(N__20955));
    defparam \RSMRST_PWRGD.count_13_LC_2_2_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_13_LC_2_2_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_13_LC_2_2_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_13_LC_2_2_5  (
            .in0(N__25409),
            .in1(N__14429),
            .in2(_gnd_net_),
            .in3(N__14417),
            .lcout(\RSMRST_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .clk(N__32316),
            .ce(),
            .sr(N__20955));
    defparam \RSMRST_PWRGD.count_14_LC_2_2_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_14_LC_2_2_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_14_LC_2_2_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_14_LC_2_2_6  (
            .in0(N__25424),
            .in1(N__14414),
            .in2(_gnd_net_),
            .in3(N__14402),
            .lcout(\RSMRST_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .clk(N__32316),
            .ce(),
            .sr(N__20955));
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_2_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_2_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_2_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_2_7  (
            .in0(_gnd_net_),
            .in1(N__25193),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_15_LC_2_3_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_15_LC_2_3_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_esr_15_LC_2_3_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \RSMRST_PWRGD.count_esr_15_LC_2_3_0  (
            .in0(_gnd_net_),
            .in1(N__14392),
            .in2(_gnd_net_),
            .in3(N__14399),
            .lcout(\RSMRST_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32354),
            .ce(N__17732),
            .sr(N__20959));
    defparam \PCH_PWRGD.count_12_LC_2_4_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_12_LC_2_4_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_12_LC_2_4_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_12_LC_2_4_0  (
            .in0(N__14372),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32318),
            .ce(N__15139),
            .sr(N__14959));
    defparam \PCH_PWRGD.count_RNIGJUB4_12_LC_2_4_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIGJUB4_12_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIGJUB4_12_LC_2_4_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \PCH_PWRGD.count_RNIGJUB4_12_LC_2_4_1  (
            .in0(N__14378),
            .in1(N__15101),
            .in2(_gnd_net_),
            .in3(N__14371),
            .lcout(\PCH_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIMC9U1_LC_2_4_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIMC9U1_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIMC9U1_LC_2_4_2 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_c_RNIMC9U1_LC_2_4_2  (
            .in0(N__14359),
            .in1(N__15328),
            .in2(N__14750),
            .in3(N__14957),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIKFM84_5_LC_2_4_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIKFM84_5_LC_2_4_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIKFM84_5_LC_2_4_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.count_RNIKFM84_5_LC_2_4_3  (
            .in0(_gnd_net_),
            .in1(N__14561),
            .in2(N__14555),
            .in3(N__15099),
            .lcout(\PCH_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI58BH4_10_LC_2_4_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI58BH4_10_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI58BH4_10_LC_2_4_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \PCH_PWRGD.count_RNI58BH4_10_LC_2_4_4  (
            .in0(N__15100),
            .in1(N__15155),
            .in2(_gnd_net_),
            .in3(N__15178),
            .lcout(\PCH_PWRGD.un2_count_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIPCK99_0_1_LC_2_4_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIPCK99_0_1_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIPCK99_0_1_LC_2_4_5 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \PCH_PWRGD.count_RNIPCK99_0_1_LC_2_4_5  (
            .in0(N__14667),
            .in1(N__14686),
            .in2(_gnd_net_),
            .in3(N__15233),
            .lcout(\PCH_PWRGD.N_386 ),
            .ltout(\PCH_PWRGD.N_386_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNI3U0P1_LC_2_4_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNI3U0P1_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNI3U0P1_LC_2_4_6 .LUT_INIT=16'b0000000001100000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_c_RNI3U0P1_LC_2_4_6  (
            .in0(N__14540),
            .in1(N__14507),
            .in2(N__14522),
            .in3(N__14958),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIEGTB4_11_LC_2_4_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIEGTB4_11_LC_2_4_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIEGTB4_11_LC_2_4_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \PCH_PWRGD.count_RNIEGTB4_11_LC_2_4_7  (
            .in0(N__14519),
            .in1(_gnd_net_),
            .in2(N__14513),
            .in3(N__15102),
            .lcout(\PCH_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIOGBU1_LC_2_5_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIOGBU1_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIOGBU1_LC_2_5_0 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_c_RNIOGBU1_LC_2_5_0  (
            .in0(N__15329),
            .in1(N__14474),
            .in2(N__14462),
            .in3(N__14923),
            .lcout(\PCH_PWRGD.count_rst_7 ),
            .ltout(\PCH_PWRGD.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI05DA2_7_LC_2_5_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI05DA2_7_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI05DA2_7_LC_2_5_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.count_RNI05DA2_7_LC_2_5_1  (
            .in0(_gnd_net_),
            .in1(N__14758),
            .in2(N__14477),
            .in3(N__15088),
            .lcout(\PCH_PWRGD.un2_count_1_axb_7 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_7_LC_2_5_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_7_LC_2_5_2 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_7_LC_2_5_2 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \PCH_PWRGD.count_7_LC_2_5_2  (
            .in0(N__15330),
            .in1(N__14461),
            .in2(N__14447),
            .in3(N__14925),
            .lcout(\PCH_PWRGD.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32356),
            .ce(N__15136),
            .sr(N__14929));
    defparam \PCH_PWRGD.count_RNIK6UQA_1_LC_2_5_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIK6UQA_1_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIK6UQA_1_LC_2_5_3 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \PCH_PWRGD.count_RNIK6UQA_1_LC_2_5_3  (
            .in0(N__14687),
            .in1(N__14930),
            .in2(N__14675),
            .in3(N__15228),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNID4B5D_0_LC_2_5_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNID4B5D_0_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNID4B5D_0_LC_2_5_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNID4B5D_0_LC_2_5_4  (
            .in0(N__15137),
            .in1(_gnd_net_),
            .in2(N__14768),
            .in3(N__14627),
            .lcout(\PCH_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI05DA2_0_7_LC_2_5_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI05DA2_0_7_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI05DA2_0_7_LC_2_5_5 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \PCH_PWRGD.count_RNI05DA2_0_7_LC_2_5_5  (
            .in0(N__14765),
            .in1(N__14759),
            .in2(N__14749),
            .in3(N__15089),
            .lcout(),
            .ltout(\PCH_PWRGD.count_1_i_a2_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIPCK99_1_LC_2_5_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIPCK99_1_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIPCK99_1_LC_2_5_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNIPCK99_1_LC_2_5_6  (
            .in0(N__14717),
            .in1(N__14711),
            .in2(N__14702),
            .in3(N__14699),
            .lcout(\PCH_PWRGD.count_1_i_a2_12_0 ),
            .ltout(\PCH_PWRGD.count_1_i_a2_12_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_0_LC_2_5_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_0_LC_2_5_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_0_LC_2_5_7 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \PCH_PWRGD.count_0_LC_2_5_7  (
            .in0(N__14924),
            .in1(N__14670),
            .in2(N__14630),
            .in3(N__15229),
            .lcout(\PCH_PWRGD.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32356),
            .ce(N__15136),
            .sr(N__14929));
    defparam \PCH_PWRGD.count_RNIMS1C4_15_LC_2_6_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIMS1C4_15_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIMS1C4_15_LC_2_6_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PCH_PWRGD.count_RNIMS1C4_15_LC_2_6_0  (
            .in0(N__15215),
            .in1(N__15206),
            .in2(_gnd_net_),
            .in3(N__15055),
            .lcout(\PCH_PWRGD.countZ0Z_15 ),
            .ltout(\PCH_PWRGD.countZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIIMVB4_0_13_LC_2_6_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIIMVB4_0_13_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIIMVB4_0_13_LC_2_6_1 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \PCH_PWRGD.count_RNIIMVB4_0_13_LC_2_6_1  (
            .in0(N__15200),
            .in1(N__15188),
            .in2(N__14612),
            .in3(N__15131),
            .lcout(\PCH_PWRGD.count_1_i_a2_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIIMVB4_13_LC_2_6_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIIMVB4_13_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIIMVB4_13_LC_2_6_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \PCH_PWRGD.count_RNIIMVB4_13_LC_2_6_2  (
            .in0(N__15187),
            .in1(N__15053),
            .in2(_gnd_net_),
            .in3(N__15198),
            .lcout(\PCH_PWRGD.un2_count_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI58BH4_0_10_LC_2_6_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI58BH4_0_10_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI58BH4_0_10_LC_2_6_3 .LUT_INIT=16'b0000001000010011;
    LogicCell40 \PCH_PWRGD.count_RNI58BH4_0_10_LC_2_6_3  (
            .in0(N__15054),
            .in1(N__14596),
            .in2(N__15179),
            .in3(N__15151),
            .lcout(),
            .ltout(\PCH_PWRGD.count_1_i_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI55U5D_2_LC_2_6_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI55U5D_2_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI55U5D_2_LC_2_6_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PCH_PWRGD.count_RNI55U5D_2_LC_2_6_4  (
            .in0(N__14585),
            .in1(N__14570),
            .in2(N__14564),
            .in3(N__15239),
            .lcout(\PCH_PWRGD.count_1_i_a2_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_15_LC_2_6_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_15_LC_2_6_5 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_15_LC_2_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_15_LC_2_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15214),
            .lcout(\PCH_PWRGD.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32411),
            .ce(N__15130),
            .sr(N__14961));
    defparam \PCH_PWRGD.count_13_LC_2_6_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_13_LC_2_6_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_13_LC_2_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_13_LC_2_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15199),
            .lcout(\PCH_PWRGD.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32411),
            .ce(N__15130),
            .sr(N__14961));
    defparam \PCH_PWRGD.count_10_LC_2_6_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_10_LC_2_6_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_10_LC_2_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_10_LC_2_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15174),
            .lcout(\PCH_PWRGD.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32411),
            .ce(N__15130),
            .sr(N__14961));
    defparam \PCH_PWRGD.curr_state_1_LC_2_7_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_1_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_1_LC_2_7_0 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \PCH_PWRGD.curr_state_1_LC_2_7_0  (
            .in0(N__15840),
            .in1(N__15391),
            .in2(N__15352),
            .in3(N__15375),
            .lcout(\PCH_PWRGD.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32402),
            .ce(N__16462),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_2_7_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_2_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_0_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15406),
            .lcout(\PCH_PWRGD.N_2266_i ),
            .ltout(\PCH_PWRGD.N_2266_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_0_LC_2_7_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_0_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_0_LC_2_7_2 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m4_0_0_LC_2_7_2  (
            .in0(N__15335),
            .in1(N__15798),
            .in2(N__14780),
            .in3(N__15373),
            .lcout(\PCH_PWRGD.curr_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_i_a2_LC_2_7_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_i_a2_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_i_a2_LC_2_7_3 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m6_i_i_a2_LC_2_7_3  (
            .in0(N__15392),
            .in1(N__15334),
            .in2(N__15380),
            .in3(N__15841),
            .lcout(),
            .ltout(\PCH_PWRGD.m6_i_i_a2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIC58V1_1_LC_2_7_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIC58V1_1_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIC58V1_1_LC_2_7_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.curr_state_RNIC58V1_1_LC_2_7_4  (
            .in0(_gnd_net_),
            .in1(N__14777),
            .in2(N__14771),
            .in3(N__25732),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIB48V1_0_LC_2_7_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIB48V1_0_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIB48V1_0_LC_2_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \PCH_PWRGD.curr_state_RNIB48V1_0_LC_2_7_5  (
            .in0(N__25733),
            .in1(N__15266),
            .in2(_gnd_net_),
            .in3(N__15413),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_0 ),
            .ltout(\PCH_PWRGD.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_0_a2_0_LC_2_7_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_0_a2_0_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_0_a2_0_LC_2_7_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m4_0_0_a2_0_LC_2_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15395),
            .in3(N__15390),
            .lcout(\PCH_PWRGD.curr_state_0_sqmuxa ),
            .ltout(\PCH_PWRGD.curr_state_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_0_LC_2_7_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_0_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_0_LC_2_7_7 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \PCH_PWRGD.curr_state_0_LC_2_7_7  (
            .in0(N__15374),
            .in1(N__15336),
            .in2(N__15269),
            .in3(N__15839),
            .lcout(\PCH_PWRGD.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32402),
            .ce(N__16462),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_0_LC_2_8_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_0_LC_2_8_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_0_LC_2_8_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_0_LC_2_8_0  (
            .in0(N__16369),
            .in1(N__16329),
            .in2(N__22334),
            .in3(N__16046),
            .lcout(\VPP_VDDQ.curr_state_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32430),
            .ce(N__16465),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_2_8_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_2_8_1 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_2_8_1  (
            .in0(N__16401),
            .in1(N__16108),
            .in2(N__16083),
            .in3(N__16367),
            .lcout(),
            .ltout(\VPP_VDDQ.N_53_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIMPBA_1_LC_2_8_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIMPBA_1_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIMPBA_1_LC_2_8_2 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIMPBA_1_LC_2_8_2  (
            .in0(N__25741),
            .in1(_gnd_net_),
            .in2(N__15260),
            .in3(N__15254),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_1 ),
            .ltout(\VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_1_LC_2_8_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_1_LC_2_8_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_1_LC_2_8_3 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \VPP_VDDQ.curr_state_2_1_LC_2_8_3  (
            .in0(N__16400),
            .in1(N__16109),
            .in2(N__15257),
            .in3(N__16370),
            .lcout(\VPP_VDDQ.curr_state_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32430),
            .ce(N__16465),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_LC_2_8_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_LC_2_8_4 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_LC_2_8_4  (
            .in0(N__22330),
            .in1(N__16330),
            .in2(N__16380),
            .in3(N__16045),
            .lcout(),
            .ltout(\VPP_VDDQ.m4_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_2_8_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_2_8_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(N__15248),
            .in2(N__15242),
            .in3(N__25740),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIE5D5_0_LC_2_8_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIE5D5_0_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIE5D5_0_LC_2_8_6 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIE5D5_0_LC_2_8_6  (
            .in0(N__25742),
            .in1(_gnd_net_),
            .in2(N__15518),
            .in3(N__16402),
            .lcout(\VPP_VDDQ.N_60 ),
            .ltout(\VPP_VDDQ.N_60_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNINI731_0_LC_2_8_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNINI731_0_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNINI731_0_LC_2_8_7 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNINI731_0_LC_2_8_7  (
            .in0(N__16493),
            .in1(N__16368),
            .in2(N__15515),
            .in3(N__22331),
            .lcout(\VPP_VDDQ.delayed_vddq_ok_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_2_9_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_2_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNO_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15498),
            .lcout(\VPP_VDDQ.N_60_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_2_9_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_2_9_1 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_2_9_1 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_LC_2_9_1  (
            .in0(N__15472),
            .in1(N__22323),
            .in2(N__15485),
            .in3(N__15499),
            .lcout(\VPP_VDDQ.delayed_vddq_okZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32435),
            .ce(),
            .sr(N__15512));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNIUP8M1_LC_2_9_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNIUP8M1_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNIUP8M1_LC_2_9_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNIUP8M1_LC_2_9_2  (
            .in0(N__15500),
            .in1(N__15484),
            .in2(N__22333),
            .in3(N__15473),
            .lcout(),
            .ltout(VPP_VDDQ_delayed_vddq_ok_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_PWRGD_LC_2_9_3 .C_ON=1'b0;
    defparam \POWERLED.VCCST_PWRGD_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_PWRGD_LC_2_9_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \POWERLED.VCCST_PWRGD_LC_2_9_3  (
            .in0(N__15983),
            .in1(_gnd_net_),
            .in2(N__15464),
            .in3(_gnd_net_),
            .lcout(vccst_pwrgd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_2_9_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_2_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_1_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16073),
            .lcout(\VPP_VDDQ.curr_state_2_RNIZ0Z_1 ),
            .ltout(\VPP_VDDQ.curr_state_2_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_a2_0_LC_2_9_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_a2_0_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_a2_0_LC_2_9_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_a2_0_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15443),
            .in3(N__22322),
            .lcout(N_639),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_0_LC_2_9_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_0_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_0_LC_2_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_0_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15982),
            .lcout(pch_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI1Q9V_10_LC_2_9_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNI1Q9V_10_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI1Q9V_10_LC_2_9_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI1Q9V_10_LC_2_9_7  (
            .in0(N__15692),
            .in1(N__25743),
            .in2(_gnd_net_),
            .in3(N__15707),
            .lcout(\POWERLED.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_0_LC_2_10_0 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_0_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_0_LC_2_10_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.pwm_out_RNO_0_LC_2_10_0  (
            .in0(N__25756),
            .in1(N__16570),
            .in2(_gnd_net_),
            .in3(N__15552),
            .lcout(\POWERLED.pwm_out_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_2_LC_2_10_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_2_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_2_LC_2_10_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.count_RNI_2_LC_2_10_1  (
            .in0(N__17169),
            .in1(N__17094),
            .in2(_gnd_net_),
            .in3(N__17130),
            .lcout(\POWERLED.un79_clk_100khzlt6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_7_LC_2_10_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_7_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_7_LC_2_10_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.count_RNI_7_LC_2_10_2  (
            .in0(N__17493),
            .in1(N__17526),
            .in2(_gnd_net_),
            .in3(N__16975),
            .lcout(\POWERLED.un79_clk_100khzlto15_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_15_LC_2_10_3 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_15_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_15_LC_2_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_RNI_15_LC_2_10_3  (
            .in0(N__17364),
            .in1(N__17329),
            .in2(N__17644),
            .in3(N__17293),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlto15_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_5_LC_2_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_5_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_5_LC_2_10_4 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \POWERLED.count_RNI_5_LC_2_10_4  (
            .in0(N__15575),
            .in1(N__17020),
            .in2(N__15569),
            .in3(N__17059),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlto15_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_10_LC_2_10_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_10_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_10_LC_2_10_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \POWERLED.count_RNI_10_LC_2_10_5  (
            .in0(N__15566),
            .in1(N__17454),
            .in2(N__15560),
            .in3(N__17403),
            .lcout(\POWERLED.un79_clk_100khz ),
            .ltout(\POWERLED.un79_clk_100khz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_1_LC_2_10_6 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_1_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_1_LC_2_10_6 .LUT_INIT=16'b0011001101111111;
    LogicCell40 \POWERLED.pwm_out_RNO_1_LC_2_10_6  (
            .in0(N__25757),
            .in1(N__16494),
            .in2(N__15533),
            .in3(N__16569),
            .lcout(\POWERLED.g0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNII1MT_15_LC_2_11_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNII1MT_15_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNII1MT_15_LC_2_11_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNII1MT_15_LC_2_11_0  (
            .in0(N__15656),
            .in1(N__25755),
            .in2(_gnd_net_),
            .in3(N__15664),
            .lcout(\POWERLED.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_15_LC_2_11_1 .C_ON=1'b0;
    defparam \POWERLED.count_15_LC_2_11_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_15_LC_2_11_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_15_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15668),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32459),
            .ce(N__16466),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIK32T_7_LC_2_11_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNIK32T_7_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIK32T_7_LC_2_11_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIK32T_7_LC_2_11_2  (
            .in0(N__15641),
            .in1(N__25752),
            .in2(_gnd_net_),
            .in3(N__15649),
            .lcout(\POWERLED.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_7_LC_2_11_3 .C_ON=1'b0;
    defparam \POWERLED.count_7_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_7_LC_2_11_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_7_LC_2_11_3  (
            .in0(N__15650),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32459),
            .ce(N__16466),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIM63T_8_LC_2_11_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNIM63T_8_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIM63T_8_LC_2_11_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIM63T_8_LC_2_11_4  (
            .in0(N__15626),
            .in1(N__25753),
            .in2(_gnd_net_),
            .in3(N__15634),
            .lcout(\POWERLED.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_8_LC_2_11_5 .C_ON=1'b0;
    defparam \POWERLED.count_8_LC_2_11_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_8_LC_2_11_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_8_LC_2_11_5  (
            .in0(N__15635),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32459),
            .ce(N__16466),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIO94T_9_LC_2_11_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNIO94T_9_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIO94T_9_LC_2_11_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIO94T_9_LC_2_11_6  (
            .in0(N__15611),
            .in1(N__25754),
            .in2(_gnd_net_),
            .in3(N__15619),
            .lcout(\POWERLED.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_9_LC_2_11_7 .C_ON=1'b0;
    defparam \POWERLED.count_9_LC_2_11_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_9_LC_2_11_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_9_LC_2_11_7  (
            .in0(N__15620),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32459),
            .ce(N__16466),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIERJT_13_LC_2_12_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNIERJT_13_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIERJT_13_LC_2_12_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIERJT_13_LC_2_12_0  (
            .in0(N__15593),
            .in1(N__25750),
            .in2(_gnd_net_),
            .in3(N__15601),
            .lcout(\POWERLED.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_13_LC_2_12_1 .C_ON=1'b0;
    defparam \POWERLED.count_13_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_13_LC_2_12_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_13_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15605),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32468),
            .ce(N__16468),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIGTVS_5_LC_2_12_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNIGTVS_5_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIGTVS_5_LC_2_12_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIGTVS_5_LC_2_12_2  (
            .in0(N__15746),
            .in1(N__25748),
            .in2(_gnd_net_),
            .in3(N__15754),
            .lcout(\POWERLED.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_5_LC_2_12_3 .C_ON=1'b0;
    defparam \POWERLED.count_5_LC_2_12_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_5_LC_2_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_5_LC_2_12_3  (
            .in0(N__15755),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32468),
            .ce(N__16468),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIGUKT_14_LC_2_12_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNIGUKT_14_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIGUKT_14_LC_2_12_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIGUKT_14_LC_2_12_4  (
            .in0(N__15728),
            .in1(N__25751),
            .in2(_gnd_net_),
            .in3(N__15736),
            .lcout(\POWERLED.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_14_LC_2_12_5 .C_ON=1'b0;
    defparam \POWERLED.count_14_LC_2_12_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_14_LC_2_12_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_14_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15740),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32468),
            .ce(N__16468),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNII01T_6_LC_2_12_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNII01T_6_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNII01T_6_LC_2_12_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNII01T_6_LC_2_12_6  (
            .in0(N__15713),
            .in1(N__25749),
            .in2(_gnd_net_),
            .in3(N__15721),
            .lcout(\POWERLED.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_6_LC_2_12_7 .C_ON=1'b0;
    defparam \POWERLED.count_6_LC_2_12_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_6_LC_2_12_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_6_LC_2_12_7  (
            .in0(N__15722),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32468),
            .ce(N__16468),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_2_13_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_2_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18512),
            .lcout(\POWERLED.mult1_un96_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_10_LC_2_13_2 .C_ON=1'b0;
    defparam \POWERLED.count_10_LC_2_13_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_10_LC_2_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_10_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15706),
            .lcout(\POWERLED.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32467),
            .ce(N__16467),
            .sr(_gnd_net_));
    defparam SLP_SUSn_RNIN4K9_LC_2_14_2.C_ON=1'b0;
    defparam SLP_SUSn_RNIN4K9_LC_2_14_2.SEQ_MODE=4'b0000;
    defparam SLP_SUSn_RNIN4K9_LC_2_14_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 SLP_SUSn_RNIN4K9_LC_2_14_2 (
            .in0(N__16267),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(v33a_enn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_6_LC_4_2_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_6_LC_4_2_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_6_LC_4_2_2 .LUT_INIT=16'b0000011001100110;
    LogicCell40 \HDA_STRAP.count_6_LC_4_2_2  (
            .in0(N__17696),
            .in1(N__18874),
            .in2(N__19162),
            .in3(N__19211),
            .lcout(\HDA_STRAP.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32166),
            .ce(N__25310),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_8_LC_4_2_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_8_LC_4_2_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_8_LC_4_2_3 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \HDA_STRAP.count_8_LC_4_2_3  (
            .in0(N__19209),
            .in1(N__18909),
            .in2(N__19145),
            .in3(N__17684),
            .lcout(\HDA_STRAP.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32166),
            .ce(N__25310),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_10_LC_4_2_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_10_LC_4_2_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_10_LC_4_2_4 .LUT_INIT=16'b0000011001100110;
    LogicCell40 \HDA_STRAP.count_10_LC_4_2_4  (
            .in0(N__17672),
            .in1(N__18766),
            .in2(N__19161),
            .in3(N__19210),
            .lcout(\HDA_STRAP.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32166),
            .ce(N__25310),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_11_LC_4_2_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_11_LC_4_2_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_11_LC_4_2_5 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \HDA_STRAP.count_11_LC_4_2_5  (
            .in0(N__19208),
            .in1(N__18783),
            .in2(N__19144),
            .in3(N__17663),
            .lcout(\HDA_STRAP.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32166),
            .ce(N__25310),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_4_2_6 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_4_2_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \HDA_STRAP.curr_state_RNO_0_2_LC_4_2_6  (
            .in0(_gnd_net_),
            .in1(N__19120),
            .in2(_gnd_net_),
            .in3(N__19207),
            .lcout(),
            .ltout(\HDA_STRAP.N_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_2_LC_4_2_7 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_2_LC_4_2_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_2_LC_4_2_7 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \HDA_STRAP.curr_state_2_LC_4_2_7  (
            .in0(N__15893),
            .in1(N__15905),
            .in2(N__15764),
            .in3(N__15970),
            .lcout(\HDA_STRAP.curr_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32166),
            .ce(N__25310),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIT2822_LC_4_3_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIT2822_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIT2822_LC_4_3_0 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNIT2822_LC_4_3_0  (
            .in0(N__15805),
            .in1(N__15778),
            .in2(N__15815),
            .in3(N__16492),
            .lcout(),
            .ltout(\PCH_PWRGD.delayed_vccin_okZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_LC_4_3_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_LC_4_3_1 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_LC_4_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15761),
            .in3(N__29617),
            .lcout(N_428),
            .ltout(N_428_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_1_LC_4_3_2 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_1_LC_4_3_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_1_LC_4_3_2 .LUT_INIT=16'b0110111000101010;
    LogicCell40 \HDA_STRAP.curr_state_1_LC_4_3_2  (
            .in0(N__15953),
            .in1(N__15934),
            .in2(N__15758),
            .in3(N__19214),
            .lcout(\HDA_STRAP.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32126),
            .ce(N__25308),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIH91A_0_LC_4_3_3 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIH91A_0_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIH91A_0_LC_4_3_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \HDA_STRAP.curr_state_RNIH91A_0_LC_4_3_3  (
            .in0(_gnd_net_),
            .in1(N__15949),
            .in2(_gnd_net_),
            .in3(N__15920),
            .lcout(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_4_3_4 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_4_3_4 .LUT_INIT=16'b0000001001010010;
    LogicCell40 \HDA_STRAP.curr_state_RNO_0_0_LC_4_3_4  (
            .in0(N__15951),
            .in1(N__16001),
            .in2(N__15933),
            .in3(N__19213),
            .lcout(),
            .ltout(\HDA_STRAP.m14_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_0_LC_4_3_5 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_0_LC_4_3_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_0_LC_4_3_5 .LUT_INIT=16'b1111000011111001;
    LogicCell40 \HDA_STRAP.curr_state_0_LC_4_3_5  (
            .in0(N__15935),
            .in1(N__15952),
            .in2(N__15986),
            .in3(N__15969),
            .lcout(\HDA_STRAP.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32126),
            .ce(N__25308),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIRV1F_2_LC_4_3_6 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIRV1F_2_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIRV1F_2_LC_4_3_6 .LUT_INIT=16'b0000000001011111;
    LogicCell40 \HDA_STRAP.curr_state_RNIRV1F_2_LC_4_3_6  (
            .in0(N__15950),
            .in1(_gnd_net_),
            .in2(N__15932),
            .in3(N__15904),
            .lcout(\HDA_STRAP.HDA_SDO_ATP_3_0 ),
            .ltout(\HDA_STRAP.HDA_SDO_ATP_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_4_3_7 .C_ON=1'b0;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_4_3_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_4_3_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \HDA_STRAP.HDA_SDO_ATP_LC_4_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15887),
            .in3(_gnd_net_),
            .lcout(hda_sdo_atp),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32126),
            .ce(N__25308),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_1_0_LC_4_4_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_1_0_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_1_0_LC_4_4_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_1_0_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(N__15869),
            .in2(_gnd_net_),
            .in3(N__15845),
            .lcout(\PCH_PWRGD.N_38_f0 ),
            .ltout(\PCH_PWRGD.N_38_f0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_4_4_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_4_4_1 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_4_4_1 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_LC_4_4_1  (
            .in0(N__15779),
            .in1(N__15806),
            .in2(N__15782),
            .in3(N__16495),
            .lcout(\PCH_PWRGD.delayed_vccin_ok_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32201),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_4_4_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_4_4_3 .LUT_INIT=16'b0000111010011001;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_4_4_3  (
            .in0(N__23311),
            .in1(N__33144),
            .in2(N__23267),
            .in3(N__25403),
            .lcout(),
            .ltout(\VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_4_4_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_4_4_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_4_4_4 .LUT_INIT=16'b1110001111000010;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_LC_4_4_4  (
            .in0(N__33145),
            .in1(N__23312),
            .in2(N__15767),
            .in3(N__23345),
            .lcout(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32201),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_4_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_4_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21509),
            .lcout(\POWERLED.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_4_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_4_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_4_6  (
            .in0(N__16688),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_4_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_4_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21668),
            .lcout(\POWERLED.mult1_un54_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIM9AN_1_LC_4_5_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIM9AN_1_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIM9AN_1_LC_4_5_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_2_RNIM9AN_1_LC_4_5_0  (
            .in0(N__19764),
            .in1(N__16009),
            .in2(_gnd_net_),
            .in3(N__16016),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_4_5_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_4_5_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_0_1_LC_4_5_1  (
            .in0(N__16102),
            .in1(N__16087),
            .in2(_gnd_net_),
            .in3(N__16385),
            .lcout(\VPP_VDDQ.count_2_1_sqmuxa ),
            .ltout(\VPP_VDDQ.count_2_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_0_LC_4_5_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_0_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_0_LC_4_5_2 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \VPP_VDDQ.count_2_RNI_0_LC_4_5_2  (
            .in0(N__17821),
            .in1(_gnd_net_),
            .in2(N__16031),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIL8AN_0_LC_4_5_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIL8AN_0_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIL8AN_0_LC_4_5_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIL8AN_0_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(N__16022),
            .in2(N__16028),
            .in3(N__19763),
            .lcout(\VPP_VDDQ.count_2Z0Z_0 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_0_LC_4_5_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_0_LC_4_5_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_0_LC_4_5_4 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \VPP_VDDQ.count_2_0_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16025),
            .in3(N__18149),
            .lcout(\VPP_VDDQ.count_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32282),
            .ce(N__19765),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_1_LC_4_5_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_1_LC_4_5_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_1_LC_4_5_5 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \VPP_VDDQ.count_2_1_LC_4_5_5  (
            .in0(N__17816),
            .in1(_gnd_net_),
            .in2(N__18160),
            .in3(N__17787),
            .lcout(\VPP_VDDQ.count_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32282),
            .ce(N__19765),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_1_LC_4_5_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_4_5_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \VPP_VDDQ.count_2_RNI_1_LC_4_5_6  (
            .in0(N__17788),
            .in1(N__18145),
            .in2(_gnd_net_),
            .in3(N__17815),
            .lcout(\VPP_VDDQ.count_2_1_1 ),
            .ltout(\VPP_VDDQ.count_2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIM9AN_0_1_LC_4_5_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIM9AN_0_1_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIM9AN_0_1_LC_4_5_7 .LUT_INIT=16'b0000001100010001;
    LogicCell40 \VPP_VDDQ.count_2_RNIM9AN_0_1_LC_4_5_7  (
            .in0(N__16010),
            .in1(N__17820),
            .in2(N__16274),
            .in3(N__19766),
            .lcout(\VPP_VDDQ.un9_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_4_6_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_4_6_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_4_6_1  (
            .in0(N__16271),
            .in1(N__16238),
            .in2(N__16221),
            .in3(N__16177),
            .lcout(rsmrst_pwrgd_signal),
            .ltout(rsmrst_pwrgd_signal_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_4_6_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_4_6_2 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(N__21197),
            .in2(N__16148),
            .in3(N__21168),
            .lcout(),
            .ltout(\RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_0_LC_4_6_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_0_LC_4_6_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_0_LC_4_6_3 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \RSMRST_PWRGD.curr_state_0_LC_4_6_3  (
            .in0(N__21198),
            .in1(_gnd_net_),
            .in2(N__16145),
            .in3(N__20918),
            .lcout(RSMRST_PWRGD_curr_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32299),
            .ce(N__25314),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_4_6_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_4_6_4 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_4_6_4  (
            .in0(N__26804),
            .in1(N__21196),
            .in2(_gnd_net_),
            .in3(N__21167),
            .lcout(\RSMRST_PWRGD.N_264_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIFQNU_1_7_LC_4_6_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIFQNU_1_7_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIFQNU_1_7_LC_4_6_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIFQNU_1_7_LC_4_6_5  (
            .in0(N__17990),
            .in1(N__16304),
            .in2(N__17956),
            .in3(N__16283),
            .lcout(),
            .ltout(\VPP_VDDQ.un9_clk_100khz_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI0JCD2_1_LC_4_6_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI0JCD2_1_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI0JCD2_1_LC_4_6_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNI0JCD2_1_LC_4_6_6  (
            .in0(N__19829),
            .in1(N__16118),
            .in2(N__16112),
            .in3(N__19619),
            .lcout(\VPP_VDDQ.N_1_i ),
            .ltout(\VPP_VDDQ.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_a2_1_LC_4_6_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_a2_1_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_a2_1_LC_4_6_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_a2_1_LC_4_6_7  (
            .in0(N__16088),
            .in1(_gnd_net_),
            .in2(N__16049),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.N_664 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_9_LC_4_7_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_9_LC_4_7_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_9_LC_4_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_9_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18004),
            .lcout(\VPP_VDDQ.count_2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32284),
            .ce(N__19776),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI1KAM_0_LC_4_7_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI1KAM_0_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI1KAM_0_LC_4_7_1 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI1KAM_0_LC_4_7_1  (
            .in0(N__16409),
            .in1(N__16384),
            .in2(N__16340),
            .in3(N__16491),
            .lcout(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_2_RNI1KAMZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIFQNU_7_LC_4_7_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIFQNU_7_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIFQNU_7_LC_4_7_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIFQNU_7_LC_4_7_2  (
            .in0(_gnd_net_),
            .in1(N__18050),
            .in2(N__16316),
            .in3(N__16297),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIJ0QU_9_LC_4_7_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIJ0QU_9_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIJ0QU_9_LC_4_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIJ0QU_9_LC_4_7_3  (
            .in0(N__18005),
            .in1(N__16313),
            .in2(_gnd_net_),
            .in3(N__19779),
            .lcout(\VPP_VDDQ.count_2Z0Z_9 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIFQNU_0_7_LC_4_7_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIFQNU_0_7_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIFQNU_0_7_LC_4_7_4 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \VPP_VDDQ.count_2_RNIFQNU_0_7_LC_4_7_4  (
            .in0(N__19778),
            .in1(N__18049),
            .in2(N__16307),
            .in3(N__16298),
            .lcout(\VPP_VDDQ.un9_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_7_LC_4_7_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_7_LC_4_7_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_7_LC_4_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_7_LC_4_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18043),
            .lcout(\VPP_VDDQ.count_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32284),
            .ce(N__19776),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI52L41_11_LC_4_7_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI52L41_11_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI52L41_11_LC_4_7_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_2_RNI52L41_11_LC_4_7_6  (
            .in0(N__19777),
            .in1(N__16289),
            .in2(_gnd_net_),
            .in3(N__17939),
            .lcout(\VPP_VDDQ.count_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_11_LC_4_7_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_11_LC_4_7_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_11_LC_4_7_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_2_11_LC_4_7_7  (
            .in0(N__17938),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32284),
            .ce(N__19776),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_15_LC_4_8_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_15_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_15_LC_4_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_2_RNI_15_LC_4_8_0  (
            .in0(N__17872),
            .in1(N__17923),
            .in2(N__17900),
            .in3(N__18217),
            .lcout(\VPP_VDDQ.un9_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI75M41_12_LC_4_8_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI75M41_12_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI75M41_12_LC_4_8_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNI75M41_12_LC_4_8_1  (
            .in0(N__17912),
            .in1(N__16592),
            .in2(_gnd_net_),
            .in3(N__19800),
            .lcout(\VPP_VDDQ.count_2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_12_LC_4_8_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_12_LC_4_8_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_12_LC_4_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_12_LC_4_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17911),
            .lcout(\VPP_VDDQ.count_2_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32397),
            .ce(N__19799),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI98N41_13_LC_4_8_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI98N41_13_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI98N41_13_LC_4_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNI98N41_13_LC_4_8_3  (
            .in0(N__17885),
            .in1(N__16586),
            .in2(_gnd_net_),
            .in3(N__19801),
            .lcout(\VPP_VDDQ.count_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_13_LC_4_8_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_13_LC_4_8_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_13_LC_4_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_13_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17884),
            .lcout(\VPP_VDDQ.count_2_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32397),
            .ce(N__19799),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIBBO41_14_LC_4_8_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIBBO41_14_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIBBO41_14_LC_4_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIBBO41_14_LC_4_8_5  (
            .in0(N__17861),
            .in1(N__16580),
            .in2(_gnd_net_),
            .in3(N__19802),
            .lcout(\VPP_VDDQ.count_2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_14_LC_4_8_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_14_LC_4_8_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_14_LC_4_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_14_LC_4_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17860),
            .lcout(\VPP_VDDQ.count_2_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32397),
            .ce(N__19799),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIDEP41_15_LC_4_8_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIDEP41_15_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIDEP41_15_LC_4_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_2_RNIDEP41_15_LC_4_8_7  (
            .in0(N__19753),
            .in1(N__18110),
            .in2(_gnd_net_),
            .in3(N__18121),
            .lcout(\VPP_VDDQ.count_2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_0_LC_4_9_0 .C_ON=1'b0;
    defparam \POWERLED.curr_state_0_LC_4_9_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.curr_state_0_LC_4_9_0 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \POWERLED.curr_state_0_LC_4_9_0  (
            .in0(N__17603),
            .in1(N__16574),
            .in2(_gnd_net_),
            .in3(N__16532),
            .lcout(\POWERLED.curr_state_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32406),
            .ce(N__16461),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI7EJU_3_LC_4_9_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI7EJU_3_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI7EJU_3_LC_4_9_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_2_RNI7EJU_3_LC_4_9_1  (
            .in0(N__19772),
            .in1(N__17720),
            .in2(_gnd_net_),
            .in3(N__17767),
            .lcout(\VPP_VDDQ.count_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIBKLU_5_LC_4_9_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIBKLU_5_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIBKLU_5_LC_4_9_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.count_2_RNIBKLU_5_LC_4_9_2  (
            .in0(N__17849),
            .in1(N__19773),
            .in2(_gnd_net_),
            .in3(N__17749),
            .lcout(\VPP_VDDQ.count_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIHTOU_8_LC_4_9_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIHTOU_8_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIHTOU_8_LC_4_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_2_RNIHTOU_8_LC_4_9_3  (
            .in0(N__19774),
            .in1(N__17840),
            .in2(_gnd_net_),
            .in3(N__18029),
            .lcout(\VPP_VDDQ.count_2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIS3FU_10_LC_4_9_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIS3FU_10_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIS3FU_10_LC_4_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNIS3FU_10_LC_4_9_4  (
            .in0(N__17831),
            .in1(N__17974),
            .in2(_gnd_net_),
            .in3(N__19775),
            .lcout(\VPP_VDDQ.count_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_4_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_4_9_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(N__16684),
            .in2(_gnd_net_),
            .in3(N__16754),
            .lcout(\POWERLED.mult1_un124_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_9_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_9_7  (
            .in0(N__16683),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un117_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_10_0  (
            .in0(_gnd_net_),
            .in1(N__21530),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_10_0_),
            .carryout(\POWERLED.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(N__16643),
            .in2(N__16631),
            .in3(N__16619),
            .lcout(\POWERLED.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(N__16750),
            .in2(N__16616),
            .in3(N__16604),
            .lcout(\POWERLED.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(N__16670),
            .in2(N__16736),
            .in3(N__16601),
            .lcout(\POWERLED.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(N__16724),
            .in2(N__16682),
            .in3(N__16598),
            .lcout(\POWERLED.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_10_5  (
            .in0(N__18371),
            .in1(N__16760),
            .in2(N__16715),
            .in3(N__16595),
            .lcout(\POWERLED.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_10_6  (
            .in0(N__16700),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16763),
            .lcout(\POWERLED.mult1_un124_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_4_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_4_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_4_10_7  (
            .in0(N__16711),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16669),
            .lcout(\POWERLED.mult1_un124_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_11_0  (
            .in0(_gnd_net_),
            .in1(N__21502),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_11_0_),
            .carryout(\POWERLED.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(N__20378),
            .in2(N__16858),
            .in3(N__16739),
            .lcout(\POWERLED.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(N__16854),
            .in2(N__16841),
            .in3(N__16727),
            .lcout(\POWERLED.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(N__16829),
            .in2(N__16790),
            .in3(N__16718),
            .lcout(\POWERLED.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(N__16820),
            .in2(N__16789),
            .in3(N__16703),
            .lcout(\POWERLED.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_11_5  (
            .in0(N__16668),
            .in1(N__16811),
            .in2(N__16859),
            .in3(N__16694),
            .lcout(\POWERLED.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_11_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_11_6  (
            .in0(N__16802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16691),
            .lcout(\POWERLED.mult1_un117_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16782),
            .lcout(\POWERLED.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_4_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_4_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(N__21482),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(\POWERLED.mult1_un110_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_4_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_4_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__20399),
            .in2(N__16876),
            .in3(N__16832),
            .lcout(\POWERLED.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_4_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_4_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(N__16872),
            .in2(N__16937),
            .in3(N__16823),
            .lcout(\POWERLED.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_4_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_4_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(N__16925),
            .in2(N__18410),
            .in3(N__16814),
            .lcout(\POWERLED.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_4_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_4_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(N__18408),
            .in2(N__16916),
            .in3(N__16805),
            .lcout(\POWERLED.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_4_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_4_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_4_12_5  (
            .in0(N__16781),
            .in1(N__16904),
            .in2(N__16877),
            .in3(N__16796),
            .lcout(\POWERLED.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_4_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_4_12_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_4_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16895),
            .in3(N__16793),
            .lcout(\POWERLED.mult1_un110_sum_s_8 ),
            .ltout(\POWERLED.mult1_un110_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_12_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16940),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un110_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_4_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_4_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__21758),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\POWERLED.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_4_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_4_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__18437),
            .in2(N__18427),
            .in3(N__16928),
            .lcout(\POWERLED.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_4_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_4_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__18423),
            .in2(N__18329),
            .in3(N__16919),
            .lcout(\POWERLED.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_4_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_4_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__18317),
            .in2(N__18508),
            .in3(N__16907),
            .lcout(\POWERLED.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_4_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_4_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__18504),
            .in2(N__18548),
            .in3(N__16898),
            .lcout(\POWERLED.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_4_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_4_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_4_13_5  (
            .in0(N__18404),
            .in1(N__18536),
            .in2(N__18428),
            .in3(N__16886),
            .lcout(\POWERLED.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_4_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_4_13_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18527),
            .in3(N__16883),
            .lcout(\POWERLED.mult1_un103_sum_s_8 ),
            .ltout(\POWERLED.mult1_un103_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_4_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_4_13_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16880),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_4_14_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_4_14_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_4_14_0  (
            .in0(N__17261),
            .in1(N__18290),
            .in2(N__17231),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_cry_0_i ),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_4_14_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_4_14_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_4_14_1  (
            .in0(N__17222),
            .in1(N__18443),
            .in2(N__17195),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5036_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_0 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_4_14_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_4_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__18281),
            .in2(N__17150),
            .in3(N__17183),
            .lcout(\POWERLED.N_5037_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_1 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_4_14_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_4_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__18272),
            .in2(N__17111),
            .in3(N__17141),
            .lcout(\POWERLED.N_5038_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_2 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_4_14_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_4_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__18449),
            .in2(N__17075),
            .in3(N__17102),
            .lcout(\POWERLED.N_5039_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_3 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_4_14_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_4_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_4_14_5  (
            .in0(_gnd_net_),
            .in1(N__18476),
            .in2(N__17033),
            .in3(N__17066),
            .lcout(\POWERLED.N_5040_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_4 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_4_14_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_4_14_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_4_14_6  (
            .in0(N__17024),
            .in1(N__18335),
            .in2(N__16994),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5041_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_5 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_4_14_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_4_14_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_4_14_7  (
            .in0(N__16982),
            .in1(N__16958),
            .in2(N__16949),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5042_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_6 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_4_15_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_4_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__17507),
            .in2(N__17546),
            .in3(N__17534),
            .lcout(\POWERLED.N_5043_i ),
            .ltout(),
            .carryin(bfn_4_15_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_4_15_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_4_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__17474),
            .in2(N__18386),
            .in3(N__17501),
            .lcout(\POWERLED.N_5044_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_8 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_4_15_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_4_15_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_4_15_2  (
            .in0(N__17468),
            .in1(N__17420),
            .in2(N__17435),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5045_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_9 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_4_15_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_4_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(N__17573),
            .in2(N__17384),
            .in3(N__17414),
            .lcout(\POWERLED.N_5046_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_10 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_4_15_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_4_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__18557),
            .in2(N__17345),
            .in3(N__17375),
            .lcout(\POWERLED.N_5047_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_11 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_4_15_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_4_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__17303),
            .in2(N__18593),
            .in3(N__17333),
            .lcout(\POWERLED.N_5048_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_12 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_4_15_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_4_15_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_4_15_6  (
            .in0(N__17297),
            .in1(N__17267),
            .in2(N__17567),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5049_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_13 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_4_15_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_4_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(N__20366),
            .in2(N__17621),
            .in3(N__17648),
            .lcout(\POWERLED.N_5050_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_14 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_16_0 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17612),
            .lcout(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_16_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18637),
            .lcout(\POWERLED.mult1_un89_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_16_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20603),
            .lcout(\POWERLED.mult1_un68_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_0_c_LC_5_1_0 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_0_c_LC_5_1_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_0_c_LC_5_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_0_c_LC_5_1_0  (
            .in0(_gnd_net_),
            .in1(N__19259),
            .in2(N__19163),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_1_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_1_LC_5_1_1 .C_ON=1'b1;
    defparam \HDA_STRAP.count_1_LC_5_1_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_1_LC_5_1_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_1_LC_5_1_1  (
            .in0(_gnd_net_),
            .in1(N__19273),
            .in2(_gnd_net_),
            .in3(N__17558),
            .lcout(\HDA_STRAP.countZ0Z_1 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_0 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_1 ),
            .clk(N__32053),
            .ce(N__25309),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_2_LC_5_1_2 .C_ON=1'b1;
    defparam \HDA_STRAP.count_2_LC_5_1_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_2_LC_5_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_2_LC_5_1_2  (
            .in0(_gnd_net_),
            .in1(N__18829),
            .in2(_gnd_net_),
            .in3(N__17555),
            .lcout(\HDA_STRAP.countZ0Z_2 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_1 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_2 ),
            .clk(N__32053),
            .ce(N__25309),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_3_LC_5_1_3 .C_ON=1'b1;
    defparam \HDA_STRAP.count_3_LC_5_1_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_3_LC_5_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_3_LC_5_1_3  (
            .in0(_gnd_net_),
            .in1(N__18814),
            .in2(_gnd_net_),
            .in3(N__17552),
            .lcout(\HDA_STRAP.countZ0Z_3 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_2 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_3 ),
            .clk(N__32053),
            .ce(N__25309),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_4_LC_5_1_4 .C_ON=1'b1;
    defparam \HDA_STRAP.count_4_LC_5_1_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_4_LC_5_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_4_LC_5_1_4  (
            .in0(_gnd_net_),
            .in1(N__18842),
            .in2(_gnd_net_),
            .in3(N__17549),
            .lcout(\HDA_STRAP.countZ0Z_4 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_3 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_4 ),
            .clk(N__32053),
            .ce(N__25309),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_5_LC_5_1_5 .C_ON=1'b1;
    defparam \HDA_STRAP.count_5_LC_5_1_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_5_LC_5_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_5_LC_5_1_5  (
            .in0(_gnd_net_),
            .in1(N__18803),
            .in2(_gnd_net_),
            .in3(N__17699),
            .lcout(\HDA_STRAP.countZ0Z_5 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_4 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_5 ),
            .clk(N__32053),
            .ce(N__25309),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_5_1_6 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_5_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_5_1_6  (
            .in0(_gnd_net_),
            .in1(N__18873),
            .in2(_gnd_net_),
            .in3(N__17690),
            .lcout(\HDA_STRAP.un1_count_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_5 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_7_LC_5_1_7 .C_ON=1'b1;
    defparam \HDA_STRAP.count_7_LC_5_1_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_7_LC_5_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_7_LC_5_1_7  (
            .in0(_gnd_net_),
            .in1(N__18692),
            .in2(_gnd_net_),
            .in3(N__17687),
            .lcout(\HDA_STRAP.countZ0Z_7 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_6 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_7 ),
            .clk(N__32053),
            .ce(N__25309),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_5_2_0 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_5_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_5_2_0  (
            .in0(_gnd_net_),
            .in1(N__18911),
            .in2(_gnd_net_),
            .in3(N__17678),
            .lcout(\HDA_STRAP.un1_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_5_2_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_9_LC_5_2_1 .C_ON=1'b1;
    defparam \HDA_STRAP.count_9_LC_5_2_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_9_LC_5_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_9_LC_5_2_1  (
            .in0(_gnd_net_),
            .in1(N__18731),
            .in2(_gnd_net_),
            .in3(N__17675),
            .lcout(\HDA_STRAP.countZ0Z_9 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_8 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_9 ),
            .clk(N__32220),
            .ce(N__25315),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_5_2_2 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_5_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_5_2_2  (
            .in0(_gnd_net_),
            .in1(N__18765),
            .in2(_gnd_net_),
            .in3(N__17666),
            .lcout(\HDA_STRAP.un1_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_9 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_5_2_3 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_5_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_5_2_3  (
            .in0(_gnd_net_),
            .in1(N__18791),
            .in2(_gnd_net_),
            .in3(N__17657),
            .lcout(\HDA_STRAP.un1_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_10 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_12_LC_5_2_4 .C_ON=1'b1;
    defparam \HDA_STRAP.count_12_LC_5_2_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_12_LC_5_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_12_LC_5_2_4  (
            .in0(_gnd_net_),
            .in1(N__18719),
            .in2(_gnd_net_),
            .in3(N__17654),
            .lcout(\HDA_STRAP.countZ0Z_12 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_11 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_12 ),
            .clk(N__32220),
            .ce(N__25315),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_13_LC_5_2_5 .C_ON=1'b1;
    defparam \HDA_STRAP.count_13_LC_5_2_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_13_LC_5_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_13_LC_5_2_5  (
            .in0(_gnd_net_),
            .in1(N__18706),
            .in2(_gnd_net_),
            .in3(N__17651),
            .lcout(\HDA_STRAP.countZ0Z_13 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_12 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_13 ),
            .clk(N__32220),
            .ce(N__25315),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_14_LC_5_2_6 .C_ON=1'b1;
    defparam \HDA_STRAP.count_14_LC_5_2_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_14_LC_5_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_14_LC_5_2_6  (
            .in0(_gnd_net_),
            .in1(N__18890),
            .in2(_gnd_net_),
            .in3(N__17711),
            .lcout(\HDA_STRAP.countZ0Z_14 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_13 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_14 ),
            .clk(N__32220),
            .ce(N__25315),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_15_LC_5_2_7 .C_ON=1'b1;
    defparam \HDA_STRAP.count_15_LC_5_2_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_15_LC_5_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_15_LC_5_2_7  (
            .in0(_gnd_net_),
            .in1(N__18854),
            .in2(_gnd_net_),
            .in3(N__17708),
            .lcout(\HDA_STRAP.countZ0Z_15 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_14 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_15 ),
            .clk(N__32220),
            .ce(N__25315),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_5_3_0 .C_ON=1'b1;
    defparam \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_5_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(N__19076),
            .in2(_gnd_net_),
            .in3(N__17705),
            .lcout(\HDA_STRAP.un1_count_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_17_LC_5_3_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_17_LC_5_3_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_17_LC_5_3_1 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \HDA_STRAP.count_17_LC_5_3_1  (
            .in0(N__19140),
            .in1(N__19234),
            .in2(N__19212),
            .in3(N__17702),
            .lcout(\HDA_STRAP.countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32226),
            .ce(N__25312),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_0_LC_5_4_0 .C_ON=1'b0;
    defparam \COUNTER.counter_0_LC_5_4_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_0_LC_5_4_0 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \COUNTER.counter_0_LC_5_4_0  (
            .in0(N__19059),
            .in1(_gnd_net_),
            .in2(N__22550),
            .in3(_gnd_net_),
            .lcout(\COUNTER.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32471),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_5_LC_5_4_2 .C_ON=1'b0;
    defparam \COUNTER.counter_5_LC_5_4_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_5_LC_5_4_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \COUNTER.counter_5_LC_5_4_2  (
            .in0(N__22543),
            .in1(N__18920),
            .in2(_gnd_net_),
            .in3(N__18934),
            .lcout(\COUNTER.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32471),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_2_LC_5_4_3 .C_ON=1'b0;
    defparam \COUNTER.counter_2_LC_5_4_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_2_LC_5_4_3 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_2_LC_5_4_3  (
            .in0(N__19014),
            .in1(N__18998),
            .in2(_gnd_net_),
            .in3(N__22547),
            .lcout(\COUNTER.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32471),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_RNO_LC_5_4_4 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_5_4_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_2_c_RNO_LC_5_4_4  (
            .in0(N__19321),
            .in1(N__19354),
            .in2(N__19340),
            .in3(N__19369),
            .lcout(\COUNTER.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_RNO_LC_5_4_5 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_5_4_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_RNO_LC_5_4_5  (
            .in0(N__18984),
            .in1(N__18957),
            .in2(N__19016),
            .in3(N__19058),
            .lcout(\COUNTER.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_RNO_LC_5_4_6 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_5_4_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \COUNTER.un4_counter_1_c_RNO_LC_5_4_6  (
            .in0(N__19384),
            .in1(N__19410),
            .in2(N__19039),
            .in3(N__18933),
            .lcout(\COUNTER.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_4_LC_5_4_7 .C_ON=1'b0;
    defparam \COUNTER.counter_4_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_4_LC_5_4_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_4_LC_5_4_7  (
            .in0(N__18944),
            .in1(N__18958),
            .in2(_gnd_net_),
            .in3(N__22548),
            .lcout(\COUNTER.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32471),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_5_5_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_5_5_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RSMRST_PWRGD.count_esr_RNO_0_15_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(N__20945),
            .in2(_gnd_net_),
            .in3(N__25402),
            .lcout(\RSMRST_PWRGD.N_92_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_RNO_LC_5_5_2 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_5_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_3_c_RNO_LC_5_5_2  (
            .in0(N__19465),
            .in1(N__19288),
            .in2(N__19307),
            .in3(N__19450),
            .lcout(\COUNTER.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_LC_5_5_4 .C_ON=1'b0;
    defparam \COUNTER.counter_1_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_1_LC_5_5_4 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \COUNTER.counter_1_LC_5_5_4  (
            .in0(N__19038),
            .in1(N__22538),
            .in2(_gnd_net_),
            .in3(N__19061),
            .lcout(\COUNTER.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32228),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_3_LC_5_5_6 .C_ON=1'b0;
    defparam \COUNTER.counter_3_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_3_LC_5_5_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_3_LC_5_5_6  (
            .in0(N__18968),
            .in1(N__18986),
            .in2(_gnd_net_),
            .in3(N__22539),
            .lcout(\COUNTER.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32228),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_6_LC_5_5_7 .C_ON=1'b0;
    defparam \COUNTER.counter_6_LC_5_5_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_6_LC_5_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \COUNTER.counter_6_LC_5_5_7  (
            .in0(N__22537),
            .in1(N__19394),
            .in2(_gnd_net_),
            .in3(N__19414),
            .lcout(\COUNTER.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32228),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_RNO_LC_5_6_6 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_5_6_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_6_c_RNO_LC_5_6_6  (
            .in0(N__19603),
            .in1(N__19555),
            .in2(N__19574),
            .in3(N__19588),
            .lcout(\COUNTER.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_5_6_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_5_6_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_5_6_7  (
            .in0(N__26805),
            .in1(N__21195),
            .in2(_gnd_net_),
            .in3(N__21169),
            .lcout(N_555),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_3_LC_5_7_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_3_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_3_LC_5_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_3_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17768),
            .lcout(\VPP_VDDQ.count_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32283),
            .ce(N__19780),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_5_LC_5_7_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_5_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_5_LC_5_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_5_LC_5_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17750),
            .lcout(\VPP_VDDQ.count_2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32283),
            .ce(N__19780),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_8_LC_5_7_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_8_LC_5_7_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_8_LC_5_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_8_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18028),
            .lcout(\VPP_VDDQ.count_2_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32283),
            .ce(N__19780),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_10_LC_5_7_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_10_LC_5_7_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_10_LC_5_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_10_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17975),
            .lcout(\VPP_VDDQ.count_2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32283),
            .ce(N__19780),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_5_8_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_5_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(N__17822),
            .in2(N__17795),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_5_8_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_5_8_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_5_8_1  (
            .in0(N__18193),
            .in1(N__19685),
            .in2(_gnd_net_),
            .in3(N__17771),
            .lcout(\VPP_VDDQ.count_2_1_2 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_5_8_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_5_8_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_5_8_2  (
            .in0(N__18201),
            .in1(N__19630),
            .in2(_gnd_net_),
            .in3(N__17756),
            .lcout(\VPP_VDDQ.count_2_1_3 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_5_8_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_5_8_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_5_8_3  (
            .in0(N__18194),
            .in1(N__19859),
            .in2(_gnd_net_),
            .in3(N__17753),
            .lcout(\VPP_VDDQ.count_2_1_4 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_5_8_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_5_8_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_5_8_4  (
            .in0(N__18202),
            .in1(N__19672),
            .in2(_gnd_net_),
            .in3(N__17738),
            .lcout(\VPP_VDDQ.count_2_1_5 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIDNMU_LC_5_8_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIDNMU_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIDNMU_LC_5_8_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIDNMU_LC_5_8_5  (
            .in0(N__18195),
            .in1(N__19880),
            .in2(_gnd_net_),
            .in3(N__17735),
            .lcout(\VPP_VDDQ.count_2_1_6 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_5_8_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_5_8_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_5_8_6  (
            .in0(N__18203),
            .in1(N__18059),
            .in2(_gnd_net_),
            .in3(N__18032),
            .lcout(\VPP_VDDQ.count_2_1_7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_5_8_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_5_8_7 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_5_8_7  (
            .in0(N__18196),
            .in1(_gnd_net_),
            .in2(N__19657),
            .in3(N__18017),
            .lcout(\VPP_VDDQ.count_2_1_8 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_5_9_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_5_9_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_5_9_0  (
            .in0(N__18205),
            .in1(N__18014),
            .in2(_gnd_net_),
            .in3(N__17993),
            .lcout(\VPP_VDDQ.count_2_1_9 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_5_9_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_5_9_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_5_9_1  (
            .in0(N__18197),
            .in1(N__17986),
            .in2(_gnd_net_),
            .in3(N__17960),
            .lcout(\VPP_VDDQ.count_2_1_10 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_5_9_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_5_9_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_5_9_2  (
            .in0(N__18204),
            .in1(N__17957),
            .in2(_gnd_net_),
            .in3(N__17927),
            .lcout(\VPP_VDDQ.count_2_1_11 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_5_9_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_5_9_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_5_9_3  (
            .in0(N__18198),
            .in1(N__17924),
            .in2(_gnd_net_),
            .in3(N__17903),
            .lcout(\VPP_VDDQ.count_2_1_12 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_5_9_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_5_9_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_5_9_4  (
            .in0(N__18206),
            .in1(N__17899),
            .in2(_gnd_net_),
            .in3(N__17876),
            .lcout(\VPP_VDDQ.count_2_1_13 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_5_9_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_5_9_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_5_9_5  (
            .in0(N__18199),
            .in1(N__17873),
            .in2(_gnd_net_),
            .in3(N__17852),
            .lcout(\VPP_VDDQ.count_2_1_14 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_5_9_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_5_9_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_5_9_6  (
            .in0(N__18218),
            .in1(N__18200),
            .in2(_gnd_net_),
            .in3(N__18125),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_15_LC_5_9_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_15_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_15_LC_5_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_15_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18122),
            .lcout(\VPP_VDDQ.count_2_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32350),
            .ce(N__19781),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_5_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_5_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__21551),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\POWERLED.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_5_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_5_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__20387),
            .in2(N__18261),
            .in3(N__18104),
            .lcout(\POWERLED.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_5_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_5_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__18101),
            .in2(N__18263),
            .in3(N__18095),
            .lcout(\POWERLED.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_5_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_5_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__18092),
            .in2(N__18373),
            .in3(N__18086),
            .lcout(\POWERLED.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_5_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_5_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__18083),
            .in2(N__18372),
            .in3(N__18077),
            .lcout(\POWERLED.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_5_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_5_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_5_10_5  (
            .in0(N__20062),
            .in1(N__18074),
            .in2(N__18262),
            .in3(N__18068),
            .lcout(\POWERLED.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_5_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_5_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_5_10_6  (
            .in0(N__18065),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18266),
            .lcout(\POWERLED.mult1_un131_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18361),
            .lcout(\POWERLED.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__21587),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\POWERLED.mult1_un145_sum_cry_2_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__19890),
            .in2(N__20183),
            .in3(N__18239),
            .lcout(\POWERLED.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_2_c ),
            .carryout(\POWERLED.mult1_un145_sum_cry_3_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__20015),
            .in2(N__19895),
            .in3(N__18236),
            .lcout(\POWERLED.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_3_c ),
            .carryout(\POWERLED.mult1_un145_sum_cry_4_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__19917),
            .in2(N__20000),
            .in3(N__18233),
            .lcout(\POWERLED.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_4_c ),
            .carryout(\POWERLED.mult1_un145_sum_cry_5_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__19979),
            .in2(N__19924),
            .in3(N__18230),
            .lcout(\POWERLED.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_5_c ),
            .carryout(\POWERLED.mult1_un145_sum_cry_6_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_11_5  (
            .in0(N__20132),
            .in1(N__19894),
            .in2(N__19964),
            .in3(N__18227),
            .lcout(\POWERLED.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_6_c ),
            .carryout(\POWERLED.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_11_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_11_6  (
            .in0(N__19946),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18224),
            .lcout(\POWERLED.mult1_un145_sum_s_8 ),
            .ltout(\POWERLED.mult1_un145_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18221),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_5_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_5_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(N__26558),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(\POWERLED.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_5_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_5_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__22754),
            .in2(N__18310),
            .in3(N__20258),
            .lcout(G_2150),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_0 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_5_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_5_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__18306),
            .in2(N__20351),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_5_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_5_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__20259),
            .in2(N__20333),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_5_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_5_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__20315),
            .in2(N__20266),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_5_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_5_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(N__20300),
            .in2(N__18311),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_5_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_5_12_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_5_12_6  (
            .in0(N__20285),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18293),
            .lcout(\POWERLED.un85_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20235),
            .lcout(\POWERLED.un85_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_13_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20141),
            .lcout(\POWERLED.un85_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_13_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19928),
            .lcout(\POWERLED.mult1_un138_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_5_13_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_5_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20267),
            .lcout(\POWERLED.un85_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_5_13_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_5_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21739),
            .lcout(\POWERLED.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_5_13_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_5_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18499),
            .lcout(\POWERLED.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18409),
            .lcout(\POWERLED.mult1_un103_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_13_7  (
            .in0(N__18374),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un124_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__21740),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\POWERLED.mult1_un96_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__18566),
            .in2(N__18610),
            .in3(N__18320),
            .lcout(\POWERLED.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__18606),
            .in2(N__18470),
            .in3(N__18551),
            .lcout(\POWERLED.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(N__18458),
            .in2(N__18638),
            .in3(N__18539),
            .lcout(\POWERLED.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__18636),
            .in2(N__18674),
            .in3(N__18530),
            .lcout(\POWERLED.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_14_5  (
            .in0(N__18500),
            .in1(N__18662),
            .in2(N__18611),
            .in3(N__18518),
            .lcout(\POWERLED.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_14_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18653),
            .in3(N__18515),
            .lcout(\POWERLED.mult1_un96_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_14_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_14_7  (
            .in0(N__20072),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un131_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__21715),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\POWERLED.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__21788),
            .in2(N__18583),
            .in3(N__18461),
            .lcout(\POWERLED.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__18579),
            .in2(N__20519),
            .in3(N__18452),
            .lcout(\POWERLED.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__20498),
            .in2(N__20654),
            .in3(N__18665),
            .lcout(\POWERLED.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(N__20653),
            .in2(N__20483),
            .in3(N__18656),
            .lcout(\POWERLED.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_15_5  (
            .in0(N__18632),
            .in1(N__20711),
            .in2(N__18584),
            .in3(N__18644),
            .lcout(\POWERLED.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_15_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20678),
            .in3(N__18641),
            .lcout(\POWERLED.mult1_un89_sum_s_8 ),
            .ltout(\POWERLED.mult1_un89_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_15_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18614),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_5_16_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_5_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_5_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20743),
            .lcout(\POWERLED.mult1_un75_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_16_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20647),
            .lcout(\POWERLED.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_5_16_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_5_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_5_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21716),
            .lcout(\POWERLED.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_5_16_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_5_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_5_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20648),
            .lcout(\POWERLED.mult1_un82_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_5_LC_6_1_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_5_LC_6_1_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_5_LC_6_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_5_LC_6_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21977),
            .lcout(\POWERLED.count_off_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31836),
            .ce(N__23545),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_6_LC_6_1_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_6_LC_6_1_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_6_LC_6_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_6_LC_6_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22052),
            .lcout(\POWERLED.count_off_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31836),
            .ce(N__23545),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_6_2_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_6_2_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \HDA_STRAP.count_RNIDLB61_6_LC_6_2_1  (
            .in0(N__18910),
            .in1(N__18889),
            .in2(N__18878),
            .in3(N__18853),
            .lcout(\HDA_STRAP.un4_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI2L821_2_LC_6_2_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI2L821_2_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI2L821_2_LC_6_2_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \HDA_STRAP.count_RNI2L821_2_LC_6_2_3  (
            .in0(N__18841),
            .in1(N__18830),
            .in2(N__18818),
            .in3(N__18802),
            .lcout(\HDA_STRAP.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIH7IR1_10_LC_6_2_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIH7IR1_10_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIH7IR1_10_LC_6_2_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \HDA_STRAP.count_RNIH7IR1_10_LC_6_2_4  (
            .in0(N__18790),
            .in1(N__18767),
            .in2(_gnd_net_),
            .in3(N__19220),
            .lcout(),
            .ltout(\HDA_STRAP.un4_count_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_6_2_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_6_2_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_6_2_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \HDA_STRAP.count_RNIB5IA5_2_LC_6_2_5  (
            .in0(N__18746),
            .in1(N__18680),
            .in2(N__18740),
            .in3(N__18737),
            .lcout(\HDA_STRAP.un4_count ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_6_2_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_6_2_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \HDA_STRAP.count_RNIBJB61_7_LC_6_2_6  (
            .in0(N__18730),
            .in1(N__18718),
            .in2(N__18707),
            .in3(N__18691),
            .lcout(\HDA_STRAP.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_0_LC_6_3_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_0_LC_6_3_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_0_LC_6_3_1 .LUT_INIT=16'b0000011001100110;
    LogicCell40 \HDA_STRAP.count_0_LC_6_3_1  (
            .in0(N__19254),
            .in1(N__19150),
            .in2(N__19160),
            .in3(N__19198),
            .lcout(\HDA_STRAP.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32225),
            .ce(N__25313),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_RNO_LC_6_3_2 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_6_3_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_7_c_RNO_LC_6_3_2  (
            .in0(N__19502),
            .in1(N__19481),
            .in2(N__19541),
            .in3(N__19520),
            .lcout(\COUNTER.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_6_3_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_6_3_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \HDA_STRAP.count_RNI4CB61_17_LC_6_3_3  (
            .in0(N__19074),
            .in1(N__19274),
            .in2(N__19258),
            .in3(N__19235),
            .lcout(\HDA_STRAP.un4_count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_16_LC_6_3_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_16_LC_6_3_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_16_LC_6_3_6 .LUT_INIT=16'b0000011101110000;
    LogicCell40 \HDA_STRAP.count_16_LC_6_3_6  (
            .in0(N__19197),
            .in1(N__19146),
            .in2(N__19085),
            .in3(N__19075),
            .lcout(\HDA_STRAP.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32225),
            .ce(N__25313),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_c_LC_6_4_0 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_c_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_c_LC_6_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.counter_1_cry_1_c_LC_6_4_0  (
            .in0(_gnd_net_),
            .in1(N__19060),
            .in2(N__19040),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(\COUNTER.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_6_4_1 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_6_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_6_4_1  (
            .in0(_gnd_net_),
            .in1(N__19015),
            .in2(_gnd_net_),
            .in3(N__18989),
            .lcout(\COUNTER.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_1 ),
            .carryout(\COUNTER.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_6_4_2 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_6_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_6_4_2  (
            .in0(_gnd_net_),
            .in1(N__18985),
            .in2(_gnd_net_),
            .in3(N__18962),
            .lcout(\COUNTER.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_2 ),
            .carryout(\COUNTER.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_6_4_3 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_6_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_6_4_3  (
            .in0(_gnd_net_),
            .in1(N__18959),
            .in2(_gnd_net_),
            .in3(N__18938),
            .lcout(\COUNTER.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_3 ),
            .carryout(\COUNTER.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_6_4_4 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_6_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_6_4_4  (
            .in0(_gnd_net_),
            .in1(N__18935),
            .in2(_gnd_net_),
            .in3(N__18914),
            .lcout(\COUNTER.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_4 ),
            .carryout(\COUNTER.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_6_4_5 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_6_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_6_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19415),
            .in3(N__19388),
            .lcout(\COUNTER.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_5 ),
            .carryout(\COUNTER.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_7_LC_6_4_6 .C_ON=1'b1;
    defparam \COUNTER.counter_7_LC_6_4_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_7_LC_6_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_7_LC_6_4_6  (
            .in0(_gnd_net_),
            .in1(N__19385),
            .in2(_gnd_net_),
            .in3(N__19373),
            .lcout(\COUNTER.counterZ0Z_7 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_6 ),
            .carryout(\COUNTER.counter_1_cry_7 ),
            .clk(N__32224),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_8_LC_6_4_7 .C_ON=1'b1;
    defparam \COUNTER.counter_8_LC_6_4_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_8_LC_6_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_8_LC_6_4_7  (
            .in0(_gnd_net_),
            .in1(N__19370),
            .in2(_gnd_net_),
            .in3(N__19358),
            .lcout(\COUNTER.counterZ0Z_8 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_7 ),
            .carryout(\COUNTER.counter_1_cry_8 ),
            .clk(N__32224),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_9_LC_6_5_0 .C_ON=1'b1;
    defparam \COUNTER.counter_9_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_9_LC_6_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_9_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(N__19355),
            .in2(_gnd_net_),
            .in3(N__19343),
            .lcout(\COUNTER.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_6_5_0_),
            .carryout(\COUNTER.counter_1_cry_9 ),
            .clk(N__32227),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_10_LC_6_5_1 .C_ON=1'b1;
    defparam \COUNTER.counter_10_LC_6_5_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_10_LC_6_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_10_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(N__19339),
            .in2(_gnd_net_),
            .in3(N__19325),
            .lcout(\COUNTER.counterZ0Z_10 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_9 ),
            .carryout(\COUNTER.counter_1_cry_10 ),
            .clk(N__32227),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_11_LC_6_5_2 .C_ON=1'b1;
    defparam \COUNTER.counter_11_LC_6_5_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_11_LC_6_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_11_LC_6_5_2  (
            .in0(_gnd_net_),
            .in1(N__19322),
            .in2(_gnd_net_),
            .in3(N__19310),
            .lcout(\COUNTER.counterZ0Z_11 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_10 ),
            .carryout(\COUNTER.counter_1_cry_11 ),
            .clk(N__32227),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_12_LC_6_5_3 .C_ON=1'b1;
    defparam \COUNTER.counter_12_LC_6_5_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_12_LC_6_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_12_LC_6_5_3  (
            .in0(_gnd_net_),
            .in1(N__19306),
            .in2(_gnd_net_),
            .in3(N__19292),
            .lcout(\COUNTER.counterZ0Z_12 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_11 ),
            .carryout(\COUNTER.counter_1_cry_12 ),
            .clk(N__32227),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_13_LC_6_5_4 .C_ON=1'b1;
    defparam \COUNTER.counter_13_LC_6_5_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_13_LC_6_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_13_LC_6_5_4  (
            .in0(_gnd_net_),
            .in1(N__19289),
            .in2(_gnd_net_),
            .in3(N__19277),
            .lcout(\COUNTER.counterZ0Z_13 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_12 ),
            .carryout(\COUNTER.counter_1_cry_13 ),
            .clk(N__32227),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_14_LC_6_5_5 .C_ON=1'b1;
    defparam \COUNTER.counter_14_LC_6_5_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_14_LC_6_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_14_LC_6_5_5  (
            .in0(_gnd_net_),
            .in1(N__19466),
            .in2(_gnd_net_),
            .in3(N__19454),
            .lcout(\COUNTER.counterZ0Z_14 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_13 ),
            .carryout(\COUNTER.counter_1_cry_14 ),
            .clk(N__32227),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_15_LC_6_5_6 .C_ON=1'b1;
    defparam \COUNTER.counter_15_LC_6_5_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_15_LC_6_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_15_LC_6_5_6  (
            .in0(_gnd_net_),
            .in1(N__19451),
            .in2(_gnd_net_),
            .in3(N__19439),
            .lcout(\COUNTER.counterZ0Z_15 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_14 ),
            .carryout(\COUNTER.counter_1_cry_15 ),
            .clk(N__32227),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_16_LC_6_5_7 .C_ON=1'b1;
    defparam \COUNTER.counter_16_LC_6_5_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_16_LC_6_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_16_LC_6_5_7  (
            .in0(_gnd_net_),
            .in1(N__21035),
            .in2(_gnd_net_),
            .in3(N__19436),
            .lcout(\COUNTER.counterZ0Z_16 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_15 ),
            .carryout(\COUNTER.counter_1_cry_16 ),
            .clk(N__32227),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_17_LC_6_6_0 .C_ON=1'b1;
    defparam \COUNTER.counter_17_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_17_LC_6_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_17_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__21062),
            .in2(_gnd_net_),
            .in3(N__19433),
            .lcout(\COUNTER.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(\COUNTER.counter_1_cry_17 ),
            .clk(N__32180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_18_LC_6_6_1 .C_ON=1'b1;
    defparam \COUNTER.counter_18_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_18_LC_6_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_18_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__21049),
            .in2(_gnd_net_),
            .in3(N__19430),
            .lcout(\COUNTER.counterZ0Z_18 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_17 ),
            .carryout(\COUNTER.counter_1_cry_18 ),
            .clk(N__32180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_19_LC_6_6_2 .C_ON=1'b1;
    defparam \COUNTER.counter_19_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_19_LC_6_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_19_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__21074),
            .in2(_gnd_net_),
            .in3(N__19427),
            .lcout(\COUNTER.counterZ0Z_19 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_18 ),
            .carryout(\COUNTER.counter_1_cry_19 ),
            .clk(N__32180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_20_LC_6_6_3 .C_ON=1'b1;
    defparam \COUNTER.counter_20_LC_6_6_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_20_LC_6_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_20_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__21011),
            .in2(_gnd_net_),
            .in3(N__19424),
            .lcout(\COUNTER.counterZ0Z_20 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_19 ),
            .carryout(\COUNTER.counter_1_cry_20 ),
            .clk(N__32180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_21_LC_6_6_4 .C_ON=1'b1;
    defparam \COUNTER.counter_21_LC_6_6_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_21_LC_6_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_21_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(N__20998),
            .in2(_gnd_net_),
            .in3(N__19421),
            .lcout(\COUNTER.counterZ0Z_21 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_20 ),
            .carryout(\COUNTER.counter_1_cry_21 ),
            .clk(N__32180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_22_LC_6_6_5 .C_ON=1'b1;
    defparam \COUNTER.counter_22_LC_6_6_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_22_LC_6_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_22_LC_6_6_5  (
            .in0(_gnd_net_),
            .in1(N__20984),
            .in2(_gnd_net_),
            .in3(N__19418),
            .lcout(\COUNTER.counterZ0Z_22 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_21 ),
            .carryout(\COUNTER.counter_1_cry_22 ),
            .clk(N__32180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_23_LC_6_6_6 .C_ON=1'b1;
    defparam \COUNTER.counter_23_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_23_LC_6_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_23_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(N__21023),
            .in2(_gnd_net_),
            .in3(N__19607),
            .lcout(\COUNTER.counterZ0Z_23 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_22 ),
            .carryout(\COUNTER.counter_1_cry_23 ),
            .clk(N__32180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_24_LC_6_6_7 .C_ON=1'b1;
    defparam \COUNTER.counter_24_LC_6_6_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_24_LC_6_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_24_LC_6_6_7  (
            .in0(_gnd_net_),
            .in1(N__19604),
            .in2(_gnd_net_),
            .in3(N__19592),
            .lcout(\COUNTER.counterZ0Z_24 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_23 ),
            .carryout(\COUNTER.counter_1_cry_24 ),
            .clk(N__32180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_25_LC_6_7_0 .C_ON=1'b1;
    defparam \COUNTER.counter_25_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_25_LC_6_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_25_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(N__19589),
            .in2(_gnd_net_),
            .in3(N__19577),
            .lcout(\COUNTER.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(\COUNTER.counter_1_cry_25 ),
            .clk(N__32052),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_26_LC_6_7_1 .C_ON=1'b1;
    defparam \COUNTER.counter_26_LC_6_7_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_26_LC_6_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_26_LC_6_7_1  (
            .in0(_gnd_net_),
            .in1(N__19573),
            .in2(_gnd_net_),
            .in3(N__19559),
            .lcout(\COUNTER.counterZ0Z_26 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_25 ),
            .carryout(\COUNTER.counter_1_cry_26 ),
            .clk(N__32052),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_27_LC_6_7_2 .C_ON=1'b1;
    defparam \COUNTER.counter_27_LC_6_7_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_27_LC_6_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_27_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(N__19556),
            .in2(_gnd_net_),
            .in3(N__19544),
            .lcout(\COUNTER.counterZ0Z_27 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_26 ),
            .carryout(\COUNTER.counter_1_cry_27 ),
            .clk(N__32052),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_28_LC_6_7_3 .C_ON=1'b1;
    defparam \COUNTER.counter_28_LC_6_7_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_28_LC_6_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_28_LC_6_7_3  (
            .in0(_gnd_net_),
            .in1(N__19537),
            .in2(_gnd_net_),
            .in3(N__19523),
            .lcout(\COUNTER.counterZ0Z_28 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_27 ),
            .carryout(\COUNTER.counter_1_cry_28 ),
            .clk(N__32052),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_29_LC_6_7_4 .C_ON=1'b1;
    defparam \COUNTER.counter_29_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_29_LC_6_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_29_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(N__19519),
            .in2(_gnd_net_),
            .in3(N__19505),
            .lcout(\COUNTER.counterZ0Z_29 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_28 ),
            .carryout(\COUNTER.counter_1_cry_29 ),
            .clk(N__32052),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_30_LC_6_7_5 .C_ON=1'b1;
    defparam \COUNTER.counter_30_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_30_LC_6_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_30_LC_6_7_5  (
            .in0(_gnd_net_),
            .in1(N__19501),
            .in2(_gnd_net_),
            .in3(N__19487),
            .lcout(\COUNTER.counterZ0Z_30 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_29 ),
            .carryout(\COUNTER.counter_1_cry_30 ),
            .clk(N__32052),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_31_LC_6_7_6 .C_ON=1'b0;
    defparam \COUNTER.counter_31_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_31_LC_6_7_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.counter_31_LC_6_7_6  (
            .in0(_gnd_net_),
            .in1(N__19480),
            .in2(_gnd_net_),
            .in3(N__19484),
            .lcout(\COUNTER.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32052),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_4_LC_6_8_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_4_LC_6_8_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_4_LC_6_8_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_2_4_LC_6_8_0  (
            .in0(N__19868),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32206),
            .ce(N__19798),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_6_LC_6_8_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_6_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_6_LC_6_8_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_2_6_LC_6_8_1  (
            .in0(N__19840),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32206),
            .ce(N__19798),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIREAN_6_LC_6_8_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIREAN_6_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIREAN_6_LC_6_8_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.count_2_RNIREAN_6_LC_6_8_2  (
            .in0(N__19852),
            .in1(N__19784),
            .in2(_gnd_net_),
            .in3(N__19839),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI9HKU_4_LC_6_8_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI9HKU_4_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI9HKU_4_LC_6_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_2_RNI9HKU_4_LC_6_8_3  (
            .in0(N__19783),
            .in1(N__19874),
            .in2(_gnd_net_),
            .in3(N__19867),
            .lcout(\VPP_VDDQ.count_2Z0Z_4 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIREAN_0_6_LC_6_8_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIREAN_0_6_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIREAN_0_6_LC_6_8_4 .LUT_INIT=16'b0000000100001101;
    LogicCell40 \VPP_VDDQ.count_2_RNIREAN_0_6_LC_6_8_4  (
            .in0(N__19853),
            .in1(N__19785),
            .in2(N__19844),
            .in3(N__19841),
            .lcout(\VPP_VDDQ.un9_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_2_LC_6_8_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_2_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_2_LC_6_8_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_2_2_LC_6_8_5  (
            .in0(N__19811),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32206),
            .ce(N__19798),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI5BIU_2_LC_6_8_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI5BIU_2_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI5BIU_2_LC_6_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNI5BIU_2_LC_6_8_6  (
            .in0(N__19817),
            .in1(N__19810),
            .in2(_gnd_net_),
            .in3(N__19782),
            .lcout(\VPP_VDDQ.count_2Z0Z_2 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_2_LC_6_8_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_2_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_2_LC_6_8_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNI_2_LC_6_8_7  (
            .in0(N__19679),
            .in1(N__19661),
            .in2(N__19640),
            .in3(N__19637),
            .lcout(\VPP_VDDQ.un9_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_6_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_6_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(N__21569),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(\POWERLED.mult1_un138_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_6_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_6_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__20420),
            .in2(N__20037),
            .in3(N__20009),
            .lcout(\POWERLED.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_6_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_6_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(N__20006),
            .in2(N__20039),
            .in3(N__19991),
            .lcout(\POWERLED.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_6_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_6_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(N__20063),
            .in2(N__19988),
            .in3(N__19973),
            .lcout(\POWERLED.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_6_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_6_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__19970),
            .in2(N__20071),
            .in3(N__19955),
            .lcout(\POWERLED.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_6_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_6_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_6_10_5  (
            .in0(N__19916),
            .in1(N__19952),
            .in2(N__20038),
            .in3(N__19940),
            .lcout(\POWERLED.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_6_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_6_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_6_10_6  (
            .in0(N__19937),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19931),
            .lcout(\POWERLED.mult1_un138_sum_s_8 ),
            .ltout(\POWERLED.mult1_un138_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_10_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19898),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_2_LC_6_11_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_1_2_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_2_LC_6_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_2_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(N__32955),
            .in2(_gnd_net_),
            .in3(N__29442),
            .lcout(\POWERLED.N_613 ),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(\POWERLED.mult1_un152_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(N__20106),
            .in2(N__20411),
            .in3(N__20171),
            .lcout(\POWERLED.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(N__20168),
            .in2(N__20111),
            .in3(N__20162),
            .lcout(\POWERLED.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(N__20133),
            .in2(N__20159),
            .in3(N__20150),
            .lcout(\POWERLED.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_11_4  (
            .in0(_gnd_net_),
            .in1(N__20147),
            .in2(N__20140),
            .in3(N__20114),
            .lcout(\POWERLED.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_11_5  (
            .in0(N__20227),
            .in1(N__20110),
            .in2(N__20096),
            .in3(N__20084),
            .lcout(\POWERLED.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_11_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_11_6  (
            .in0(N__20081),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20075),
            .lcout(\POWERLED.mult1_un152_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_6_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_6_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_6_11_7  (
            .in0(N__20067),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_6_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_6_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_6_12_0  (
            .in0(_gnd_net_),
            .in1(N__30929),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_12_0_),
            .carryout(\POWERLED.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_6_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_6_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_6_12_1  (
            .in0(_gnd_net_),
            .in1(N__20196),
            .in2(N__22592),
            .in3(N__20342),
            .lcout(\POWERLED.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_6_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_6_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(N__20339),
            .in2(N__20203),
            .in3(N__20324),
            .lcout(\POWERLED.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_6_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_6_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_6_12_3  (
            .in0(_gnd_net_),
            .in1(N__20321),
            .in2(N__20237),
            .in3(N__20309),
            .lcout(\POWERLED.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_6_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_6_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_6_12_4  (
            .in0(_gnd_net_),
            .in1(N__20306),
            .in2(N__20236),
            .in3(N__20294),
            .lcout(\POWERLED.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_6_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_6_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_6_12_5  (
            .in0(N__20257),
            .in1(N__20291),
            .in2(N__20204),
            .in3(N__20279),
            .lcout(\POWERLED.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_6_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_6_12_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_6_12_6  (
            .in0(N__20276),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20270),
            .lcout(\POWERLED.mult1_un159_sum_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20228),
            .lcout(\POWERLED.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_13_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21565),
            .lcout(\POWERLED.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_13_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21544),
            .lcout(\POWERLED.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_6_13_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_6_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_6_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21580),
            .lcout(\POWERLED.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_6_13_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_6_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_6_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21757),
            .lcout(\POWERLED.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_13_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_13_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_13_4  (
            .in0(N__21523),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_6_13_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_6_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_6_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21478),
            .lcout(\POWERLED.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_6_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_6_13_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_6_13_6  (
            .in0(N__21615),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un61_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21614),
            .lcout(\POWERLED.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(N__21829),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_14_0_),
            .carryout(\POWERLED.mult1_un68_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(N__21764),
            .in2(N__20461),
            .in3(N__20354),
            .lcout(\POWERLED.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_14_2  (
            .in0(_gnd_net_),
            .in1(N__20457),
            .in2(N__21431),
            .in3(N__20471),
            .lcout(\POWERLED.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(N__21407),
            .in2(N__21626),
            .in3(N__20468),
            .lcout(\POWERLED.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(N__21625),
            .in2(N__21389),
            .in3(N__20465),
            .lcout(\POWERLED.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_14_5  (
            .in0(N__20591),
            .in1(N__21365),
            .in2(N__20462),
            .in3(N__20444),
            .lcout(\POWERLED.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_14_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(N__21344),
            .in2(_gnd_net_),
            .in3(N__20441),
            .lcout(\POWERLED.mult1_un68_sum_s_8 ),
            .ltout(\POWERLED.mult1_un68_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20438),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(N__21688),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_15_0_),
            .carryout(\POWERLED.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_15_1  (
            .in0(_gnd_net_),
            .in1(N__21818),
            .in2(N__20554),
            .in3(N__20435),
            .lcout(\POWERLED.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_15_2  (
            .in0(_gnd_net_),
            .in1(N__20550),
            .in2(N__20432),
            .in3(N__20423),
            .lcout(\POWERLED.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_15_3  (
            .in0(_gnd_net_),
            .in1(N__20612),
            .in2(N__20599),
            .in3(N__20606),
            .lcout(\POWERLED.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_15_4  (
            .in0(_gnd_net_),
            .in1(N__20595),
            .in2(N__20573),
            .in3(N__20564),
            .lcout(\POWERLED.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_15_5  (
            .in0(N__20738),
            .in1(N__20561),
            .in2(N__20555),
            .in3(N__20537),
            .lcout(\POWERLED.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_15_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20534),
            .in3(N__20525),
            .lcout(\POWERLED.mult1_un75_sum_s_8 ),
            .ltout(\POWERLED.mult1_un75_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_15_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20522),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_16_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21806),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_16_0_),
            .carryout(\POWERLED.mult1_un82_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_16_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_16_1  (
            .in0(_gnd_net_),
            .in1(N__20627),
            .in2(N__20695),
            .in3(N__20510),
            .lcout(\POWERLED.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_16_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_16_2  (
            .in0(_gnd_net_),
            .in1(N__20691),
            .in2(N__20507),
            .in3(N__20492),
            .lcout(\POWERLED.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_16_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_16_3  (
            .in0(_gnd_net_),
            .in1(N__20489),
            .in2(N__20744),
            .in3(N__20474),
            .lcout(\POWERLED.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_16_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_16_4  (
            .in0(_gnd_net_),
            .in1(N__20742),
            .in2(N__20720),
            .in3(N__20705),
            .lcout(\POWERLED.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_16_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_16_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_16_5  (
            .in0(N__20649),
            .in1(N__20702),
            .in2(N__20696),
            .in3(N__20669),
            .lcout(\POWERLED.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_16_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_16_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20666),
            .in3(N__20657),
            .lcout(\POWERLED.mult1_un82_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_16_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21692),
            .lcout(\POWERLED.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_9_LC_7_2_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_9_LC_7_2_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_9_LC_7_2_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_9_LC_7_2_0  (
            .in0(N__20873),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32045),
            .ce(N__23546),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIN3TIG_9_LC_7_2_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIN3TIG_9_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIN3TIG_9_LC_7_2_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNIN3TIG_9_LC_7_2_1  (
            .in0(N__20621),
            .in1(N__23541),
            .in2(_gnd_net_),
            .in3(N__20872),
            .lcout(\POWERLED.count_offZ0Z_9 ),
            .ltout(\POWERLED.count_offZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_10_LC_7_2_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_10_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_10_LC_7_2_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_10_LC_7_2_2  (
            .in0(N__20794),
            .in1(N__20854),
            .in2(N__20615),
            .in3(N__20824),
            .lcout(\POWERLED.un34_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI0E2HG_10_LC_7_2_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI0E2HG_10_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI0E2HG_10_LC_7_2_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNI0E2HG_10_LC_7_2_3  (
            .in0(N__20771),
            .in1(N__20839),
            .in2(_gnd_net_),
            .in3(N__23542),
            .lcout(\POWERLED.count_offZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_10_LC_7_2_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_10_LC_7_2_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_10_LC_7_2_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_10_LC_7_2_4  (
            .in0(N__20840),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32045),
            .ce(N__23546),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI9LFFG_11_LC_7_2_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI9LFFG_11_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI9LFFG_11_LC_7_2_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNI9LFFG_11_LC_7_2_5  (
            .in0(N__20765),
            .in1(N__20809),
            .in2(_gnd_net_),
            .in3(N__23543),
            .lcout(\POWERLED.count_offZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_11_LC_7_2_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_11_LC_7_2_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_11_LC_7_2_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_11_LC_7_2_6  (
            .in0(N__20810),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32045),
            .ce(N__23546),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIBOGFG_12_LC_7_2_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIBOGFG_12_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIBOGFG_12_LC_7_2_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIBOGFG_12_LC_7_2_7  (
            .in0(N__21083),
            .in1(N__21098),
            .in2(_gnd_net_),
            .in3(N__23544),
            .lcout(\POWERLED.count_offZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_7_3_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_7_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_LC_7_3_0  (
            .in0(_gnd_net_),
            .in1(N__23396),
            .in2(N__22090),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_3_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI5IAA7_LC_7_3_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI5IAA7_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI5IAA7_LC_7_3_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_RNI5IAA7_LC_7_3_1  (
            .in0(N__26130),
            .in1(N__21919),
            .in2(_gnd_net_),
            .in3(N__20759),
            .lcout(\POWERLED.count_off_1_2 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_1_cZ0 ),
            .carryout(\POWERLED.un3_count_off_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_7_3_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_7_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_7_3_2  (
            .in0(_gnd_net_),
            .in1(N__23210),
            .in2(_gnd_net_),
            .in3(N__20756),
            .lcout(\POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_2 ),
            .carryout(\POWERLED.un3_count_off_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_7_3_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_7_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_7_3_3  (
            .in0(_gnd_net_),
            .in1(N__23606),
            .in2(_gnd_net_),
            .in3(N__20753),
            .lcout(\POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_3 ),
            .carryout(\POWERLED.un3_count_off_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI8ODA7_LC_7_3_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI8ODA7_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI8ODA7_LC_7_3_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_4_c_RNI8ODA7_LC_7_3_4  (
            .in0(N__26126),
            .in1(N__21959),
            .in2(_gnd_net_),
            .in3(N__20750),
            .lcout(\POWERLED.count_off_1_5 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_4 ),
            .carryout(\POWERLED.un3_count_off_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI9QEA7_LC_7_3_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI9QEA7_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI9QEA7_LC_7_3_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_5_c_RNI9QEA7_LC_7_3_5  (
            .in0(N__26128),
            .in1(N__22036),
            .in2(_gnd_net_),
            .in3(N__20747),
            .lcout(\POWERLED.count_off_1_6 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_5 ),
            .carryout(\POWERLED.un3_count_off_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNIASFA7_LC_7_3_6 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNIASFA7_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNIASFA7_LC_7_3_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_6_c_RNIASFA7_LC_7_3_6  (
            .in0(N__26127),
            .in1(N__23191),
            .in2(_gnd_net_),
            .in3(N__20888),
            .lcout(\POWERLED.count_off_1_7 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_6 ),
            .carryout(\POWERLED.un3_count_off_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNIBUGA7_LC_7_3_7 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNIBUGA7_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNIBUGA7_LC_7_3_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_7_c_RNIBUGA7_LC_7_3_7  (
            .in0(N__26129),
            .in1(N__23167),
            .in2(_gnd_net_),
            .in3(N__20885),
            .lcout(\POWERLED.count_off_1_8 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_7 ),
            .carryout(\POWERLED.un3_count_off_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNIC0IA7_LC_7_4_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNIC0IA7_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNIC0IA7_LC_7_4_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_8_c_RNIC0IA7_LC_7_4_0  (
            .in0(N__26119),
            .in1(N__20882),
            .in2(_gnd_net_),
            .in3(N__20861),
            .lcout(\POWERLED.count_off_1_9 ),
            .ltout(),
            .carryin(bfn_7_4_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNID2JA7_LC_7_4_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNID2JA7_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNID2JA7_LC_7_4_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_9_c_RNID2JA7_LC_7_4_1  (
            .in0(N__26122),
            .in1(_gnd_net_),
            .in2(N__20858),
            .in3(N__20828),
            .lcout(\POWERLED.count_off_1_10 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_9 ),
            .carryout(\POWERLED.un3_count_off_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIL8097_LC_7_4_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIL8097_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIL8097_LC_7_4_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_10_c_RNIL8097_LC_7_4_2  (
            .in0(N__26120),
            .in1(N__20825),
            .in2(_gnd_net_),
            .in3(N__20798),
            .lcout(\POWERLED.count_off_1_11 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_10 ),
            .carryout(\POWERLED.un3_count_off_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIMA197_LC_7_4_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIMA197_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIMA197_LC_7_4_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_11_c_RNIMA197_LC_7_4_3  (
            .in0(N__26123),
            .in1(N__20795),
            .in2(_gnd_net_),
            .in3(N__20780),
            .lcout(\POWERLED.count_off_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_11 ),
            .carryout(\POWERLED.un3_count_off_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNINC297_LC_7_4_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNINC297_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNINC297_LC_7_4_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_12_c_RNINC297_LC_7_4_4  (
            .in0(N__26121),
            .in1(N__22117),
            .in2(_gnd_net_),
            .in3(N__20777),
            .lcout(\POWERLED.count_off_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_12 ),
            .carryout(\POWERLED.un3_count_off_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIOE397_LC_7_4_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIOE397_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIOE397_LC_7_4_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_13_c_RNIOE397_LC_7_4_5  (
            .in0(N__26124),
            .in1(N__22105),
            .in2(_gnd_net_),
            .in3(N__20774),
            .lcout(\POWERLED.count_off_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_13 ),
            .carryout(\POWERLED.un3_count_off_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIPG497_LC_7_4_6 .C_ON=1'b0;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIPG497_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIPG497_LC_7_4_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_14_c_RNIPG497_LC_7_4_6  (
            .in0(N__22124),
            .in1(N__26125),
            .in2(_gnd_net_),
            .in3(N__21101),
            .lcout(\POWERLED.un3_count_off_1_cry_14_c_RNIPGZ0Z497 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_12_LC_7_4_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_12_LC_7_4_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_12_LC_7_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_12_LC_7_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21097),
            .lcout(\POWERLED.count_off_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32046),
            .ce(N__23537),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_LC_7_5_0 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_LC_7_5_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_LC_7_5_0 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \COUNTER.tmp_0_LC_7_5_0  (
            .in0(N__25620),
            .in1(_gnd_net_),
            .in2(N__22524),
            .in3(_gnd_net_),
            .lcout(clk_100Khz_signalkeep_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32349),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_en_LC_7_5_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_en_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_en_LC_7_5_1 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \POWERLED.func_state_en_LC_7_5_1  (
            .in0(N__29557),
            .in1(N__25619),
            .in2(N__30739),
            .in3(N__22504),
            .lcout(\POWERLED.func_state_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_RNO_LC_7_5_2 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_7_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_4_c_RNO_LC_7_5_2  (
            .in0(N__21073),
            .in1(N__21061),
            .in2(N__21050),
            .in3(N__21034),
            .lcout(\COUNTER.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_RNO_LC_7_5_3 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_7_5_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_5_c_RNO_LC_7_5_3  (
            .in0(N__21022),
            .in1(N__21010),
            .in2(N__20999),
            .in3(N__20983),
            .lcout(\COUNTER.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_14_LC_7_6_0 .C_ON=1'b0;
    defparam \POWERLED.G_14_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_14_LC_7_6_0 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \POWERLED.G_14_LC_7_6_0  (
            .in0(N__21213),
            .in1(N__20910),
            .in2(N__20972),
            .in3(N__25399),
            .lcout(G_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_1_LC_7_6_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_1_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_1_LC_7_6_3 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \RSMRST_PWRGD.curr_state_1_LC_7_6_3  (
            .in0(N__26824),
            .in1(N__21216),
            .in2(N__20917),
            .in3(N__21152),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32179),
            .ce(N__25311),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_7_6_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_7_6_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_fast_LC_7_6_4  (
            .in0(N__21148),
            .in1(N__26821),
            .in2(_gnd_net_),
            .in3(N__21217),
            .lcout(RSMRSTn_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32179),
            .ce(N__25311),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_7_6_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_7_6_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_7_6_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_7_6_5  (
            .in0(N__26822),
            .in1(N__21215),
            .in2(_gnd_net_),
            .in3(N__21151),
            .lcout(RSMRSTn_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32179),
            .ce(N__25311),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep2_LC_7_6_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep2_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep2_LC_7_6_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_rep2_LC_7_6_6  (
            .in0(N__21149),
            .in1(N__26823),
            .in2(_gnd_net_),
            .in3(N__21218),
            .lcout(RSMRSTn_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32179),
            .ce(N__25311),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_7_6_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_7_6_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_LC_7_6_7  (
            .in0(N__26820),
            .in1(N__21214),
            .in2(_gnd_net_),
            .in3(N__21150),
            .lcout(rsmrstn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32179),
            .ce(N__25311),
            .sr(_gnd_net_));
    defparam \POWERLED.N_430_i_LC_7_7_0 .C_ON=1'b0;
    defparam \POWERLED.N_430_i_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.N_430_i_LC_7_7_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.N_430_i_LC_7_7_0  (
            .in0(N__26747),
            .in1(N__26367),
            .in2(N__27617),
            .in3(N__25658),
            .lcout(\POWERLED.N_430_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.VCCST_EN_i_0_o2_LC_7_7_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.VCCST_EN_i_0_o2_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.VCCST_EN_i_0_o2_LC_7_7_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \PCH_PWRGD.VCCST_EN_i_0_o2_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__30575),
            .in2(_gnd_net_),
            .in3(N__29844),
            .lcout(VCCST_EN_i_1),
            .ltout(VCCST_EN_i_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_LC_7_7_3 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_LC_7_7_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_LC_7_7_3  (
            .in0(N__21113),
            .in1(N__28813),
            .in2(N__21119),
            .in3(N__28590),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_o_N_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_LC_7_7_4 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_LC_7_7_4 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_LC_7_7_4  (
            .in0(N__21107),
            .in1(N__25988),
            .in2(N__21116),
            .in3(N__23738),
            .lcout(\POWERLED.un1_func_state25_6_0_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_0_o2_LC_7_7_5 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_0_o2_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_0_o2_LC_7_7_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \POWERLED.un1_func_state25_6_0_0_o2_LC_7_7_5  (
            .in0(N__30420),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26748),
            .lcout(\POWERLED.N_432 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_3_2_LC_7_7_6 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_3_2_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_3_2_LC_7_7_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_3_2_LC_7_7_6  (
            .in0(N__27575),
            .in1(N__30577),
            .in2(N__26756),
            .in3(N__30421),
            .lcout(\POWERLED.un1_func_state25_6_0_o_N_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBVNS_0_LC_7_7_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_0_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_0_LC_7_7_7 .LUT_INIT=16'b0100100000000000;
    LogicCell40 \POWERLED.func_state_RNIBVNS_0_LC_7_7_7  (
            .in0(N__30576),
            .in1(N__27574),
            .in2(N__30422),
            .in3(N__26235),
            .lcout(\POWERLED.func_state_RNIBVNSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI78D82_1_LC_7_8_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI78D82_1_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI78D82_1_LC_7_8_0 .LUT_INIT=16'b0100000001110000;
    LogicCell40 \POWERLED.func_state_RNI78D82_1_LC_7_8_0  (
            .in0(N__22426),
            .in1(N__21257),
            .in2(N__30074),
            .in3(N__25655),
            .lcout(),
            .ltout(\POWERLED.func_state_1_ss0_i_0_0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3H2K3_1_LC_7_8_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3H2K3_1_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3H2K3_1_LC_7_8_1 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \POWERLED.func_state_RNI3H2K3_1_LC_7_8_1  (
            .in0(N__28814),
            .in1(N__21251),
            .in2(N__21260),
            .in3(N__25874),
            .lcout(\POWERLED.N_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.N_215_i_0_o2_0_LC_7_8_2 .C_ON=1'b0;
    defparam \POWERLED.N_215_i_0_o2_0_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.N_215_i_0_o2_0_LC_7_8_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \POWERLED.N_215_i_0_o2_0_LC_7_8_2  (
            .in0(N__30388),
            .in1(N__30722),
            .in2(N__27663),
            .in3(N__26752),
            .lcout(\POWERLED.N_423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIMJ6IF_1_LC_7_8_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIMJ6IF_1_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIMJ6IF_1_LC_7_8_3 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \POWERLED.func_state_RNIMJ6IF_1_LC_7_8_3  (
            .in0(N__21241),
            .in1(N__33067),
            .in2(N__21230),
            .in3(N__22396),
            .lcout(func_state_RNIMJ6IF_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBVNS_1_0_LC_7_8_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_1_0_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_1_0_LC_7_8_4 .LUT_INIT=16'b0110000000000000;
    LogicCell40 \POWERLED.func_state_RNIBVNS_1_0_LC_7_8_4  (
            .in0(N__30389),
            .in1(N__30723),
            .in2(N__27664),
            .in3(N__28815),
            .lcout(\POWERLED.N_673 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIP4521_0_1_LC_7_8_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIP4521_0_1_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIP4521_0_1_LC_7_8_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \POWERLED.func_state_RNIP4521_0_1_LC_7_8_5  (
            .in0(N__25656),
            .in1(N__27640),
            .in2(N__26383),
            .in3(N__30022),
            .lcout(\POWERLED.N_542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_0_a2_5_LC_7_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_0_a2_5_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_0_a2_5_LC_7_8_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_0_a2_5_LC_7_8_6  (
            .in0(N__26753),
            .in1(N__25657),
            .in2(N__27665),
            .in3(N__26371),
            .lcout(\POWERLED.N_671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_LC_7_8_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_1_LC_7_8_7 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \POWERLED.func_state_1_LC_7_8_7  (
            .in0(N__21229),
            .in1(N__33068),
            .in2(N__21245),
            .in3(N__22397),
            .lcout(\POWERLED.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32205),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6SKJ1_11_LC_7_9_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6SKJ1_11_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6SKJ1_11_LC_7_9_0 .LUT_INIT=16'b1000000011001100;
    LogicCell40 \POWERLED.dutycycle_RNI6SKJ1_11_LC_7_9_0  (
            .in0(N__29862),
            .in1(N__30266),
            .in2(N__29742),
            .in3(N__24703),
            .lcout(),
            .ltout(\POWERLED.N_512_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5TUF2_11_LC_7_9_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5TUF2_11_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5TUF2_11_LC_7_9_1 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \POWERLED.dutycycle_RNI5TUF2_11_LC_7_9_1  (
            .in0(N__24704),
            .in1(N__27452),
            .in2(N__21302),
            .in3(N__30014),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_39_and_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIRUFD6_11_LC_7_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIRUFD6_11_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIRUFD6_11_LC_7_9_2 .LUT_INIT=16'b0010001000101010;
    LogicCell40 \POWERLED.dutycycle_RNIRUFD6_11_LC_7_9_2  (
            .in0(N__32629),
            .in1(N__32812),
            .in2(N__21299),
            .in3(N__21296),
            .lcout(\POWERLED.dutycycle_en_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI24KO1_10_LC_7_9_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI24KO1_10_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI24KO1_10_LC_7_9_3 .LUT_INIT=16'b0000100010101010;
    LogicCell40 \POWERLED.dutycycle_RNI24KO1_10_LC_7_9_3  (
            .in0(N__27878),
            .in1(N__33086),
            .in2(N__24815),
            .in3(N__27834),
            .lcout(\POWERLED.N_508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI24KO1_11_LC_7_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI24KO1_11_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI24KO1_11_LC_7_9_5 .LUT_INIT=16'b0100000011110000;
    LogicCell40 \POWERLED.dutycycle_RNI24KO1_11_LC_7_9_5  (
            .in0(N__24702),
            .in1(N__33085),
            .in2(N__27892),
            .in3(N__27833),
            .lcout(\POWERLED.N_514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5TUF2_10_LC_7_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5TUF2_10_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5TUF2_10_LC_7_9_6 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \POWERLED.dutycycle_RNI5TUF2_10_LC_7_9_6  (
            .in0(N__24813),
            .in1(N__30073),
            .in2(N__27461),
            .in3(N__23801),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_33_and_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIRUFD6_10_LC_7_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIRUFD6_10_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIRUFD6_10_LC_7_9_7 .LUT_INIT=16'b0000010011001100;
    LogicCell40 \POWERLED.dutycycle_RNIRUFD6_10_LC_7_9_7  (
            .in0(N__21290),
            .in1(N__32630),
            .in2(N__21284),
            .in3(N__32813),
            .lcout(\POWERLED.dutycycle_en_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIJTQIG_7_LC_7_10_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIJTQIG_7_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIJTQIG_7_LC_7_10_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNIJTQIG_7_LC_7_10_0  (
            .in0(N__21266),
            .in1(N__23520),
            .in2(_gnd_net_),
            .in3(N__21280),
            .lcout(\POWERLED.count_offZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_7_LC_7_10_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_7_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_7_LC_7_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_7_LC_7_10_1  (
            .in0(N__21281),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32322),
            .ce(N__23538),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIL0SIG_8_LC_7_10_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIL0SIG_8_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIL0SIG_8_LC_7_10_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNIL0SIG_8_LC_7_10_2  (
            .in0(N__21320),
            .in1(N__23521),
            .in2(_gnd_net_),
            .in3(N__21331),
            .lcout(\POWERLED.count_offZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_8_LC_7_10_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_8_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_8_LC_7_10_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_8_LC_7_10_3  (
            .in0(N__21332),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32322),
            .ce(N__23538),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_10_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_10_4 .LUT_INIT=16'b1111101000000101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_10_4  (
            .in0(N__22812),
            .in1(_gnd_net_),
            .in2(N__22790),
            .in3(N__21853),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_10_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_10_5 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(N__22813),
            .in2(N__21857),
            .in3(N__22789),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22811),
            .lcout(\POWERLED.un1_dutycycle_53_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__21658),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\POWERLED.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_11_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21596),
            .in3(N__21314),
            .lcout(\POWERLED.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__22871),
            .in2(N__22853),
            .in3(N__21311),
            .lcout(\POWERLED.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__25182),
            .in2(N__22709),
            .in3(N__21308),
            .lcout(\POWERLED.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__25194),
            .in2(N__22688),
            .in3(N__21305),
            .lcout(\POWERLED.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_7_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_7_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_7_11_5  (
            .in0(N__22632),
            .in1(N__22667),
            .in2(N__21455),
            .in3(N__21461),
            .lcout(\POWERLED.mult1_un61_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_11_6 .C_ON=1'b0;
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21458),
            .lcout(\POWERLED.mult1_un54_sum_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_7_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_7_11_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_7_11_7  (
            .in0(N__22665),
            .in1(N__22666),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__21779),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\POWERLED.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__21446),
            .in2(N__22615),
            .in3(N__21419),
            .lcout(\POWERLED.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_7_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_7_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__22611),
            .in2(N__21416),
            .in3(N__21398),
            .lcout(\POWERLED.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_7_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_7_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(N__21395),
            .in2(N__22637),
            .in3(N__21377),
            .lcout(\POWERLED.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_7_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_7_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__22636),
            .in2(N__21374),
            .in3(N__21353),
            .lcout(\POWERLED.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_7_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_7_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_7_12_5  (
            .in0(N__21616),
            .in1(N__21350),
            .in2(N__22616),
            .in3(N__21335),
            .lcout(\POWERLED.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_7_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_7_12_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_7_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21638),
            .in3(N__21629),
            .lcout(\POWERLED.mult1_un61_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_12_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22744),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_dutycycle_53_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_0_LC_7_13_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_1_0_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_0_LC_7_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \POWERLED.dutycycle_RNI_1_0_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__26548),
            .in2(N__31028),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_dutycycle_53_axb_0 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__22844),
            .in2(N__26557),
            .in3(N__21554),
            .lcout(\POWERLED.mult1_un138_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__32949),
            .in2(N__22826),
            .in3(N__21533),
            .lcout(\POWERLED.mult1_un131_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_1 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__32858),
            .in2(N__32957),
            .in3(N__21512),
            .lcout(\POWERLED.mult1_un124_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_2 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__31169),
            .in2(N__31186),
            .in3(N__21485),
            .lcout(\POWERLED.mult1_un117_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_3 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__31321),
            .in2(N__22835),
            .in3(N__21464),
            .lcout(\POWERLED.mult1_un110_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_4 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_13_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__31314),
            .in2(N__22976),
            .in3(N__21743),
            .lcout(\POWERLED.mult1_un103_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_5 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_13_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__22988),
            .in2(N__24809),
            .in3(N__21719),
            .lcout(\POWERLED.mult1_un96_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_6 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__24701),
            .in2(N__24203),
            .in3(N__21698),
            .lcout(\POWERLED.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__26973),
            .in2(N__22952),
            .in3(N__21695),
            .lcout(\POWERLED.mult1_un82_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_8 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__24093),
            .in2(N__22898),
            .in3(N__21677),
            .lcout(\POWERLED.mult1_un75_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__27747),
            .in2(N__24254),
            .in3(N__21674),
            .lcout(\POWERLED.mult1_un68_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__27506),
            .in2(N__23063),
            .in3(N__21671),
            .lcout(\POWERLED.mult1_un61_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__24094),
            .in2(N__24278),
            .in3(N__21644),
            .lcout(\POWERLED.mult1_un54_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_14_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__23030),
            .in2(N__27763),
            .in3(N__21641),
            .lcout(\POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_14_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(N__21812),
            .in2(N__27519),
            .in3(N__21866),
            .lcout(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_14 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__27510),
            .in2(N__21839),
            .in3(N__21863),
            .lcout(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\POWERLED.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_15_1 .C_ON=1'b0;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.CO2_THRU_LUT4_0_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21860),
            .lcout(\POWERLED.CO2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_14_LC_7_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_14_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_14_LC_7_15_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_14_LC_7_15_2  (
            .in0(N__27746),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23096),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_7_15_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_7_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21830),
            .lcout(\POWERLED.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_15_LC_7_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_15_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_15_LC_7_15_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_15_LC_7_15_4  (
            .in0(N__27745),
            .in1(N__27511),
            .in2(_gnd_net_),
            .in3(N__23095),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_15_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21802),
            .lcout(\POWERLED.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI12AS_8_LC_7_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI12AS_8_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI12AS_8_LC_7_15_6 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \POWERLED.dutycycle_RNI12AS_8_LC_7_15_6  (
            .in0(N__30602),
            .in1(N__24441),
            .in2(_gnd_net_),
            .in3(N__29894),
            .lcout(\POWERLED.N_599 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_7_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_7_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21778),
            .lcout(\POWERLED.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI99TE_13_LC_7_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI99TE_13_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI99TE_13_LC_7_16_0 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \POWERLED.dutycycle_RNI99TE_13_LC_7_16_0  (
            .in0(N__21878),
            .in1(N__30550),
            .in2(_gnd_net_),
            .in3(N__27677),
            .lcout(),
            .ltout(\POWERLED.N_598_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIAB7B1_13_LC_7_16_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIAB7B1_13_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIAB7B1_13_LC_7_16_1 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \POWERLED.dutycycle_RNIAB7B1_13_LC_7_16_1  (
            .in0(N__27236),
            .in1(N__24115),
            .in2(N__21893),
            .in3(N__27836),
            .lcout(),
            .ltout(\POWERLED.N_450_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI35P35_13_LC_7_16_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI35P35_13_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI35P35_13_LC_7_16_2 .LUT_INIT=16'b0111001100000000;
    LogicCell40 \POWERLED.dutycycle_RNI35P35_13_LC_7_16_2  (
            .in0(N__22352),
            .in1(N__32843),
            .in2(N__21890),
            .in3(N__32673),
            .lcout(\POWERLED.dutycycle_en_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI24KO1_8_LC_7_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI24KO1_8_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI24KO1_8_LC_7_16_3 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \POWERLED.dutycycle_RNI24KO1_8_LC_7_16_3  (
            .in0(N__27235),
            .in1(N__21887),
            .in2(N__24623),
            .in3(N__27835),
            .lcout(),
            .ltout(\POWERLED.N_449_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIRT5H5_8_LC_7_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIRT5H5_8_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIRT5H5_8_LC_7_16_4 .LUT_INIT=16'b0111001100000000;
    LogicCell40 \POWERLED.dutycycle_RNIRT5H5_8_LC_7_16_4  (
            .in0(N__22351),
            .in1(N__32842),
            .in2(N__21881),
            .in3(N__32672),
            .lcout(\POWERLED.dutycycle_RNIRT5H5Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_13_LC_7_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_7_16_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.dutycycle_RNI_1_13_LC_7_16_6  (
            .in0(N__24114),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_2376_i ),
            .ltout(\POWERLED.N_2376_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_12_LC_7_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_12_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_12_LC_7_16_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_12_LC_7_16_7  (
            .in0(N__24443),
            .in1(N__24875),
            .in2(N__21872),
            .in3(N__23036),
            .lcout(\POWERLED.N_612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIG4L3G_0_LC_8_2_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIG4L3G_0_LC_8_2_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIG4L3G_0_LC_8_2_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIG4L3G_0_LC_8_2_0  (
            .in0(N__21950),
            .in1(N__21944),
            .in2(_gnd_net_),
            .in3(N__23483),
            .lcout(\POWERLED.count_offZ0Z_0 ),
            .ltout(\POWERLED.count_offZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_1_LC_8_2_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_1_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_1_LC_8_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.count_off_RNI_1_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21869),
            .in3(N__23392),
            .lcout(\POWERLED.count_off_RNIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIFNOIG_5_LC_8_2_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIFNOIG_5_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIFNOIG_5_LC_8_2_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIFNOIG_5_LC_8_2_2  (
            .in0(N__21989),
            .in1(N__21970),
            .in2(_gnd_net_),
            .in3(N__23485),
            .lcout(\POWERLED.count_offZ0Z_5 ),
            .ltout(\POWERLED.count_offZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_0_1_LC_8_2_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_0_1_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_0_1_LC_8_2_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.count_off_RNI_0_1_LC_8_2_3  (
            .in0(N__21920),
            .in1(N__22037),
            .in2(N__21953),
            .in3(N__23391),
            .lcout(\POWERLED.un34_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_0_LC_8_2_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_0_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_0_LC_8_2_4 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \POWERLED.count_off_0_LC_8_2_4  (
            .in0(N__26132),
            .in1(_gnd_net_),
            .in2(N__22091),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32265),
            .ce(N__23518),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIEAAR6_0_LC_8_2_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIEAAR6_0_LC_8_2_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIEAAR6_0_LC_8_2_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.count_off_RNIEAAR6_0_LC_8_2_5  (
            .in0(_gnd_net_),
            .in1(N__22085),
            .in2(_gnd_net_),
            .in3(N__26131),
            .lcout(\POWERLED.count_off_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_2_LC_8_2_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_2_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_2_LC_8_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_2_LC_8_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21928),
            .lcout(\POWERLED.count_off_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32265),
            .ce(N__23518),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI9ELIG_2_LC_8_2_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI9ELIG_2_LC_8_2_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI9ELIG_2_LC_8_2_7 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \POWERLED.count_off_RNI9ELIG_2_LC_8_2_7  (
            .in0(N__23484),
            .in1(N__21938),
            .in2(N__21932),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_offZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_15_LC_8_3_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_15_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_15_LC_8_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_15_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22138),
            .lcout(\POWERLED.count_off_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32279),
            .ce(N__23489),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIDRHFG_13_LC_8_3_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIDRHFG_13_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIDRHFG_13_LC_8_3_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIDRHFG_13_LC_8_3_1  (
            .in0(N__21899),
            .in1(N__21907),
            .in2(_gnd_net_),
            .in3(N__23487),
            .lcout(\POWERLED.count_offZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_13_LC_8_3_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_13_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_13_LC_8_3_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_13_LC_8_3_2  (
            .in0(N__21908),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32279),
            .ce(N__23489),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIFUIFG_14_LC_8_3_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIFUIFG_14_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIFUIFG_14_LC_8_3_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIFUIFG_14_LC_8_3_3  (
            .in0(N__22145),
            .in1(N__22153),
            .in2(_gnd_net_),
            .in3(N__23488),
            .lcout(\POWERLED.count_offZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_14_LC_8_3_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_14_LC_8_3_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_14_LC_8_3_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_14_LC_8_3_4  (
            .in0(N__22154),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32279),
            .ce(N__23489),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIH1KFG_15_LC_8_3_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIH1KFG_15_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIH1KFG_15_LC_8_3_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_off_RNIH1KFG_15_LC_8_3_5  (
            .in0(N__22139),
            .in1(N__22130),
            .in2(_gnd_net_),
            .in3(N__23490),
            .lcout(\POWERLED.count_offZ0Z_15 ),
            .ltout(\POWERLED.count_offZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_15_LC_8_3_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_15_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_15_LC_8_3_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_15_LC_8_3_6  (
            .in0(N__22118),
            .in1(N__22106),
            .in2(N__22094),
            .in3(N__22089),
            .lcout(\POWERLED.un34_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIHQPIG_6_LC_8_3_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIHQPIG_6_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIHQPIG_6_LC_8_3_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNIHQPIG_6_LC_8_3_7  (
            .in0(N__22064),
            .in1(N__23486),
            .in2(_gnd_net_),
            .in3(N__22048),
            .lcout(\POWERLED.count_offZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_LC_8_4_0 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_0_c_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_LC_8_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_LC_8_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22025),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(\COUNTER.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_LC_8_4_1 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_1_c_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_LC_8_4_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_1_c_LC_8_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22013),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_0 ),
            .carryout(\COUNTER.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_LC_8_4_2 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_2_c_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_LC_8_4_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_2_c_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22001),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_1 ),
            .carryout(\COUNTER.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_LC_8_4_3 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_3_c_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_LC_8_4_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_3_c_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22229),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_2 ),
            .carryout(\COUNTER.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_LC_8_4_4 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_4_c_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_LC_8_4_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_4_c_LC_8_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22214),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_3 ),
            .carryout(\COUNTER.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_LC_8_4_5 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_5_c_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_LC_8_4_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_5_c_LC_8_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22205),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_4 ),
            .carryout(\COUNTER.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_LC_8_4_6 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_6_c_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_LC_8_4_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_6_c_LC_8_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22196),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_5 ),
            .carryout(\COUNTER.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_LC_8_4_7 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_7_c_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_LC_8_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_7_c_LC_8_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22181),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_6 ),
            .carryout(COUNTER_un4_counter_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_8_5_0.C_ON=1'b0;
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_8_5_0.SEQ_MODE=4'b0000;
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_8_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 COUNTER_un4_counter_7_THRU_LUT4_0_LC_8_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22166),
            .lcout(COUNTER_un4_counter_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOGRS_0_0_LC_8_5_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOGRS_0_0_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOGRS_0_0_LC_8_5_2 .LUT_INIT=16'b0110000000000000;
    LogicCell40 \POWERLED.func_state_RNIOGRS_0_0_LC_8_5_2  (
            .in0(N__30736),
            .in1(N__30414),
            .in2(N__22252),
            .in3(N__28847),
            .lcout(),
            .ltout(\POWERLED.N_673_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIE48E2_1_LC_8_5_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIE48E2_1_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIE48E2_1_LC_8_5_3 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \POWERLED.func_state_RNIE48E2_1_LC_8_5_3  (
            .in0(N__22160),
            .in1(N__23657),
            .in2(N__22163),
            .in3(N__30075),
            .lcout(\POWERLED.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.g0_11_LC_8_5_4 .C_ON=1'b0;
    defparam \POWERLED.g0_11_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.g0_11_LC_8_5_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \POWERLED.g0_11_LC_8_5_4  (
            .in0(N__30737),
            .in1(N__30415),
            .in2(N__22253),
            .in3(N__26745),
            .lcout(\POWERLED.N_423_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_fast_LC_8_5_5 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_fast_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_fast_LC_8_5_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.tmp_0_fast_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(N__23656),
            .in2(_gnd_net_),
            .in3(N__22521),
            .lcout(clk_100Khz_signalkeep_3_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32281),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_0_LC_8_5_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_0_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_0_LC_8_5_6 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_0_LC_8_5_6  (
            .in0(N__30738),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30416),
            .lcout(N_247),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_LC_8_6_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_0_LC_8_6_0 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \POWERLED.func_state_0_LC_8_6_0  (
            .in0(N__23678),
            .in1(N__22271),
            .in2(N__33084),
            .in3(N__22265),
            .lcout(\POWERLED.func_stateZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32384),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_2_1_LC_8_6_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_2_1_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_2_1_LC_8_6_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.func_state_RNI_2_1_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__28832),
            .in2(_gnd_net_),
            .in3(N__30049),
            .lcout(\POWERLED.N_633 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_5_LC_8_6_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_5_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_5_LC_8_6_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_5_LC_8_6_2  (
            .in0(N__31309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29231),
            .lcout(\POWERLED.un1_dutycycle_164_0_a3_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.slp_s3n_signal_i_0_o2_2_LC_8_6_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.slp_s3n_signal_i_0_o2_2_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.slp_s3n_signal_i_0_o2_2_LC_8_6_3 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \PCH_PWRGD.slp_s3n_signal_i_0_o2_2_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27151),
            .in3(N__30412),
            .lcout(v5s_enn),
            .ltout(v5s_enn_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.g0_19_LC_8_6_4 .C_ON=1'b0;
    defparam \POWERLED.g0_19_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.g0_19_LC_8_6_4 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \POWERLED.g0_19_LC_8_6_4  (
            .in0(N__30727),
            .in1(N__25578),
            .in2(N__22274),
            .in3(N__22503),
            .lcout(\POWERLED.func_state_en_0_0 ),
            .ltout(\POWERLED.func_state_en_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI6BR4J_0_LC_8_6_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI6BR4J_0_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI6BR4J_0_LC_8_6_5 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \POWERLED.func_state_RNI6BR4J_0_LC_8_6_5  (
            .in0(N__22264),
            .in1(N__33063),
            .in2(N__22256),
            .in3(N__23677),
            .lcout(\POWERLED.func_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_m1_e_0_LC_8_6_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_m1_e_0_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_m1_e_0_LC_8_6_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \POWERLED.dutycycle_m1_e_0_LC_8_6_6  (
            .in0(N__30413),
            .in1(_gnd_net_),
            .in2(N__22251),
            .in3(N__30735),
            .lcout(\POWERLED.dutycycle_N_3_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_rep1_LC_8_6_7 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_rep1_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_rep1_LC_8_6_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \COUNTER.tmp_0_rep1_LC_8_6_7  (
            .in0(N__25579),
            .in1(N__22522),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(clk_100Khz_signalkeep_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32384),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIU8AB2_0_LC_8_7_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIU8AB2_0_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIU8AB2_0_LC_8_7_0 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \POWERLED.func_state_RNIU8AB2_0_LC_8_7_0  (
            .in0(N__22388),
            .in1(N__32768),
            .in2(N__25873),
            .in3(N__26280),
            .lcout(\POWERLED.func_state_1_m0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI7LSV8_0_LC_8_7_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI7LSV8_0_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI7LSV8_0_LC_8_7_1 .LUT_INIT=16'b1111000001000000;
    LogicCell40 \POWERLED.func_state_RNI7LSV8_0_LC_8_7_1  (
            .in0(N__31590),
            .in1(N__26240),
            .in2(N__32667),
            .in3(N__22358),
            .lcout(\POWERLED.func_state_RNI7LSV8Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5SKJ1_1_LC_8_7_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5SKJ1_1_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5SKJ1_1_LC_8_7_2 .LUT_INIT=16'b1111111100110010;
    LogicCell40 \POWERLED.func_state_RNI5SKJ1_1_LC_8_7_2  (
            .in0(N__29654),
            .in1(N__29558),
            .in2(N__29743),
            .in3(N__28925),
            .lcout(\POWERLED.func_state_RNI5SKJ1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_1_LC_8_7_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_1_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_1_LC_8_7_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.func_state_RNI_1_1_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__25864),
            .in2(_gnd_net_),
            .in3(N__29980),
            .lcout(\POWERLED.N_617 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_0_LC_8_7_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_0_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_0_LC_8_7_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_0_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__22332),
            .in2(_gnd_net_),
            .in3(N__33077),
            .lcout(N_626),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_0_LC_8_7_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_0_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_0_LC_8_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_1_0_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26425),
            .lcout(func_state_RNI_2_0),
            .ltout(func_state_RNI_2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_LC_8_7_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_LC_8_7_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \POWERLED.func_state_RNI_1_LC_8_7_6  (
            .in0(N__29981),
            .in1(_gnd_net_),
            .in2(N__22283),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_435 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.N_215_i_0_o2_LC_8_7_7 .C_ON=1'b0;
    defparam \POWERLED.N_215_i_0_o2_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.N_215_i_0_o2_LC_8_7_7 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \POWERLED.N_215_i_0_o2_LC_8_7_7  (
            .in0(N__26746),
            .in1(N__26366),
            .in2(N__27582),
            .in3(N__25577),
            .lcout(\POWERLED.N_430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIQHVM3_0_LC_8_8_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIQHVM3_0_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIQHVM3_0_LC_8_8_0 .LUT_INIT=16'b0000000011110011;
    LogicCell40 \POWERLED.func_state_RNIQHVM3_0_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__22442),
            .in2(N__26015),
            .in3(N__22280),
            .lcout(\POWERLED.func_state_1_m2_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_1_LC_8_8_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_1_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_1_LC_8_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.func_state_RNI5DLR_1_LC_8_8_1  (
            .in0(N__30705),
            .in1(N__28791),
            .in2(N__30409),
            .in3(N__30012),
            .lcout(\POWERLED.dutycycle_1_0_iv_i_0_a2_0_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_LC_8_8_2 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_LC_8_8_2 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_LC_8_8_2  (
            .in0(N__27625),
            .in1(N__30708),
            .in2(_gnd_net_),
            .in3(N__30387),
            .lcout(\POWERLED.N_443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBVNS_0_0_LC_8_8_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_0_0_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_0_0_LC_8_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.func_state_RNIBVNS_0_0_LC_8_8_3  (
            .in0(N__30706),
            .in1(N__28790),
            .in2(N__30410),
            .in3(N__27624),
            .lcout(\POWERLED.N_540_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIP4521_1_LC_8_8_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIP4521_1_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIP4521_1_LC_8_8_4 .LUT_INIT=16'b1101110011111111;
    LogicCell40 \POWERLED.func_state_RNIP4521_1_LC_8_8_4  (
            .in0(N__30013),
            .in1(N__22436),
            .in2(N__23831),
            .in3(N__29267),
            .lcout(),
            .ltout(\POWERLED.func_state_1_m2s2_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNINDFD3_1_LC_8_8_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNINDFD3_1_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNINDFD3_1_LC_8_8_5 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \POWERLED.func_state_RNINDFD3_1_LC_8_8_5  (
            .in0(N__32744),
            .in1(N__22430),
            .in2(N__22415),
            .in3(N__26276),
            .lcout(\POWERLED.N_74 ),
            .ltout(\POWERLED.N_74_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI4TUGC_1_LC_8_8_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI4TUGC_1_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI4TUGC_1_LC_8_8_6 .LUT_INIT=16'b1110000011101111;
    LogicCell40 \POWERLED.func_state_RNI4TUGC_1_LC_8_8_6  (
            .in0(N__22373),
            .in1(N__22412),
            .in2(N__22406),
            .in3(N__22403),
            .lcout(\POWERLED.func_state_1_m2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIGCDO1_0_LC_8_8_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIGCDO1_0_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIGCDO1_0_LC_8_8_7 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \POWERLED.func_state_RNIGCDO1_0_LC_8_8_7  (
            .in0(N__30707),
            .in1(N__22387),
            .in2(N__30411),
            .in3(N__26275),
            .lcout(\POWERLED.N_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIFBNT_LC_8_9_0 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIFBNT_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIFBNT_LC_8_9_0 .LUT_INIT=16'b1010111110101010;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNIFBNT_LC_8_9_0  (
            .in0(N__26029),
            .in1(_gnd_net_),
            .in2(N__23885),
            .in3(N__27861),
            .lcout(),
            .ltout(\POWERLED.dutycycle_1_0_iv_i_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIS27B2_LC_8_9_1 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIS27B2_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIS27B2_LC_8_9_1 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNIS27B2_LC_8_9_1  (
            .in0(N__26742),
            .in1(N__22367),
            .in2(N__22361),
            .in3(N__25582),
            .lcout(\POWERLED.N_71 ),
            .ltout(\POWERLED.N_71_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIVSVI5_2_LC_8_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIVSVI5_2_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIVSVI5_2_LC_8_9_2 .LUT_INIT=16'b0100111011001100;
    LogicCell40 \POWERLED.dutycycle_RNIVSVI5_2_LC_8_9_2  (
            .in0(N__22574),
            .in1(N__22558),
            .in2(N__22598),
            .in3(N__32626),
            .lcout(\POWERLED.dutycycleZ0Z_0 ),
            .ltout(\POWERLED.dutycycleZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_9_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_9_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22595),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_2_LC_8_9_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_2_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_2_LC_8_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_3_2_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__32913),
            .in2(_gnd_net_),
            .in3(N__30018),
            .lcout(),
            .ltout(\POWERLED.N_426_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIIASA2_2_LC_8_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIIASA2_2_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIIASA2_2_LC_8_9_5 .LUT_INIT=16'b0011001110111111;
    LogicCell40 \POWERLED.dutycycle_RNIIASA2_2_LC_8_9_5  (
            .in0(N__29572),
            .in1(N__32783),
            .in2(N__22577),
            .in3(N__29489),
            .lcout(\POWERLED.dutycycle_eena_1 ),
            .ltout(\POWERLED.dutycycle_eena_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_2_LC_8_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_2_LC_8_9_6 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_2_LC_8_9_6 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \POWERLED.dutycycle_2_LC_8_9_6  (
            .in0(N__22568),
            .in1(N__22559),
            .in2(N__22562),
            .in3(N__32627),
            .lcout(\POWERLED.dutycycleZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32450),
            .ce(),
            .sr(N__31754));
    defparam \POWERLED.G_141_LC_8_9_7 .C_ON=1'b0;
    defparam \POWERLED.G_141_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_141_LC_8_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.G_141_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__25581),
            .in2(_gnd_net_),
            .in3(N__22523),
            .lcout(G_141),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_7_LC_8_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_7_LC_8_10_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_7_LC_8_10_0 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \POWERLED.dutycycle_7_LC_8_10_0  (
            .in0(N__22460),
            .in1(N__26771),
            .in2(N__32628),
            .in3(N__22454),
            .lcout(\POWERLED.dutycycleZ1Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32412),
            .ce(),
            .sr(N__31731));
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1G_LC_8_10_1 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1G_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1G_LC_8_10_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1G_LC_8_10_1  (
            .in0(N__23861),
            .in1(N__27234),
            .in2(N__30721),
            .in3(N__27623),
            .lcout(\POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1GZ0 ),
            .ltout(\POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1GZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNICSH47_7_LC_8_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNICSH47_7_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNICSH47_7_LC_8_10_2 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.dutycycle_RNICSH47_7_LC_8_10_2  (
            .in0(N__32575),
            .in1(N__22453),
            .in2(N__22445),
            .in3(N__26770),
            .lcout(\POWERLED.dutycycleZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.g0_5_LC_8_10_3 .C_ON=1'b0;
    defparam \POWERLED.g0_5_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.g0_5_LC_8_10_3 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \POWERLED.g0_5_LC_8_10_3  (
            .in0(N__30672),
            .in1(N__30288),
            .in2(_gnd_net_),
            .in3(N__27621),
            .lcout(\POWERLED.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBVNS_2_0_LC_8_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_2_0_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_2_0_LC_8_10_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.func_state_RNIBVNS_2_0_LC_8_10_6  (
            .in0(N__27622),
            .in1(N__30671),
            .in2(N__30314),
            .in3(N__28816),
            .lcout(\POWERLED.func_state_RNIBVNS_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22745),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\POWERLED.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_8_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_8_11_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22721),
            .in3(N__22712),
            .lcout(\POWERLED.mult1_un47_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_8_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_8_11_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22763),
            .in3(N__22700),
            .lcout(\POWERLED.mult1_un47_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_8_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_8_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__25195),
            .in2(N__22697),
            .in3(N__22679),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_8_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_8_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__25183),
            .in2(N__22676),
            .in3(N__22652),
            .lcout(\POWERLED.mult1_un47_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_8_11_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_8_11_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22649),
            .in3(N__22640),
            .lcout(\POWERLED.mult1_un54_sum_s_8 ),
            .ltout(\POWERLED.mult1_un54_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_8_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_8_11_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22619),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_8_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_8_11_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_8_11_7  (
            .in0(N__22869),
            .in1(N__22870),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_0_LC_8_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_0_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_0_LC_8_12_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_0_LC_8_12_0  (
            .in0(N__26552),
            .in1(N__30925),
            .in2(_gnd_net_),
            .in3(N__31400),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_LC_8_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_LC_8_12_1 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_LC_8_12_1  (
            .in0(N__31401),
            .in1(_gnd_net_),
            .in2(N__27098),
            .in3(N__31013),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNIZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_8_LC_8_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_8_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_8_LC_8_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_2_8_LC_8_12_2  (
            .in0(N__31298),
            .in1(N__31406),
            .in2(N__22838),
            .in3(N__24607),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_LC_8_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_LC_8_12_3 .LUT_INIT=16'b1100011011000110;
    LogicCell40 \POWERLED.dutycycle_RNI_2_LC_8_12_3  (
            .in0(N__30926),
            .in1(N__31297),
            .in2(N__31430),
            .in3(N__32953),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_3_LC_8_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_8_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNI_1_3_LC_8_12_4  (
            .in0(N__31014),
            .in1(N__31405),
            .in2(_gnd_net_),
            .in3(N__27073),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_12_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_12_5 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22817),
            .in3(N__22785),
            .lcout(\POWERLED.mult1_un47_sum_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_8_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_8_12_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__30927),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_7_LC_8_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_7_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_7_LC_8_12_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_7_LC_8_12_7  (
            .in0(N__27074),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30144),
            .lcout(\POWERLED.N_510 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIRPVQ5_13_LC_8_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIRPVQ5_13_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIRPVQ5_13_LC_8_13_0 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \POWERLED.dutycycle_RNIRPVQ5_13_LC_8_13_0  (
            .in0(N__24062),
            .in1(N__22915),
            .in2(N__22934),
            .in3(N__31566),
            .lcout(\POWERLED.dutycycleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_13_LC_8_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_13_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_13_LC_8_13_1 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \POWERLED.dutycycle_13_LC_8_13_1  (
            .in0(N__31567),
            .in1(N__24061),
            .in2(N__22919),
            .in3(N__22930),
            .lcout(\POWERLED.dutycycleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32466),
            .ce(),
            .sr(N__31721));
    defparam \POWERLED.dutycycle_9_LC_8_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_9_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_9_LC_8_13_2 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \POWERLED.dutycycle_9_LC_8_13_2  (
            .in0(N__23849),
            .in1(N__27248),
            .in2(N__22889),
            .in3(N__31568),
            .lcout(\POWERLED.dutycycleZ1Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32466),
            .ce(),
            .sr(N__31721));
    defparam \POWERLED.dutycycle_RNI_1_10_LC_8_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_10_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_10_LC_8_13_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_10_LC_8_13_3  (
            .in0(N__27346),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24796),
            .lcout(\POWERLED.un1_dutycycle_53_41_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_8_LC_8_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_8_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_8_LC_8_13_4 .LUT_INIT=16'b1111000011000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_8_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__27345),
            .in2(N__24618),
            .in3(N__24860),
            .lcout(\POWERLED.un1_dutycycle_53_40_0 ),
            .ltout(\POWERLED.un1_dutycycle_53_40_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_13_LC_8_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_13_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_13_LC_8_13_5 .LUT_INIT=16'b0011001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_2_13_LC_8_13_5  (
            .in0(N__24111),
            .in1(N__22907),
            .in2(N__22901),
            .in3(N__24473),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNITR8L6_9_LC_8_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNITR8L6_9_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNITR8L6_9_LC_8_13_6 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \POWERLED.dutycycle_RNITR8L6_9_LC_8_13_6  (
            .in0(N__23848),
            .in1(N__27247),
            .in2(N__22888),
            .in3(N__31565),
            .lcout(\POWERLED.dutycycleZ0Z_4 ),
            .ltout(\POWERLED.dutycycleZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_8_LC_8_13_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_8_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_8_LC_8_13_7 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_8_LC_8_13_7  (
            .in0(N__27065),
            .in1(_gnd_net_),
            .in2(N__22874),
            .in3(N__24599),
            .lcout(\POWERLED.un1_dutycycle_53_31_a5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_8_LC_8_14_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_8_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_8_LC_8_14_0 .LUT_INIT=16'b1110110011001000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_8_LC_8_14_0  (
            .in0(N__31020),
            .in1(N__31425),
            .in2(N__27106),
            .in3(N__24604),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_8 ),
            .ltout(\POWERLED.dutycycle_RNI_0Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_LC_8_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_LC_8_14_1 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_LC_8_14_1  (
            .in0(N__27341),
            .in1(_gnd_net_),
            .in2(N__22994),
            .in3(N__31149),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNIZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_7_LC_8_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_7_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_7_LC_8_14_2 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \POWERLED.dutycycle_RNI_1_7_LC_8_14_2  (
            .in0(N__27096),
            .in1(N__31148),
            .in2(N__22991),
            .in3(N__24794),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_5_LC_8_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_5_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_5_LC_8_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNI_0_5_LC_8_14_3  (
            .in0(N__27342),
            .in1(N__31150),
            .in2(N__31322),
            .in3(N__22982),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_4_LC_8_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_4_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_4_LC_8_14_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \POWERLED.dutycycle_RNI_0_4_LC_8_14_4  (
            .in0(N__24425),
            .in1(N__31424),
            .in2(_gnd_net_),
            .in3(N__27340),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_31_a4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_6_LC_8_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_6_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_6_LC_8_14_5 .LUT_INIT=16'b0001000100011011;
    LogicCell40 \POWERLED.dutycycle_RNI_1_6_LC_8_14_5  (
            .in0(N__31147),
            .in1(N__22958),
            .in2(N__22967),
            .in3(N__22964),
            .lcout(\POWERLED.un1_dutycycle_53_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_8_LC_8_14_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_8_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_8_LC_8_14_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_9_8_LC_8_14_6  (
            .in0(N__31019),
            .in1(N__31423),
            .in2(N__27105),
            .in3(N__24603),
            .lcout(\POWERLED.un1_dutycycle_53_31_a0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_12_LC_8_14_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_12_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_12_LC_8_14_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNI_12_LC_8_14_7  (
            .in0(N__27343),
            .in1(N__26963),
            .in2(N__24368),
            .in3(N__24608),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNITTAN6_14_LC_8_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNITTAN6_14_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNITTAN6_14_LC_8_15_0 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \POWERLED.dutycycle_RNITTAN6_14_LC_8_15_0  (
            .in0(N__22942),
            .in1(N__27913),
            .in2(N__23960),
            .in3(N__31583),
            .lcout(\POWERLED.dutycycleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_14_LC_8_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_14_LC_8_15_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_14_LC_8_15_1 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \POWERLED.dutycycle_14_LC_8_15_1  (
            .in0(N__31585),
            .in1(N__23956),
            .in2(N__27917),
            .in3(N__22943),
            .lcout(\POWERLED.dutycycleZ1Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32472),
            .ce(),
            .sr(N__31781));
    defparam \POWERLED.dutycycle_15_LC_8_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_15_LC_8_15_2 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_15_LC_8_15_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \POWERLED.dutycycle_15_LC_8_15_2  (
            .in0(N__27962),
            .in1(N__31586),
            .in2(N__23054),
            .in3(N__23935),
            .lcout(\POWERLED.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32472),
            .ce(),
            .sr(N__31781));
    defparam \POWERLED.dutycycle_RNI_12_8_LC_8_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_12_8_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_12_8_LC_8_15_3 .LUT_INIT=16'b1010101000100000;
    LogicCell40 \POWERLED.dutycycle_RNI_12_8_LC_8_15_3  (
            .in0(N__24866),
            .in1(N__24332),
            .in2(N__24542),
            .in3(N__24472),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_12Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_15_LC_8_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_15_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_15_LC_8_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_15_LC_8_15_4  (
            .in0(N__27512),
            .in1(N__26952),
            .in2(N__23066),
            .in3(N__24677),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIV0CN6_15_LC_8_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIV0CN6_15_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIV0CN6_15_LC_8_15_5 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \POWERLED.dutycycle_RNIV0CN6_15_LC_8_15_5  (
            .in0(N__31584),
            .in1(N__23050),
            .in2(N__23936),
            .in3(N__27961),
            .lcout(\POWERLED.dutycycleZ0Z_14 ),
            .ltout(\POWERLED.dutycycleZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_15_LC_8_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_8_15_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_15_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23042),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_2381_i ),
            .ltout(\POWERLED.N_2381_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_14_LC_8_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_14_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_14_LC_8_15_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_14_LC_8_15_7  (
            .in0(N__24678),
            .in1(N__27754),
            .in2(N__23039),
            .in3(N__29335),
            .lcout(\POWERLED.un2_count_clk_17_0_0_a2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_11_LC_8_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_11_LC_8_16_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_11_LC_8_16_0 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \POWERLED.dutycycle_11_LC_8_16_0  (
            .in0(N__23009),
            .in1(N__23020),
            .in2(N__31592),
            .in3(N__24137),
            .lcout(\POWERLED.dutycycleZ1Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32479),
            .ce(),
            .sr(N__31750));
    defparam \POWERLED.dutycycle_RNI_13_LC_8_16_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_13_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_13_LC_8_16_2 .LUT_INIT=16'b1010101001011010;
    LogicCell40 \POWERLED.dutycycle_RNI_13_LC_8_16_2  (
            .in0(N__24113),
            .in1(N__27755),
            .in2(N__23108),
            .in3(N__24449),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIFDK47_11_LC_8_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIFDK47_11_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIFDK47_11_LC_8_16_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \POWERLED.dutycycle_RNIFDK47_11_LC_8_16_3  (
            .in0(N__24136),
            .in1(N__31575),
            .in2(N__23021),
            .in3(N__23008),
            .lcout(\POWERLED.dutycycleZ0Z_9 ),
            .ltout(\POWERLED.dutycycleZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_11_LC_8_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_8_16_4 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \POWERLED.dutycycle_RNI_2_11_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23114),
            .in3(N__24767),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_2Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_12_LC_8_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_8_16_5 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \POWERLED.dutycycle_RNI_3_12_LC_8_16_5  (
            .in0(N__24348),
            .in1(N__26978),
            .in2(N__23111),
            .in3(N__24442),
            .lcout(\POWERLED.un1_dutycycle_53_2_1 ),
            .ltout(\POWERLED.un1_dutycycle_53_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_13_LC_8_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_8_16_6 .LUT_INIT=16'b1010000000100000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_13_LC_8_16_6  (
            .in0(N__24112),
            .in1(N__24349),
            .in2(N__23099),
            .in3(N__24364),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI63141_10_LC_9_2_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_9_2_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_RNI63141_10_LC_9_2_0  (
            .in0(N__24980),
            .in1(N__25052),
            .in2(N__25523),
            .in3(N__25070),
            .lcout(),
            .ltout(\VPP_VDDQ.un6_count_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_2_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_2_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_2_1  (
            .in0(N__23078),
            .in1(N__23084),
            .in2(N__23087),
            .in3(N__23072),
            .lcout(VPP_VDDQ_un6_count),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_9_2_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_9_2_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_RNIVJP51_3_LC_9_2_2  (
            .in0(N__24998),
            .in1(N__25016),
            .in2(N__24962),
            .in3(N__25034),
            .lcout(\VPP_VDDQ.un6_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_9_2_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_9_2_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \VPP_VDDQ.count_RNIFC141_11_LC_9_2_3  (
            .in0(N__25544),
            .in1(N__24509),
            .in2(N__25499),
            .in3(N__24941),
            .lcout(\VPP_VDDQ.un6_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_2_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_2_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_2_4  (
            .in0(N__25223),
            .in1(N__25454),
            .in2(N__25103),
            .in3(N__25475),
            .lcout(\VPP_VDDQ.un6_count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNIMTB22_0_LC_9_3_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNIMTB22_0_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNIMTB22_0_LC_9_3_1 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \VPP_VDDQ.curr_state_RNIMTB22_0_LC_9_3_1  (
            .in0(N__23339),
            .in1(N__23289),
            .in2(_gnd_net_),
            .in3(N__23251),
            .lcout(\VPP_VDDQ.N_64_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_1_LC_9_3_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_1_LC_9_3_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_1_LC_9_3_2 .LUT_INIT=16'b0011000000111010;
    LogicCell40 \VPP_VDDQ.curr_state_1_LC_9_3_2  (
            .in0(N__23254),
            .in1(N__23360),
            .in2(N__23302),
            .in3(N__23341),
            .lcout(VPP_VDDQ_curr_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32280),
            .ce(N__25316),
            .sr(_gnd_net_));
    defparam \POWERLED.G_30_0_LC_9_3_4 .C_ON=1'b0;
    defparam \POWERLED.G_30_0_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_30_0_LC_9_3_4 .LUT_INIT=16'b0101011100000000;
    LogicCell40 \POWERLED.G_30_0_LC_9_3_4  (
            .in0(N__23252),
            .in1(N__23338),
            .in2(N__23301),
            .in3(N__25400),
            .lcout(),
            .ltout(\POWERLED.G_30Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_30_LC_9_3_5 .C_ON=1'b0;
    defparam \POWERLED.G_30_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_30_LC_9_3_5 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \POWERLED.G_30_LC_9_3_5  (
            .in0(N__23297),
            .in1(N__23253),
            .in2(N__23363),
            .in3(N__23359),
            .lcout(G_30),
            .ltout(G_30_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_9_3_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_9_3_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \VPP_VDDQ.count_esr_RNO_0_15_LC_9_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23348),
            .in3(N__25401),
            .lcout(\VPP_VDDQ.N_92_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_0_LC_9_3_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_0_LC_9_3_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_0_LC_9_3_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \VPP_VDDQ.curr_state_0_LC_9_3_7  (
            .in0(N__23340),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23296),
            .lcout(VPP_VDDQ_curr_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32280),
            .ce(N__25316),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_3_LC_9_4_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_3_LC_9_4_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_3_LC_9_4_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_off_3_LC_9_4_0  (
            .in0(N__26100),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23224),
            .lcout(\POWERLED.count_off_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32269),
            .ce(N__23519),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIBHMIG_3_LC_9_4_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIBHMIG_3_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIBHMIG_3_LC_9_4_1 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \POWERLED.count_off_RNIBHMIG_3_LC_9_4_1  (
            .in0(N__23234),
            .in1(N__23511),
            .in2(N__23228),
            .in3(N__26097),
            .lcout(\POWERLED.count_offZ0Z_3 ),
            .ltout(\POWERLED.count_offZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_3_LC_9_4_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_3_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_3_LC_9_4_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_3_LC_9_4_2  (
            .in0(N__23198),
            .in1(N__23602),
            .in2(N__23174),
            .in3(N__23171),
            .lcout(),
            .ltout(\POWERLED.un34_clk_100khz_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_0_10_LC_9_4_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_0_10_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_0_10_LC_9_4_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.count_off_RNI_0_10_LC_9_4_3  (
            .in0(N__23144),
            .in1(N__23138),
            .in2(N__23126),
            .in3(N__23123),
            .lcout(\POWERLED.count_off_RNI_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIDKNIG_4_LC_9_4_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIDKNIG_4_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIDKNIG_4_LC_9_4_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \POWERLED.count_off_RNIDKNIG_4_LC_9_4_4  (
            .in0(N__26098),
            .in1(N__23570),
            .in2(N__23539),
            .in3(N__23588),
            .lcout(\POWERLED.count_offZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_4_LC_9_4_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_4_LC_9_4_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_4_LC_9_4_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_off_4_LC_9_4_5  (
            .in0(_gnd_net_),
            .in1(N__23587),
            .in2(_gnd_net_),
            .in3(N__26101),
            .lcout(\POWERLED.count_off_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32269),
            .ce(N__23519),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_1_LC_9_4_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_1_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_1_LC_9_4_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_off_1_LC_9_4_6  (
            .in0(N__26099),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23563),
            .lcout(\POWERLED.count_off_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32269),
            .ce(N__23519),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIH5L3G_1_LC_9_4_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIH5L3G_1_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIH5L3G_1_LC_9_4_7 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \POWERLED.count_off_RNIH5L3G_1_LC_9_4_7  (
            .in0(N__23564),
            .in1(N__23552),
            .in2(N__23540),
            .in3(N__26096),
            .lcout(\POWERLED.count_offZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_S3n_RNI5DLR_LC_9_5_0.C_ON=1'b0;
    defparam SLP_S3n_RNI5DLR_LC_9_5_0.SEQ_MODE=4'b0000;
    defparam SLP_S3n_RNI5DLR_LC_9_5_0.LUT_INIT=16'b1001100111111111;
    LogicCell40 SLP_S3n_RNI5DLR_LC_9_5_0 (
            .in0(N__30354),
            .in1(N__30734),
            .in2(_gnd_net_),
            .in3(N__28850),
            .lcout(),
            .ltout(N_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_fast_RNI8TRB2_LC_9_5_1 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_fast_RNI8TRB2_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_0_fast_RNI8TRB2_LC_9_5_1 .LUT_INIT=16'b1101000011110010;
    LogicCell40 \COUNTER.tmp_0_fast_RNI8TRB2_LC_9_5_1  (
            .in0(N__26734),
            .in1(N__26342),
            .in2(N__23372),
            .in3(N__23655),
            .lcout(),
            .ltout(N_8_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep2_RNIDD505_LC_9_5_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep2_RNIDD505_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep2_RNIDD505_LC_9_5_2 .LUT_INIT=16'b0000001000110011;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_rep2_RNIDD505_LC_9_5_2  (
            .in0(N__29893),
            .in1(N__23627),
            .in2(N__23369),
            .in3(N__30118),
            .lcout(POWERLED_g2_1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.g0_5_1_LC_9_5_3 .C_ON=1'b0;
    defparam \POWERLED.g0_5_1_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.g0_5_1_LC_9_5_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.g0_5_1_LC_9_5_3  (
            .in0(N__30733),
            .in1(N__30353),
            .in2(N__26754),
            .in3(N__27177),
            .lcout(),
            .ltout(\POWERLED.g0_5Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIA2VR1_0_LC_9_5_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIA2VR1_0_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIA2VR1_0_LC_9_5_4 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \POWERLED.func_state_RNIA2VR1_0_LC_9_5_4  (
            .in0(N__25580),
            .in1(N__25866),
            .in2(N__23366),
            .in3(N__28849),
            .lcout(),
            .ltout(\POWERLED.N_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIUKM0G_1_LC_9_5_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIUKM0G_1_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIUKM0G_1_LC_9_5_5 .LUT_INIT=16'b0000100000111011;
    LogicCell40 \POWERLED.func_state_RNIUKM0G_1_LC_9_5_5  (
            .in0(N__23699),
            .in1(N__23693),
            .in2(N__23681),
            .in3(N__23663),
            .lcout(\POWERLED.func_state_1_m2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIGN2N5_1_LC_9_5_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIGN2N5_1_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIGN2N5_1_LC_9_5_6 .LUT_INIT=16'b0011001100110111;
    LogicCell40 \POWERLED.func_state_RNIGN2N5_1_LC_9_5_6  (
            .in0(N__23669),
            .in1(N__25867),
            .in2(N__23639),
            .in3(N__23786),
            .lcout(\POWERLED.func_state_1_m2_N_3_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.g0_17_LC_9_5_7 .C_ON=1'b0;
    defparam \POWERLED.g0_17_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.g0_17_LC_9_5_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.g0_17_LC_9_5_7  (
            .in0(N__26735),
            .in1(N__23654),
            .in2(N__26365),
            .in3(N__27176),
            .lcout(\POWERLED.N_671_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_S3n_RNI5DLR_0_LC_9_6_0.C_ON=1'b0;
    defparam SLP_S3n_RNI5DLR_0_LC_9_6_0.SEQ_MODE=4'b0000;
    defparam SLP_S3n_RNI5DLR_0_LC_9_6_0.LUT_INIT=16'b0011000011000000;
    LogicCell40 SLP_S3n_RNI5DLR_0_LC_9_6_0 (
            .in0(_gnd_net_),
            .in1(N__30352),
            .in2(N__26239),
            .in3(N__30732),
            .lcout(),
            .ltout(G_7_i_a4_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_RNI75Q52_LC_9_6_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_RNI75Q52_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_RNI75Q52_LC_9_6_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_rep1_RNI75Q52_LC_9_6_1  (
            .in0(N__27172),
            .in1(N__26285),
            .in2(N__23630),
            .in3(N__26349),
            .lcout(\RSMRST_PWRGD.G_7_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIPGQN2_4_3_LC_9_6_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIPGQN2_4_3_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIPGQN2_4_3_LC_9_6_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.count_clk_RNIPGQN2_4_3_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__28133),
            .in2(_gnd_net_),
            .in3(N__28112),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2MQD_0_LC_9_6_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2MQD_0_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2MQD_0_LC_9_6_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.func_state_RNI2MQD_0_LC_9_6_3  (
            .in0(N__30348),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26231),
            .lcout(\POWERLED.N_533 ),
            .ltout(\POWERLED.N_533_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI98AF2_1_LC_9_6_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI98AF2_1_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI98AF2_1_LC_9_6_4 .LUT_INIT=16'b0011001100110000;
    LogicCell40 \POWERLED.func_state_RNI98AF2_1_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__23612),
            .in2(N__23621),
            .in3(N__27171),
            .lcout(\POWERLED.un1_clk_100khz_51_and_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIA70J1_1_LC_9_6_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIA70J1_1_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIA70J1_1_LC_9_6_5 .LUT_INIT=16'b0000010100010101;
    LogicCell40 \POWERLED.func_state_RNIA70J1_1_LC_9_6_5  (
            .in0(N__23618),
            .in1(N__29655),
            .in2(N__30377),
            .in3(N__29726),
            .lcout(\POWERLED.un1_clk_100khz_51_and_i_3_0_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOI5P1_0_5_LC_9_6_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOI5P1_0_5_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOI5P1_0_5_LC_9_6_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \POWERLED.dutycycle_RNIOI5P1_0_5_LC_9_6_6  (
            .in0(N__23747),
            .in1(N__29423),
            .in2(N__25969),
            .in3(N__25934),
            .lcout(\POWERLED.un1_dutycycle_172_m3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_3_1_LC_9_6_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_3_1_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_3_1_LC_9_6_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.func_state_RNI_3_1_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(N__25865),
            .in2(_gnd_net_),
            .in3(N__30115),
            .lcout(\POWERLED.func_state_RNI_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI1TUN2_7_LC_9_7_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI1TUN2_7_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI1TUN2_7_LC_9_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNI1TUN2_7_LC_9_7_0  (
            .in0(N__29099),
            .in1(N__23720),
            .in2(_gnd_net_),
            .in3(N__28264),
            .lcout(\POWERLED.count_clkZ0Z_7 ),
            .ltout(\POWERLED.count_clkZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_0_LC_9_7_1 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_0_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_0_LC_9_7_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_0_LC_9_7_1  (
            .in0(N__30116),
            .in1(N__23728),
            .in2(N__23741),
            .in3(N__28624),
            .lcout(\POWERLED.un1_func_state25_6_0_o_N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIPGQN2_7_LC_9_7_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIPGQN2_7_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIPGQN2_7_LC_9_7_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.count_clk_RNIPGQN2_7_LC_9_7_2  (
            .in0(N__23729),
            .in1(N__28300),
            .in2(N__28628),
            .in3(N__26281),
            .lcout(\POWERLED.N_490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_7_LC_9_7_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_7_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_7_LC_9_7_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_7_LC_9_7_3  (
            .in0(N__28265),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32385),
            .ce(N__29117),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_5_LC_9_7_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_5_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_5_LC_9_7_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \POWERLED.dutycycle_RNI_2_5_LC_9_7_4  (
            .in0(N__31308),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30117),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_2Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIV0AS_5_LC_9_7_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIV0AS_5_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIV0AS_5_LC_9_7_5 .LUT_INIT=16'b0010011100000101;
    LogicCell40 \POWERLED.dutycycle_RNIV0AS_5_LC_9_7_5  (
            .in0(N__29536),
            .in1(N__23819),
            .in2(N__23714),
            .in3(N__29408),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_52_and_i_0_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIGV3L6_5_LC_9_7_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIGV3L6_5_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIGV3L6_5_LC_9_7_6 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \POWERLED.dutycycle_RNIGV3L6_5_LC_9_7_6  (
            .in0(N__23711),
            .in1(N__23774),
            .in2(N__23702),
            .in3(N__29537),
            .lcout(),
            .ltout(\POWERLED.N_448_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIS28SB_1_LC_9_7_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIS28SB_1_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIS28SB_1_LC_9_7_7 .LUT_INIT=16'b1010001000000000;
    LogicCell40 \POWERLED.func_state_RNIS28SB_1_LC_9_7_7  (
            .in0(N__23768),
            .in1(N__32740),
            .in2(N__23789),
            .in3(N__32593),
            .lcout(\POWERLED.func_state_RNIS28SBZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2O4A1_0_LC_9_8_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2O4A1_0_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2O4A1_0_LC_9_8_0 .LUT_INIT=16'b0100100000000000;
    LogicCell40 \POWERLED.func_state_RNI2O4A1_0_LC_9_8_0  (
            .in0(N__30696),
            .in1(N__27173),
            .in2(N__30347),
            .in3(N__26230),
            .lcout(\POWERLED.N_656_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_LC_9_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_LC_9_8_1 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \POWERLED.dutycycle_RNI_5_LC_9_8_1  (
            .in0(N__31589),
            .in1(N__28801),
            .in2(_gnd_net_),
            .in3(N__31306),
            .lcout(),
            .ltout(\POWERLED.N_133_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQAA33_0_5_LC_9_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQAA33_0_5_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQAA33_0_5_LC_9_8_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \POWERLED.dutycycle_RNIQAA33_0_5_LC_9_8_2  (
            .in0(N__23815),
            .in1(_gnd_net_),
            .in2(N__23777),
            .in3(N__23756),
            .lcout(\POWERLED.un1_dutycycle_172_m4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIO5723_1_LC_9_8_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIO5723_1_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIO5723_1_LC_9_8_3 .LUT_INIT=16'b1100110111111111;
    LogicCell40 \POWERLED.func_state_RNIO5723_1_LC_9_8_3  (
            .in0(N__29699),
            .in1(N__29573),
            .in2(N__29668),
            .in3(N__32745),
            .lcout(\POWERLED.dutycycle_eena_14_c ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_2_LC_9_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_2_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_2_LC_9_8_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_2_LC_9_8_4  (
            .in0(N__30318),
            .in1(N__30709),
            .in2(N__32956),
            .in3(N__27174),
            .lcout(),
            .ltout(\POWERLED.N_488_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQAA33_5_LC_9_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQAA33_5_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQAA33_5_LC_9_8_5 .LUT_INIT=16'b1011101110111000;
    LogicCell40 \POWERLED.dutycycle_RNIQAA33_5_LC_9_8_5  (
            .in0(N__25946),
            .in1(N__26627),
            .in2(N__23759),
            .in3(N__31305),
            .lcout(\POWERLED.un1_dutycycle_172_m2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2MQD_0_1_LC_9_8_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2MQD_0_1_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2MQD_0_1_LC_9_8_6 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \POWERLED.func_state_RNI2MQD_0_1_LC_9_8_6  (
            .in0(N__28800),
            .in1(N__30061),
            .in2(N__30346),
            .in3(N__28923),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_30_and_i_0_0_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIV0AS_1_LC_9_8_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIV0AS_1_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIV0AS_1_LC_9_8_7 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \POWERLED.func_state_RNIV0AS_1_LC_9_8_7  (
            .in0(N__28924),
            .in1(_gnd_net_),
            .in2(N__23750),
            .in3(N__27175),
            .lcout(\POWERLED.N_91_1_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_5_LC_9_9_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_5_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_5_LC_9_9_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_5_LC_9_9_0  (
            .in0(N__31145),
            .in1(N__29355),
            .in2(N__31307),
            .in3(N__30781),
            .lcout(\POWERLED.func_state_1_m2s2_i_0_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_8_1_LC_9_9_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_8_1_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_8_1_LC_9_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_8_1_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27227),
            .lcout(\POWERLED.func_state_RNI_8Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_6_1_LC_9_9_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_6_1_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_6_1_LC_9_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_6_1_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29274),
            .lcout(\POWERLED.N_435_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI02AS_0_1_LC_9_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI02AS_0_1_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI02AS_0_1_LC_9_9_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.func_state_RNI02AS_0_1_LC_9_9_3  (
            .in0(N__30694),
            .in1(N__28841),
            .in2(N__27185),
            .in3(N__27228),
            .lcout(\POWERLED.count_off_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_LC_9_9_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_LC_9_9_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_LC_9_9_4  (
            .in0(N__30928),
            .in1(N__29275),
            .in2(N__29230),
            .in3(N__26553),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_96_0_a3_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_3_LC_9_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_9_9_5 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \POWERLED.dutycycle_RNI_0_3_LC_9_9_5  (
            .in0(N__26623),
            .in1(N__31024),
            .in2(N__23822),
            .in3(N__31432),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_clk_100khz_32_and_i_0_o2_0_LC_9_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_clk_100khz_32_and_i_0_o2_0_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_clk_100khz_32_and_i_0_o2_0_LC_9_9_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \POWERLED.un1_clk_100khz_32_and_i_0_o2_0_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__30695),
            .in2(_gnd_net_),
            .in3(N__26755),
            .lcout(\POWERLED.N_251 ),
            .ltout(\POWERLED.N_251_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6SKJ1_10_LC_9_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6SKJ1_10_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6SKJ1_10_LC_9_9_7 .LUT_INIT=16'b1010001000100010;
    LogicCell40 \POWERLED.dutycycle_RNI6SKJ1_10_LC_9_9_7  (
            .in0(N__30317),
            .in1(N__24793),
            .in2(N__23804),
            .in3(N__29892),
            .lcout(\POWERLED.N_506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_0_LC_9_10_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_3_0_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_0_LC_9_10_0 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_0_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26547),
            .in3(N__30905),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_0 ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNIE9MT_LC_9_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNIE9MT_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNIE9MT_LC_9_10_1 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_RNIE9MT_LC_9_10_1  (
            .in0(N__26578),
            .in1(N__24029),
            .in2(N__30924),
            .in3(N__23792),
            .lcout(\POWERLED.g0_i_m2_rn_1_0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__24010),
            .in2(N__32940),
            .in3(N__23876),
            .lcout(\POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__31018),
            .in2(N__24036),
            .in3(N__23873),
            .lcout(\POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__31431),
            .in2(N__24042),
            .in3(N__23870),
            .lcout(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__31310),
            .in2(N__24038),
            .in3(N__23867),
            .lcout(\POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_4 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_9_10_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_9_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__24014),
            .in2(N__31146),
            .in3(N__23864),
            .lcout(\POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_10_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__27075),
            .in2(N__24037),
            .in3(N__23855),
            .lcout(\POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__24619),
            .in2(N__24044),
            .in3(N__23852),
            .lcout(\POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_9_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_9_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__27354),
            .in2(N__24039),
            .in3(N__23837),
            .lcout(\POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_8 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_9_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_9_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__24022),
            .in2(N__24814),
            .in3(N__23834),
            .lcout(\POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_9_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_9_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__24705),
            .in2(N__24040),
            .in3(N__24122),
            .lcout(\POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_11_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_9_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_9_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__24021),
            .in2(N__26977),
            .in3(N__24119),
            .lcout(\POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_11_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_9_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_9_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__24116),
            .in2(N__24041),
            .in3(N__24047),
            .lcout(\POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_13_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_9_11_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_9_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__27770),
            .in2(N__24043),
            .in3(N__23942),
            .lcout(\POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_13_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_9_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_9_11_7 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_9_11_7  (
            .in0(N__27524),
            .in1(_gnd_net_),
            .in2(N__29294),
            .in3(N__23939),
            .lcout(\POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.VCCST_EN_i_1_i_LC_9_12_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.VCCST_EN_i_1_i_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.VCCST_EN_i_1_i_LC_9_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \PCH_PWRGD.VCCST_EN_i_1_i_LC_9_12_1  (
            .in0(N__27672),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30666),
            .lcout(vccst_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIP1UT_4_LC_9_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIP1UT_4_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIP1UT_4_LC_9_12_3 .LUT_INIT=16'b1100111101010101;
    LogicCell40 \POWERLED.dutycycle_RNIP1UT_4_LC_9_12_3  (
            .in0(N__24222),
            .in1(N__31564),
            .in2(N__23900),
            .in3(N__32607),
            .lcout(\POWERLED.dutycycle_RNIP1UTZ0Z_4 ),
            .ltout(\POWERLED.dutycycle_RNIP1UTZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIDH8E6_4_LC_9_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIDH8E6_4_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIDH8E6_4_LC_9_12_4 .LUT_INIT=16'b0000111110001101;
    LogicCell40 \POWERLED.dutycycle_RNIDH8E6_4_LC_9_12_4  (
            .in0(N__32834),
            .in1(N__24223),
            .in2(N__23888),
            .in3(N__24239),
            .lcout(\POWERLED.dutycycleZ0Z_5 ),
            .ltout(\POWERLED.dutycycleZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_LC_9_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_LC_9_12_5 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__31122),
            .in2(N__24242),
            .in3(N__27355),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIF86R3_4_LC_9_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIF86R3_4_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIF86R3_4_LC_9_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.dutycycle_RNIF86R3_4_LC_9_12_6  (
            .in0(N__27932),
            .in1(N__26900),
            .in2(N__27457),
            .in3(N__29812),
            .lcout(\POWERLED.dutycycle_RNIF86R3Z0Z_4 ),
            .ltout(\POWERLED.dutycycle_RNIF86R3Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_4_LC_9_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_4_LC_9_12_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_4_LC_9_12_7 .LUT_INIT=16'b0011101000110011;
    LogicCell40 \POWERLED.dutycycle_4_LC_9_12_7  (
            .in0(N__24224),
            .in1(N__24233),
            .in2(N__24227),
            .in3(N__32835),
            .lcout(\POWERLED.dutycycleZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32419),
            .ce(),
            .sr(N__31757));
    defparam \POWERLED.dutycycle_8_LC_9_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_8_LC_9_13_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_8_LC_9_13_0 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \POWERLED.dutycycle_8_LC_9_13_0  (
            .in0(N__24164),
            .in1(N__24175),
            .in2(N__31563),
            .in3(N__24188),
            .lcout(\POWERLED.dutycycleZ1Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32449),
            .ce(),
            .sr(N__31771));
    defparam \POWERLED.dutycycle_RNI_3_8_LC_9_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_8_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_8_LC_9_13_1 .LUT_INIT=16'b1010111111111010;
    LogicCell40 \POWERLED.dutycycle_RNI_3_8_LC_9_13_1  (
            .in0(N__24606),
            .in1(_gnd_net_),
            .in2(N__27097),
            .in3(N__31144),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_31_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_11_LC_9_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_9_13_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_11_LC_9_13_2  (
            .in0(N__24143),
            .in1(N__24706),
            .in2(N__24212),
            .in3(N__24209),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIRNTO5_8_LC_9_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIRNTO5_8_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIRNTO5_8_LC_9_13_3 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \POWERLED.dutycycle_RNIRNTO5_8_LC_9_13_3  (
            .in0(N__24187),
            .in1(N__31508),
            .in2(N__24179),
            .in3(N__24163),
            .lcout(\POWERLED.dutycycleZ0Z_3 ),
            .ltout(\POWERLED.dutycycleZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_8_LC_9_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_8_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_8_LC_9_13_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_6_8_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24149),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_10_8 ),
            .ltout(\POWERLED.dutycycle_RNI_10_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_8_LC_9_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_8_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_8_LC_9_13_5 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \POWERLED.dutycycle_RNI_8_8_LC_9_13_5  (
            .in0(N__24605),
            .in1(N__24320),
            .in2(N__24146),
            .in3(N__24326),
            .lcout(\POWERLED.un1_dutycycle_53_9_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_7_LC_9_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_7_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_7_LC_9_13_6 .LUT_INIT=16'b0000010111000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_7_LC_9_13_6  (
            .in0(N__27364),
            .in1(N__31399),
            .in2(N__31154),
            .in3(N__27066),
            .lcout(\POWERLED.un1_dutycycle_53_9_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_3_LC_9_13_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_9_13_7 .LUT_INIT=16'b0000001110100000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_3_LC_9_13_7  (
            .in0(N__31398),
            .in1(N__31023),
            .in2(N__27371),
            .in3(N__31140),
            .lcout(\POWERLED.un1_dutycycle_53_9_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_12_LC_9_14_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_12_LC_9_14_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_12_LC_9_14_0 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \POWERLED.dutycycle_12_LC_9_14_0  (
            .in0(N__31580),
            .in1(N__24298),
            .in2(N__26996),
            .in3(N__24314),
            .lcout(\POWERLED.dutycycleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32463),
            .ce(),
            .sr(N__31767));
    defparam \POWERLED.dutycycle_RNIHGL47_12_LC_9_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIHGL47_12_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIHGL47_12_LC_9_14_1 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \POWERLED.dutycycle_RNIHGL47_12_LC_9_14_1  (
            .in0(N__26992),
            .in1(N__24313),
            .in2(N__24299),
            .in3(N__31579),
            .lcout(\POWERLED.dutycycleZ0Z_7 ),
            .ltout(\POWERLED.dutycycleZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_12_LC_9_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_9_14_2 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \POWERLED.dutycycle_RNI_2_12_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24284),
            .in3(N__24778),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_9_a0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_8_LC_9_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_8_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_8_LC_9_14_3 .LUT_INIT=16'b1101111100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_11_8_LC_9_14_3  (
            .in0(N__24427),
            .in1(N__24468),
            .in2(N__24281),
            .in3(N__24830),
            .lcout(\POWERLED.un1_dutycycle_53_10_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_14_LC_9_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_14_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_14_LC_9_14_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_1_14_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__27743),
            .in2(_gnd_net_),
            .in3(N__24700),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_11_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_10_LC_9_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_10_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_10_LC_9_14_5 .LUT_INIT=16'b1010010111010010;
    LogicCell40 \POWERLED.dutycycle_RNI_0_10_LC_9_14_5  (
            .in0(N__24777),
            .in1(N__24266),
            .in2(N__24260),
            .in3(N__24491),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_14_LC_9_14_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_9_14_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_14_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24257),
            .in3(N__27744),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_LC_9_14_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_LC_9_14_7 .LUT_INIT=16'b1010101010100010;
    LogicCell40 \POWERLED.dutycycle_RNI_10_LC_9_14_7  (
            .in0(N__27344),
            .in1(N__24426),
            .in2(N__24795),
            .in3(N__24467),
            .lcout(\POWERLED.un1_dutycycle_53_45_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_LC_9_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_LC_9_15_0 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_LC_9_15_0  (
            .in0(N__31151),
            .in1(N__31421),
            .in2(N__27375),
            .in3(N__27085),
            .lcout(\POWERLED.un1_dutycycle_53_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_8_LC_9_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_8_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_8_LC_9_15_1 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_8_LC_9_15_1  (
            .in0(N__31422),
            .in1(N__31152),
            .in2(N__27104),
            .in3(N__24612),
            .lcout(\POWERLED.un1_dutycycle_53_35_1 ),
            .ltout(\POWERLED.un1_dutycycle_53_35_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_7_LC_9_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_7_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_7_LC_9_15_2 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_7_LC_9_15_2  (
            .in0(N__27359),
            .in1(N__24485),
            .in2(N__24476),
            .in3(N__27089),
            .lcout(\POWERLED.un1_dutycycle_53_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_6_LC_9_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_6_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_6_LC_9_15_3 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_6_LC_9_15_3  (
            .in0(N__24386),
            .in1(N__24858),
            .in2(N__24353),
            .in3(N__24377),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_6_LC_9_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_6_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_6_LC_9_15_4 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_6_LC_9_15_4  (
            .in0(N__31153),
            .in1(_gnd_net_),
            .in2(N__27376),
            .in3(N__24434),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_6 ),
            .ltout(\POWERLED.dutycycle_RNI_2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_6_LC_9_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_6_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_6_LC_9_15_5 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_6_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__24856),
            .in2(N__24380),
            .in3(N__24376),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_11_LC_9_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_9_15_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \POWERLED.dutycycle_RNI_1_11_LC_9_15_6  (
            .in0(N__27360),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24676),
            .lcout(\POWERLED.un1_dutycycle_53_50_a0_0 ),
            .ltout(\POWERLED.un1_dutycycle_53_50_a0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_11_LC_9_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_11_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_11_LC_9_15_7 .LUT_INIT=16'b0011000000110000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_11_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__24857),
            .in2(N__24335),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_dutycycle_53_50_a0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_10_LC_9_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_10_LC_9_16_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_10_LC_9_16_0 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \POWERLED.dutycycle_10_LC_9_16_0  (
            .in0(N__24919),
            .in1(N__24904),
            .in2(N__24890),
            .in3(N__31582),
            .lcout(\POWERLED.dutycycleZ1Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32480),
            .ce(),
            .sr(N__31780));
    defparam \POWERLED.dutycycle_RNI6P2N6_10_LC_9_16_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6P2N6_10_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6P2N6_10_LC_9_16_1 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \POWERLED.dutycycle_RNI6P2N6_10_LC_9_16_1  (
            .in0(N__31581),
            .in1(N__24920),
            .in2(N__24908),
            .in3(N__24886),
            .lcout(\POWERLED.dutycycleZ0Z_2 ),
            .ltout(\POWERLED.dutycycleZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_12_LC_9_16_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_9_16_2 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \POWERLED.dutycycle_RNI_4_12_LC_9_16_2  (
            .in0(N__27370),
            .in1(_gnd_net_),
            .in2(N__24878),
            .in3(N__26969),
            .lcout(\POWERLED.un2_count_clk_17_0_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_LC_9_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_LC_9_16_3 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \POWERLED.dutycycle_RNI_11_LC_9_16_3  (
            .in0(N__24748),
            .in1(N__27368),
            .in2(_gnd_net_),
            .in3(N__24696),
            .lcout(\POWERLED.un1_dutycycle_53_50_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_12_LC_9_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_9_16_4 .LUT_INIT=16'b0001010110101000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_12_LC_9_16_4  (
            .in0(N__24695),
            .in1(N__24747),
            .in2(N__27377),
            .in3(N__26968),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_10_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_8_LC_9_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_8_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_8_LC_9_16_5 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_8_LC_9_16_5  (
            .in0(N__24859),
            .in1(N__24821),
            .in2(N__24833),
            .in3(N__24613),
            .lcout(\POWERLED.un1_dutycycle_53_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_12_LC_9_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_9_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_12_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__24746),
            .in2(_gnd_net_),
            .in3(N__26967),
            .lcout(\POWERLED.un1_dutycycle_53_9_a1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_LC_9_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_LC_9_16_7 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \POWERLED.dutycycle_RNI_8_LC_9_16_7  (
            .in0(N__24749),
            .in1(N__27369),
            .in2(N__24707),
            .in3(N__24614),
            .lcout(\POWERLED.un1_dutycycle_53_50_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_0_LC_11_2_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_0_LC_11_2_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_0_LC_11_2_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_0_LC_11_2_0  (
            .in0(N__25418),
            .in1(N__24508),
            .in2(N__24533),
            .in3(N__24532),
            .lcout(\VPP_VDDQ.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_2_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_0 ),
            .clk(N__32332),
            .ce(),
            .sr(N__25801));
    defparam \VPP_VDDQ.count_1_LC_11_2_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_1_LC_11_2_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_1_LC_11_2_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_1_LC_11_2_1  (
            .in0(N__25404),
            .in1(N__25069),
            .in2(_gnd_net_),
            .in3(N__25055),
            .lcout(\VPP_VDDQ.countZ0Z_1 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_0 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_1 ),
            .clk(N__32332),
            .ce(),
            .sr(N__25801));
    defparam \VPP_VDDQ.count_2_LC_11_2_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_2_LC_11_2_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_LC_11_2_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_2_LC_11_2_2  (
            .in0(N__25419),
            .in1(N__25051),
            .in2(_gnd_net_),
            .in3(N__25037),
            .lcout(\VPP_VDDQ.countZ0Z_2 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_2 ),
            .clk(N__32332),
            .ce(),
            .sr(N__25801));
    defparam \VPP_VDDQ.count_3_LC_11_2_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_3_LC_11_2_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_3_LC_11_2_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_3_LC_11_2_3  (
            .in0(N__25405),
            .in1(N__25033),
            .in2(_gnd_net_),
            .in3(N__25019),
            .lcout(\VPP_VDDQ.countZ0Z_3 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_3 ),
            .clk(N__32332),
            .ce(),
            .sr(N__25801));
    defparam \VPP_VDDQ.count_4_LC_11_2_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_4_LC_11_2_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_4_LC_11_2_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_4_LC_11_2_4  (
            .in0(N__25420),
            .in1(N__25015),
            .in2(_gnd_net_),
            .in3(N__25001),
            .lcout(\VPP_VDDQ.countZ0Z_4 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_4 ),
            .clk(N__32332),
            .ce(),
            .sr(N__25801));
    defparam \VPP_VDDQ.count_5_LC_11_2_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_5_LC_11_2_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_5_LC_11_2_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_5_LC_11_2_5  (
            .in0(N__25406),
            .in1(N__24997),
            .in2(_gnd_net_),
            .in3(N__24983),
            .lcout(\VPP_VDDQ.countZ0Z_5 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_5 ),
            .clk(N__32332),
            .ce(),
            .sr(N__25801));
    defparam \VPP_VDDQ.count_6_LC_11_2_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_6_LC_11_2_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_6_LC_11_2_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_6_LC_11_2_6  (
            .in0(N__25421),
            .in1(N__24979),
            .in2(_gnd_net_),
            .in3(N__24965),
            .lcout(\VPP_VDDQ.countZ0Z_6 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_6 ),
            .clk(N__32332),
            .ce(),
            .sr(N__25801));
    defparam \VPP_VDDQ.count_7_LC_11_2_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_7_LC_11_2_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_7_LC_11_2_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_7_LC_11_2_7  (
            .in0(N__25407),
            .in1(N__24958),
            .in2(_gnd_net_),
            .in3(N__24944),
            .lcout(\VPP_VDDQ.countZ0Z_7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_7 ),
            .clk(N__32332),
            .ce(),
            .sr(N__25801));
    defparam \VPP_VDDQ.count_8_LC_11_3_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_8_LC_11_3_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_8_LC_11_3_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_8_LC_11_3_0  (
            .in0(N__25433),
            .in1(N__24940),
            .in2(_gnd_net_),
            .in3(N__24923),
            .lcout(\VPP_VDDQ.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_8 ),
            .clk(N__32333),
            .ce(),
            .sr(N__25800));
    defparam \VPP_VDDQ.count_9_LC_11_3_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_9_LC_11_3_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_9_LC_11_3_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_9_LC_11_3_1  (
            .in0(N__25417),
            .in1(N__25543),
            .in2(_gnd_net_),
            .in3(N__25526),
            .lcout(\VPP_VDDQ.countZ0Z_9 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_8 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_9 ),
            .clk(N__32333),
            .ce(),
            .sr(N__25800));
    defparam \VPP_VDDQ.count_10_LC_11_3_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_10_LC_11_3_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_10_LC_11_3_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_10_LC_11_3_2  (
            .in0(N__25430),
            .in1(N__25516),
            .in2(_gnd_net_),
            .in3(N__25502),
            .lcout(\VPP_VDDQ.countZ0Z_10 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_10 ),
            .clk(N__32333),
            .ce(),
            .sr(N__25800));
    defparam \VPP_VDDQ.count_11_LC_11_3_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_11_LC_11_3_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_11_LC_11_3_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_11_LC_11_3_3  (
            .in0(N__25415),
            .in1(N__25492),
            .in2(_gnd_net_),
            .in3(N__25478),
            .lcout(\VPP_VDDQ.countZ0Z_11 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_11 ),
            .clk(N__32333),
            .ce(),
            .sr(N__25800));
    defparam \VPP_VDDQ.count_12_LC_11_3_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_12_LC_11_3_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_12_LC_11_3_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_12_LC_11_3_4  (
            .in0(N__25431),
            .in1(N__25471),
            .in2(_gnd_net_),
            .in3(N__25457),
            .lcout(\VPP_VDDQ.countZ0Z_12 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_12 ),
            .clk(N__32333),
            .ce(),
            .sr(N__25800));
    defparam \VPP_VDDQ.count_13_LC_11_3_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_13_LC_11_3_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_13_LC_11_3_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_13_LC_11_3_5  (
            .in0(N__25416),
            .in1(N__25450),
            .in2(_gnd_net_),
            .in3(N__25436),
            .lcout(\VPP_VDDQ.countZ0Z_13 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_13 ),
            .clk(N__32333),
            .ce(),
            .sr(N__25800));
    defparam \VPP_VDDQ.count_14_LC_11_3_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_14_LC_11_3_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_14_LC_11_3_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_14_LC_11_3_6  (
            .in0(N__25432),
            .in1(N__25222),
            .in2(_gnd_net_),
            .in3(N__25205),
            .lcout(\VPP_VDDQ.countZ0Z_14 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14 ),
            .clk(N__32333),
            .ce(),
            .sr(N__25800));
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_3_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_3_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_3_7  (
            .in0(_gnd_net_),
            .in1(N__25180),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_14 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_15_LC_11_4_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_15_LC_11_4_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_esr_15_LC_11_4_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \VPP_VDDQ.count_esr_15_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(N__25096),
            .in2(_gnd_net_),
            .in3(N__25106),
            .lcout(\VPP_VDDQ.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32342),
            .ce(N__25082),
            .sr(N__25805));
    defparam \POWERLED.count_clk_RNIRJRN2_4_LC_11_5_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIRJRN2_4_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIRJRN2_4_LC_11_5_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNIRJRN2_4_LC_11_5_0  (
            .in0(N__25775),
            .in1(N__29060),
            .in2(_gnd_net_),
            .in3(N__28393),
            .lcout(\POWERLED.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_4_LC_11_5_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_4_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_4_LC_11_5_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_4_LC_11_5_1  (
            .in0(N__28394),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32334),
            .ce(N__29103),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNITMSN2_5_LC_11_5_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNITMSN2_5_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNITMSN2_5_LC_11_5_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNITMSN2_5_LC_11_5_2  (
            .in0(N__25769),
            .in1(N__29061),
            .in2(_gnd_net_),
            .in3(N__28357),
            .lcout(\POWERLED.count_clkZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_5_LC_11_5_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_5_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_5_LC_11_5_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_5_LC_11_5_3  (
            .in0(N__28358),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32334),
            .ce(N__29103),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIVPTN2_6_LC_11_5_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIVPTN2_6_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIVPTN2_6_LC_11_5_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNIVPTN2_6_LC_11_5_4  (
            .in0(N__25763),
            .in1(N__29062),
            .in2(_gnd_net_),
            .in3(N__28330),
            .lcout(\POWERLED.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_6_LC_11_5_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_6_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_6_LC_11_5_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_6_LC_11_5_5  (
            .in0(N__28331),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32334),
            .ce(N__29103),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIH9TE_10_LC_11_5_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIH9TE_10_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIH9TE_10_LC_11_5_6 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \POWERLED.count_off_RNIH9TE_10_LC_11_5_6  (
            .in0(N__26707),
            .in1(N__25634),
            .in2(_gnd_net_),
            .in3(N__25872),
            .lcout(\POWERLED.count_off_RNIH9TEZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8AQH_0_LC_11_5_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8AQH_0_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8AQH_0_LC_11_5_7 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \POWERLED.func_state_RNI8AQH_0_LC_11_5_7  (
            .in0(N__25586),
            .in1(N__28848),
            .in2(_gnd_net_),
            .in3(N__26708),
            .lcout(\POWERLED.func_state_RNI8AQHZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNINH2G2_11_LC_11_6_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNINH2G2_11_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNINH2G2_11_LC_11_6_0 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \POWERLED.count_clk_RNINH2G2_11_LC_11_6_0  (
            .in0(N__28168),
            .in1(N__29039),
            .in2(N__25886),
            .in3(N__28520),
            .lcout(\POWERLED.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_LC_11_6_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_LC_11_6_1 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \POWERLED.count_clk_RNI_0_LC_11_6_1  (
            .in0(N__28071),
            .in1(_gnd_net_),
            .in2(N__28546),
            .in3(N__28714),
            .lcout(),
            .ltout(\POWERLED.count_clk_RNIZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI118L2_1_LC_11_6_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI118L2_1_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI118L2_1_LC_11_6_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_clk_RNI118L2_1_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__25892),
            .in2(N__25898),
            .in3(N__29038),
            .lcout(\POWERLED.count_clkZ0Z_1 ),
            .ltout(\POWERLED.count_clkZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_1_LC_11_6_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_1_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_1_LC_11_6_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.count_clk_1_LC_11_6_3  (
            .in0(N__28522),
            .in1(_gnd_net_),
            .in2(N__25895),
            .in3(N__28716),
            .lcout(\POWERLED.count_clk_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32423),
            .ce(N__29118),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_0_LC_11_6_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_0_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_0_LC_11_6_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_0_LC_11_6_4  (
            .in0(N__28717),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28516),
            .lcout(\POWERLED.count_clk_RNI_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_11_LC_11_6_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_11_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_11_LC_11_6_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_clk_11_LC_11_6_5  (
            .in0(N__28521),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28169),
            .lcout(\POWERLED.count_clk_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32423),
            .ce(N__29118),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_0_LC_11_6_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_0_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_0_LC_11_6_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.count_clk_0_LC_11_6_6  (
            .in0(N__28715),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28523),
            .lcout(\POWERLED.count_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32423),
            .ce(N__29118),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_1_LC_11_6_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_1_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_1_LC_11_6_7 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \POWERLED.count_clk_RNI_1_LC_11_6_7  (
            .in0(N__28070),
            .in1(N__28377),
            .in2(N__28652),
            .in3(N__28209),
            .lcout(\POWERLED.count_clk_RNIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_1_LC_11_7_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_1_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_1_LC_11_7_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \POWERLED.func_state_RNI_0_1_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__30157),
            .in2(_gnd_net_),
            .in3(N__25871),
            .lcout(\POWERLED.func_state_RNI_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_1_LC_11_7_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_1_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_1_LC_11_7_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_1_LC_11_7_1  (
            .in0(N__28382),
            .in1(N__28310),
            .in2(N__28076),
            .in3(N__28214),
            .lcout(),
            .ltout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_8_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIPGQN2_3_3_LC_11_7_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIPGQN2_3_3_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIPGQN2_3_3_LC_11_7_2 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \POWERLED.count_clk_RNIPGQN2_3_3_LC_11_7_2  (
            .in0(N__28132),
            .in1(_gnd_net_),
            .in2(N__25808),
            .in3(N__28648),
            .lcout(\POWERLED.N_668 ),
            .ltout(\POWERLED.N_668_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNILPF34_3_LC_11_7_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNILPF34_3_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNILPF34_3_LC_11_7_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.count_clk_RNILPF34_3_LC_11_7_3  (
            .in0(N__26010),
            .in1(N__26384),
            .in2(N__26147),
            .in3(N__27644),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIEAAR6_0_LC_11_7_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIEAAR6_0_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIEAAR6_0_LC_11_7_4 .LUT_INIT=16'b1101110011101100;
    LogicCell40 \POWERLED.func_state_RNIEAAR6_0_LC_11_7_4  (
            .in0(N__26454),
            .in1(N__26144),
            .in2(N__26135),
            .in3(N__30153),
            .lcout(\POWERLED.N_123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2VV9A_0_LC_11_7_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2VV9A_0_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2VV9A_0_LC_11_7_5 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \POWERLED.func_state_RNI2VV9A_0_LC_11_7_5  (
            .in0(N__26386),
            .in1(N__26033),
            .in2(N__26014),
            .in3(N__26300),
            .lcout(\POWERLED.func_state_RNI2VV9A_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_1_LC_11_7_6 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_1_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_1_LC_11_7_6 .LUT_INIT=16'b0001101101010111;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_1_LC_11_7_6  (
            .in0(N__26455),
            .in1(N__25978),
            .in2(N__25921),
            .in3(N__30152),
            .lcout(\POWERLED.un1_func_state25_6_0_0_0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNINEAB6_1_LC_11_7_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNINEAB6_1_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNINEAB6_1_LC_11_7_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \POWERLED.func_state_RNINEAB6_1_LC_11_7_7  (
            .in0(N__25979),
            .in1(N__28088),
            .in2(N__30158),
            .in3(N__26385),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOI5P1_5_LC_11_8_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOI5P1_5_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOI5P1_5_LC_11_8_0 .LUT_INIT=16'b1101110111000000;
    LogicCell40 \POWERLED.dutycycle_RNIOI5P1_5_LC_11_8_0  (
            .in0(N__25970),
            .in1(N__29180),
            .in2(N__26180),
            .in3(N__31247),
            .lcout(\POWERLED.un1_dutycycle_172_m0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_2_LC_11_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_2_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_2_LC_11_8_1 .LUT_INIT=16'b0011010111110101;
    LogicCell40 \POWERLED.dutycycle_RNI_4_2_LC_11_8_1  (
            .in0(N__31248),
            .in1(N__32954),
            .in2(N__29312),
            .in3(N__28843),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_172_m1_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOGRS_2_LC_11_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOGRS_2_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOGRS_2_LC_11_8_2 .LUT_INIT=16'b1100110111000001;
    LogicCell40 \POWERLED.dutycycle_RNIOGRS_2_LC_11_8_2  (
            .in0(N__26175),
            .in1(N__29308),
            .in2(N__25937),
            .in3(N__31587),
            .lcout(\POWERLED.un1_dutycycle_172_m1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI34G9_1_LC_11_8_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI34G9_1_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI34G9_1_LC_11_8_3 .LUT_INIT=16'b1100110111001111;
    LogicCell40 \POWERLED.func_state_RNI34G9_1_LC_11_8_3  (
            .in0(N__26294),
            .in1(N__26709),
            .in2(N__25922),
            .in3(N__28844),
            .lcout(\POWERLED.count_clk_en_917_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_0_LC_11_8_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_0_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_0_LC_11_8_4 .LUT_INIT=16'b1100110000001010;
    LogicCell40 \POWERLED.func_state_RNI5DLR_0_LC_11_8_4  (
            .in0(N__28842),
            .in1(N__26456),
            .in2(N__26390),
            .in3(N__30105),
            .lcout(),
            .ltout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI19L28_0_LC_11_8_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI19L28_0_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI19L28_0_LC_11_8_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.func_state_RNI19L28_0_LC_11_8_5  (
            .in0(N__26606),
            .in1(N__26309),
            .in2(N__26303),
            .in3(N__28597),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_4_1_LC_11_8_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_4_1_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_4_1_LC_11_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_4_1_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26293),
            .lcout(func_state_RNI_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOGRS_0_LC_11_8_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOGRS_0_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOGRS_0_LC_11_8_7 .LUT_INIT=16'b1011111110110011;
    LogicCell40 \POWERLED.func_state_RNIOGRS_0_LC_11_8_7  (
            .in0(N__26457),
            .in1(N__26174),
            .in2(N__30145),
            .in3(N__26540),
            .lcout(\POWERLED.dutycycle_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_LC_11_9_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_LC_11_9_0 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \POWERLED.func_state_RNI_0_LC_11_9_0  (
            .in0(N__26192),
            .in1(N__30799),
            .in2(N__26459),
            .in3(N__30782),
            .lcout(\POWERLED.N_676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_0_LC_11_9_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_0_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_0_LC_11_9_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.func_state_RNI_0_0_LC_11_9_1  (
            .in0(N__30783),
            .in1(N__26453),
            .in2(_gnd_net_),
            .in3(N__26191),
            .lcout(func_state_RNI_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_0_LC_11_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_0_LC_11_9_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_0_LC_11_9_2  (
            .in0(N__31276),
            .in1(N__31090),
            .in2(N__30920),
            .in3(N__26508),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_0 ),
            .ltout(\POWERLED.dutycycle_RNI_4Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOGRS_0_2_LC_11_9_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOGRS_0_2_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOGRS_0_2_LC_11_9_3 .LUT_INIT=16'b0001010111111111;
    LogicCell40 \POWERLED.dutycycle_RNIOGRS_0_2_LC_11_9_3  (
            .in0(N__29395),
            .in1(N__30784),
            .in2(N__26183),
            .in3(N__26179),
            .lcout(\POWERLED.un1_count_off_1_sqmuxa_8_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_0_LC_11_9_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_0_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_0_LC_11_9_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_0_LC_11_9_4  (
            .in0(N__29456),
            .in1(N__31089),
            .in2(N__30919),
            .in3(N__26509),
            .lcout(),
            .ltout(\POWERLED.N_546_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_0_LC_11_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_0_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_0_LC_11_9_5 .LUT_INIT=16'b1100110011001101;
    LogicCell40 \POWERLED.dutycycle_RNI_7_0_LC_11_9_5  (
            .in0(N__29396),
            .in1(N__30839),
            .in2(N__26630),
            .in3(N__29292),
            .lcout(\POWERLED.dutycycle_RNI_7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_0_1_LC_11_9_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_0_1_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_0_1_LC_11_9_6 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \POWERLED.func_state_RNI5DLR_0_1_LC_11_9_6  (
            .in0(N__29222),
            .in1(N__30728),
            .in2(N__30284),
            .in3(N__30079),
            .lcout(\POWERLED.N_482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIG2F54_1_LC_11_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIG2F54_1_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIG2F54_1_LC_11_10_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.dutycycle_RNIG2F54_1_LC_11_10_0  (
            .in0(N__32640),
            .in1(N__26396),
            .in2(N__26588),
            .in3(N__26600),
            .lcout(\POWERLED.g0_i_m2_rn_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIE0E38_1_LC_11_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIE0E38_1_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIE0E38_1_LC_11_10_1 .LUT_INIT=16'b0000101011111010;
    LogicCell40 \POWERLED.dutycycle_RNIE0E38_1_LC_11_10_1  (
            .in0(N__26405),
            .in1(_gnd_net_),
            .in2(N__26471),
            .in3(N__26446),
            .lcout(\POWERLED.dutycycleZ0Z_1 ),
            .ltout(\POWERLED.dutycycleZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIIASA2_1_LC_11_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIIASA2_1_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIIASA2_1_LC_11_10_2 .LUT_INIT=16'b0101010111111101;
    LogicCell40 \POWERLED.dutycycle_RNIIASA2_1_LC_11_10_2  (
            .in0(N__32793),
            .in1(N__29604),
            .in2(N__26591),
            .in3(N__29485),
            .lcout(\POWERLED.dutycycle_eena_0_0 ),
            .ltout(\POWERLED.dutycycle_eena_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIUTUT3_1_LC_11_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIUTUT3_1_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIUTUT3_1_LC_11_10_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.func_state_RNIUTUT3_1_LC_11_10_3  (
            .in0(N__26579),
            .in1(N__30143),
            .in2(N__26564),
            .in3(N__32639),
            .lcout(\POWERLED.g0_i_m2_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIIASA2_0_LC_11_10_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIIASA2_0_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIIASA2_0_LC_11_10_4 .LUT_INIT=16'b0101010111111101;
    LogicCell40 \POWERLED.dutycycle_RNIIASA2_0_LC_11_10_4  (
            .in0(N__32792),
            .in1(N__26522),
            .in2(N__29618),
            .in3(N__29484),
            .lcout(\POWERLED.dutycycle_eena ),
            .ltout(\POWERLED.dutycycle_eena_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIP8K44_0_LC_11_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIP8K44_0_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIP8K44_0_LC_11_10_5 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \POWERLED.dutycycle_RNIP8K44_0_LC_11_10_5  (
            .in0(N__26870),
            .in1(N__26851),
            .in2(N__26561),
            .in3(N__32638),
            .lcout(\POWERLED.dutycycle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_LC_11_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_LC_11_10_6 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_1_LC_11_10_6 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \POWERLED.dutycycle_1_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__26470),
            .in2(N__26458),
            .in3(N__26404),
            .lcout(\POWERLED.dutycycleZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32462),
            .ce(),
            .sr(N__31772));
    defparam \POWERLED.dutycycle_0_LC_11_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_0_LC_11_10_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_0_LC_11_10_7 .LUT_INIT=16'b0111111101000000;
    LogicCell40 \POWERLED.dutycycle_0_LC_11_10_7  (
            .in0(N__26869),
            .in1(N__26858),
            .in2(N__32668),
            .in3(N__26852),
            .lcout(\POWERLED.dutycycleZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32462),
            .ce(),
            .sr(N__31772));
    defparam \POWERLED.dutycycle_RNI2MQD_7_LC_11_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2MQD_7_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2MQD_7_LC_11_11_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.dutycycle_RNI2MQD_7_LC_11_11_0  (
            .in0(N__30243),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27099),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_36_and_i_0_a2_c_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI7JPT2_7_LC_11_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI7JPT2_7_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI7JPT2_7_LC_11_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.dutycycle_RNI7JPT2_7_LC_11_11_1  (
            .in0(N__26786),
            .in1(N__26843),
            .in2(N__26831),
            .in3(N__27451),
            .lcout(\POWERLED.un1_clk_100khz_36_and_i_0_a2_1_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_1_LC_11_11_2 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_1_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_1_LC_11_11_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \VCCIN_PWRGD.un10_output_1_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__26828),
            .in2(_gnd_net_),
            .in3(N__29619),
            .lcout(\VCCIN_PWRGD.un10_outputZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_m1_0_a2_0_LC_11_11_3 .C_ON=1'b0;
    defparam \POWERLED.un1_m1_0_a2_0_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_m1_0_a2_0_LC_11_11_3 .LUT_INIT=16'b1100000001000000;
    LogicCell40 \POWERLED.un1_m1_0_a2_0_LC_11_11_3  (
            .in0(N__30580),
            .in1(N__30244),
            .in2(N__29912),
            .in3(N__26744),
            .lcout(\POWERLED.un1_clk_100khz_36_and_i_0_a2_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI99TE_7_LC_11_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI99TE_7_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI99TE_7_LC_11_11_4 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \POWERLED.dutycycle_RNI99TE_7_LC_11_11_4  (
            .in0(N__27666),
            .in1(N__30578),
            .in2(N__27107),
            .in3(N__27891),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_36_and_i_0_a2_1_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI48JN5_7_LC_11_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI48JN5_7_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI48JN5_7_LC_11_11_5 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \POWERLED.dutycycle_RNI48JN5_7_LC_11_11_5  (
            .in0(N__32811),
            .in1(N__26780),
            .in2(N__26774),
            .in3(N__29805),
            .lcout(\POWERLED.dutycycle_eena_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_clk_100khz_43_and_i_0_o2_0_LC_11_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_clk_100khz_43_and_i_0_o2_0_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_clk_100khz_43_and_i_0_o2_0_LC_11_11_6 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \POWERLED.un1_clk_100khz_43_and_i_0_o2_0_LC_11_11_6  (
            .in0(N__26743),
            .in1(N__30579),
            .in2(_gnd_net_),
            .in3(N__29900),
            .lcout(),
            .ltout(\POWERLED.N_249_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6SKJ1_4_LC_11_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6SKJ1_4_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6SKJ1_4_LC_11_11_7 .LUT_INIT=16'b0011101100101010;
    LogicCell40 \POWERLED.dutycycle_RNI6SKJ1_4_LC_11_11_7  (
            .in0(N__30258),
            .in1(N__31435),
            .in2(N__26633),
            .in3(N__30123),
            .lcout(\POWERLED.un1_clk_100khz_40_and_i_0_a2_1_0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2MQD_1_LC_11_12_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2MQD_1_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2MQD_1_LC_11_12_0 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \POWERLED.func_state_RNI2MQD_1_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30265),
            .in3(N__30146),
            .lcout(\POWERLED.func_state_RNI2MQDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI12AS_6_LC_11_12_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI12AS_6_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI12AS_6_LC_11_12_1 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \POWERLED.count_clk_RNI12AS_6_LC_11_12_1  (
            .in0(N__29898),
            .in1(_gnd_net_),
            .in2(N__29223),
            .in3(N__30670),
            .lcout(\POWERLED.N_203 ),
            .ltout(\POWERLED.N_203_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI12AS_0_1_LC_11_12_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI12AS_0_1_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI12AS_0_1_LC_11_12_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \POWERLED.func_state_RNI12AS_0_1_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26888),
            .in3(N__27879),
            .lcout(\POWERLED.N_531 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6SKJ1_3_LC_11_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6SKJ1_3_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6SKJ1_3_LC_11_12_4 .LUT_INIT=16'b1000101000001010;
    LogicCell40 \POWERLED.dutycycle_RNI6SKJ1_3_LC_11_12_4  (
            .in0(N__30239),
            .in1(N__29744),
            .in2(N__31022),
            .in3(N__29899),
            .lcout(),
            .ltout(\POWERLED.N_521_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5TUF2_3_LC_11_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5TUF2_3_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5TUF2_3_LC_11_12_5 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \POWERLED.dutycycle_RNI5TUF2_3_LC_11_12_5  (
            .in0(N__27442),
            .in1(N__31003),
            .in2(N__26885),
            .in3(N__30147),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_43_and_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIRUFD6_3_LC_11_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIRUFD6_3_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIRUFD6_3_LC_11_12_6 .LUT_INIT=16'b0011011100000000;
    LogicCell40 \POWERLED.dutycycle_RNIRUFD6_3_LC_11_12_6  (
            .in0(N__26879),
            .in1(N__32826),
            .in2(N__26882),
            .in3(N__32645),
            .lcout(\POWERLED.dutycycle_en_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI24KO1_3_LC_11_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI24KO1_3_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI24KO1_3_LC_11_12_7 .LUT_INIT=16'b0010101000001010;
    LogicCell40 \POWERLED.dutycycle_RNI24KO1_3_LC_11_12_7  (
            .in0(N__27880),
            .in1(N__31002),
            .in2(N__27825),
            .in3(N__33129),
            .lcout(\POWERLED.N_523 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6SKJ1_9_LC_11_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6SKJ1_9_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6SKJ1_9_LC_11_13_1 .LUT_INIT=16'b1101000001010000;
    LogicCell40 \POWERLED.dutycycle_RNI6SKJ1_9_LC_11_13_1  (
            .in0(N__27374),
            .in1(N__29914),
            .in2(N__30264),
            .in3(N__29748),
            .lcout(),
            .ltout(\POWERLED.N_503_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5TUF2_9_LC_11_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5TUF2_9_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5TUF2_9_LC_11_13_2 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \POWERLED.dutycycle_RNI5TUF2_9_LC_11_13_2  (
            .in0(N__30122),
            .in1(N__27373),
            .in2(N__26873),
            .in3(N__27456),
            .lcout(\POWERLED.dutycycle_eena_2_0_0_tz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI12AS_9_LC_11_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI12AS_9_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI12AS_9_LC_11_13_3 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \POWERLED.dutycycle_RNI12AS_9_LC_11_13_3  (
            .in0(N__27372),
            .in1(N__29913),
            .in2(_gnd_net_),
            .in3(N__30720),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_30_and_i_0_a2_5_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI24KO1_9_LC_11_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI24KO1_9_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI24KO1_9_LC_11_13_4 .LUT_INIT=16'b1010111010101110;
    LogicCell40 \POWERLED.dutycycle_RNI24KO1_9_LC_11_13_4  (
            .in0(N__27206),
            .in1(N__27810),
            .in2(N__27260),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.dutycycle_eena_2_d_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIRUFD6_9_LC_11_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIRUFD6_9_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIRUFD6_9_LC_11_13_5 .LUT_INIT=16'b1011001100000000;
    LogicCell40 \POWERLED.dutycycle_RNIRUFD6_9_LC_11_13_5  (
            .in0(N__27257),
            .in1(N__32827),
            .in2(N__27251),
            .in3(N__32646),
            .lcout(\POWERLED.dutycycle_RNIRUFD6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI02AS_1_LC_11_13_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI02AS_1_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI02AS_1_LC_11_13_7 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \POWERLED.func_state_RNI02AS_1_LC_11_13_7  (
            .in0(N__30687),
            .in1(N__27205),
            .in2(_gnd_net_),
            .in3(N__27184),
            .lcout(\POWERLED.N_421 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_3_LC_11_14_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_11_14_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.dutycycle_RNI_5_3_LC_11_14_0  (
            .in0(N__31434),
            .in1(N__27103),
            .in2(_gnd_net_),
            .in3(N__31021),
            .lcout(\POWERLED.N_604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI24KO1_12_LC_11_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI24KO1_12_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI24KO1_12_LC_11_14_3 .LUT_INIT=16'b0100000011110000;
    LogicCell40 \POWERLED.dutycycle_RNI24KO1_12_LC_11_14_3  (
            .in0(N__26974),
            .in1(N__33130),
            .in2(N__27901),
            .in3(N__27819),
            .lcout(),
            .ltout(\POWERLED.N_520_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIRUFD6_12_LC_11_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIRUFD6_12_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIRUFD6_12_LC_11_14_4 .LUT_INIT=16'b0011011100000000;
    LogicCell40 \POWERLED.dutycycle_RNIRUFD6_12_LC_11_14_4  (
            .in0(N__26906),
            .in1(N__32831),
            .in2(N__26999),
            .in3(N__32669),
            .lcout(\POWERLED.dutycycle_RNIRUFD6Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6SKJ1_12_LC_11_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6SKJ1_12_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6SKJ1_12_LC_11_14_5 .LUT_INIT=16'b1100010001000100;
    LogicCell40 \POWERLED.dutycycle_RNI6SKJ1_12_LC_11_14_5  (
            .in0(N__26976),
            .in1(N__30235),
            .in2(N__29759),
            .in3(N__29915),
            .lcout(),
            .ltout(\POWERLED.N_518_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5TUF2_12_LC_11_14_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5TUF2_12_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5TUF2_12_LC_11_14_6 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \POWERLED.dutycycle_RNI5TUF2_12_LC_11_14_6  (
            .in0(N__30149),
            .in1(N__26975),
            .in2(N__26909),
            .in3(N__27458),
            .lcout(\POWERLED.un1_clk_100khz_42_and_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI99TE_4_LC_11_14_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI99TE_4_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI99TE_4_LC_11_14_7 .LUT_INIT=16'b0000001000100010;
    LogicCell40 \POWERLED.dutycycle_RNI99TE_4_LC_11_14_7  (
            .in0(N__27893),
            .in1(N__31433),
            .in2(N__30665),
            .in3(N__27673),
            .lcout(\POWERLED.un1_clk_100khz_40_and_i_0_a2_1_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI24KO1_14_LC_11_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI24KO1_14_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI24KO1_14_LC_11_15_0 .LUT_INIT=16'b0100000011110000;
    LogicCell40 \POWERLED.dutycycle_RNI24KO1_14_LC_11_15_0  (
            .in0(N__27767),
            .in1(N__33128),
            .in2(N__27902),
            .in3(N__27832),
            .lcout(),
            .ltout(\POWERLED.N_526_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI36306_14_LC_11_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI36306_14_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI36306_14_LC_11_15_1 .LUT_INIT=16'b0011011100000000;
    LogicCell40 \POWERLED.dutycycle_RNI36306_14_LC_11_15_1  (
            .in0(N__27698),
            .in1(N__32832),
            .in2(N__27920),
            .in3(N__32670),
            .lcout(\POWERLED.dutycycle_RNI36306Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI24KO1_15_LC_11_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI24KO1_15_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI24KO1_15_LC_11_15_2 .LUT_INIT=16'b1000000010101010;
    LogicCell40 \POWERLED.dutycycle_RNI24KO1_15_LC_11_15_2  (
            .in0(N__27897),
            .in1(N__33127),
            .in2(N__27476),
            .in3(N__27831),
            .lcout(\POWERLED.N_529 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIE3861_14_LC_11_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIE3861_14_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIE3861_14_LC_11_15_3 .LUT_INIT=16'b1000000010101010;
    LogicCell40 \POWERLED.dutycycle_RNIE3861_14_LC_11_15_3  (
            .in0(N__30227),
            .in1(N__29757),
            .in2(N__27687),
            .in3(N__27769),
            .lcout(),
            .ltout(\POWERLED.N_524_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNID4I22_14_LC_11_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNID4I22_14_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNID4I22_14_LC_11_15_4 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \POWERLED.dutycycle_RNID4I22_14_LC_11_15_4  (
            .in0(N__27768),
            .in1(N__27459),
            .in2(N__27701),
            .in3(N__30150),
            .lcout(\POWERLED.un1_clk_100khz_47_and_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIE3861_15_LC_11_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIE3861_15_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIE3861_15_LC_11_15_5 .LUT_INIT=16'b1000000010101010;
    LogicCell40 \POWERLED.dutycycle_RNIE3861_15_LC_11_15_5  (
            .in0(N__30228),
            .in1(N__29758),
            .in2(N__27688),
            .in3(N__27520),
            .lcout(),
            .ltout(\POWERLED.N_527_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNID4I22_1_LC_11_15_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNID4I22_1_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNID4I22_1_LC_11_15_6 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \POWERLED.func_state_RNID4I22_1_LC_11_15_6  (
            .in0(N__27475),
            .in1(N__27460),
            .in2(N__27383),
            .in3(N__30151),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_48_and_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI36306_1_LC_11_15_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI36306_1_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI36306_1_LC_11_15_7 .LUT_INIT=16'b0010001000101010;
    LogicCell40 \POWERLED.func_state_RNI36306_1_LC_11_15_7  (
            .in0(N__32671),
            .in1(N__32833),
            .in2(N__27380),
            .in3(N__27968),
            .lcout(\POWERLED.dutycycle_en_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI300O2_8_LC_12_3_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI300O2_8_LC_12_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI300O2_8_LC_12_3_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNI300O2_8_LC_12_3_0  (
            .in0(N__29080),
            .in1(N__27950),
            .in2(_gnd_net_),
            .in3(N__28228),
            .lcout(\POWERLED.count_clkZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_8_LC_12_3_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_8_LC_12_3_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_8_LC_12_3_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_8_LC_12_3_1  (
            .in0(N__28229),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32261),
            .ce(N__29106),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_15_LC_12_3_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_15_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_15_LC_12_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_15_LC_12_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28463),
            .lcout(\POWERLED.count_clk_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32261),
            .ce(N__29106),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI531O2_9_LC_12_3_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI531O2_9_LC_12_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI531O2_9_LC_12_3_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNI531O2_9_LC_12_3_4  (
            .in0(N__29081),
            .in1(N__27944),
            .in2(_gnd_net_),
            .in3(N__28189),
            .lcout(\POWERLED.count_clkZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_9_LC_12_3_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_9_LC_12_3_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_9_LC_12_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_9_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28190),
            .lcout(\POWERLED.count_clk_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32261),
            .ce(N__29106),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNINDPN2_2_LC_12_3_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNINDPN2_2_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNINDPN2_2_LC_12_3_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \POWERLED.count_clk_RNINDPN2_2_LC_12_3_6  (
            .in0(_gnd_net_),
            .in1(N__27938),
            .in2(N__29104),
            .in3(N__28027),
            .lcout(\POWERLED.count_clkZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_2_LC_12_3_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_2_LC_12_3_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_2_LC_12_3_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_2_LC_12_3_7  (
            .in0(N__28028),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32261),
            .ce(N__29106),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_3_LC_12_4_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_3_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_3_LC_12_4_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_3_LC_12_4_0  (
            .in0(N__28004),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32309),
            .ce(N__29076),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIPGQN2_3_LC_12_4_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIPGQN2_3_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIPGQN2_3_LC_12_4_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNIPGQN2_3_LC_12_4_1  (
            .in0(N__28147),
            .in1(N__29082),
            .in2(_gnd_net_),
            .in3(N__28002),
            .lcout(\POWERLED.count_clkZ0Z_3 ),
            .ltout(\POWERLED.count_clkZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_3_LC_12_4_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_3_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_3_LC_12_4_2 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \POWERLED.count_clk_RNI_3_LC_12_4_2  (
            .in0(N__28044),
            .in1(N__27987),
            .in2(N__28154),
            .in3(N__28245),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_168_0_0_o2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_6_LC_12_4_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_6_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_6_LC_12_4_3 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \POWERLED.count_clk_RNI_6_LC_12_4_3  (
            .in0(N__28345),
            .in1(N__28314),
            .in2(N__28151),
            .in3(N__28110),
            .lcout(\POWERLED.count_clk_RNIZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIPGQN2_0_3_LC_12_4_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIPGQN2_0_3_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIPGQN2_0_3_LC_12_4_4 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \POWERLED.count_clk_RNIPGQN2_0_3_LC_12_4_4  (
            .in0(N__28003),
            .in1(N__28148),
            .in2(N__29105),
            .in3(N__28246),
            .lcout(),
            .ltout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIPGQN2_1_3_LC_12_4_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIPGQN2_1_3_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIPGQN2_1_3_LC_12_4_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.count_clk_RNIPGQN2_1_3_LC_12_4_5  (
            .in0(N__28346),
            .in1(N__27988),
            .in2(N__28136),
            .in3(N__28045),
            .lcout(\POWERLED.N_625 ),
            .ltout(\POWERLED.N_625_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIPGQN2_5_3_LC_12_4_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIPGQN2_5_3_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIPGQN2_5_3_LC_12_4_6 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \POWERLED.count_clk_RNIPGQN2_5_3_LC_12_4_6  (
            .in0(N__28111),
            .in1(_gnd_net_),
            .in2(N__28091),
            .in3(N__28319),
            .lcout(\POWERLED.count_clk_RNIPGQN2_5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_12_5_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_12_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(N__28721),
            .in2(N__28075),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_5_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_12_5_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_12_5_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_12_5_1  (
            .in0(N__28547),
            .in1(_gnd_net_),
            .in2(N__28049),
            .in3(N__28016),
            .lcout(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_1 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_12_5_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_12_5_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_12_5_2  (
            .in0(N__28551),
            .in1(_gnd_net_),
            .in2(N__28013),
            .in3(N__27992),
            .lcout(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_2 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_12_5_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_12_5_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_12_5_3  (
            .in0(N__28548),
            .in1(_gnd_net_),
            .in2(N__27989),
            .in3(N__28385),
            .lcout(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_3 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_12_5_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_12_5_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_12_5_4  (
            .in0(N__28552),
            .in1(_gnd_net_),
            .in2(N__28381),
            .in3(N__28349),
            .lcout(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_4 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_12_5_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_12_5_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_12_5_5  (
            .in0(N__28549),
            .in1(N__28344),
            .in2(_gnd_net_),
            .in3(N__28322),
            .lcout(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_5 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_12_5_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_12_5_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_12_5_6  (
            .in0(N__28553),
            .in1(_gnd_net_),
            .in2(N__28318),
            .in3(N__28250),
            .lcout(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_6 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_12_5_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_12_5_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_12_5_7  (
            .in0(N__28550),
            .in1(N__28247),
            .in2(_gnd_net_),
            .in3(N__28217),
            .lcout(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_7 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_12_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_12_6_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_12_6_0  (
            .in0(N__28540),
            .in1(N__28213),
            .in2(_gnd_net_),
            .in3(N__28175),
            .lcout(\POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_12_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_12_6_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_12_6_1  (
            .in0(N__28543),
            .in1(N__28406),
            .in2(_gnd_net_),
            .in3(N__28172),
            .lcout(\POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_9 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_12_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_12_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(N__28672),
            .in2(_gnd_net_),
            .in3(N__28160),
            .lcout(\POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_10 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_11_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_12_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_12_6_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_12_6_3  (
            .in0(N__28544),
            .in1(_gnd_net_),
            .in2(N__28571),
            .in3(N__28157),
            .lcout(\POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_11_cZ0 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_12_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_12_6_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_12_6_4  (
            .in0(N__28541),
            .in1(N__29144),
            .in2(_gnd_net_),
            .in3(N__28559),
            .lcout(\POWERLED.count_clk_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_12 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_13_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNITQ5G2_LC_12_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNITQ5G2_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNITQ5G2_LC_12_6_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_13_c_RNITQ5G2_LC_12_6_5  (
            .in0(N__28545),
            .in1(N__28400),
            .in2(_gnd_net_),
            .in3(N__28556),
            .lcout(\POWERLED.count_clk_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_13_cZ0 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_12_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_12_6_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_12_6_6  (
            .in0(N__28542),
            .in1(N__28448),
            .in2(_gnd_net_),
            .in3(N__28475),
            .lcout(\POWERLED.count_clk_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIVT6G2_15_LC_12_6_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIVT6G2_15_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIVT6G2_15_LC_12_6_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNIVT6G2_15_LC_12_6_7  (
            .in0(N__29075),
            .in1(N__28472),
            .in2(_gnd_net_),
            .in3(N__28459),
            .lcout(\POWERLED.count_clkZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIECHG2_10_LC_12_7_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIECHG2_10_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIECHG2_10_LC_12_7_0 .LUT_INIT=16'b1111111110101100;
    LogicCell40 \POWERLED.count_clk_RNIECHG2_10_LC_12_7_0  (
            .in0(N__28436),
            .in1(N__28414),
            .in2(N__29119),
            .in3(N__28447),
            .lcout(\POWERLED.un2_count_clk_17_0_o2_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_10_LC_12_7_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_10_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_10_LC_12_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_10_LC_12_7_1  (
            .in0(N__28429),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clkZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32380),
            .ce(N__29110),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIECHG2_0_10_LC_12_7_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIECHG2_0_10_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIECHG2_0_10_LC_12_7_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \POWERLED.count_clk_RNIECHG2_0_10_LC_12_7_2  (
            .in0(N__28991),
            .in1(N__28428),
            .in2(_gnd_net_),
            .in3(N__28415),
            .lcout(\POWERLED.un1_count_clk_2_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_14_LC_12_7_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_14_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_14_LC_12_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_14_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28695),
            .lcout(\POWERLED.count_clkZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32380),
            .ce(N__29110),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNILKND2_0_14_LC_12_7_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNILKND2_0_14_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNILKND2_0_14_LC_12_7_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \POWERLED.count_clk_RNILKND2_0_14_LC_12_7_4  (
            .in0(N__28696),
            .in1(_gnd_net_),
            .in2(N__29120),
            .in3(N__28681),
            .lcout(\POWERLED.un1_count_clk_2_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI008L2_0_LC_12_7_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI008L2_0_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI008L2_0_LC_12_7_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_clk_RNI008L2_0_LC_12_7_5  (
            .in0(N__28733),
            .in1(N__28990),
            .in2(_gnd_net_),
            .in3(N__28727),
            .lcout(\POWERLED.count_clkZ0Z_0 ),
            .ltout(\POWERLED.count_clkZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNILKND2_14_LC_12_7_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNILKND2_14_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNILKND2_14_LC_12_7_6 .LUT_INIT=16'b1111101111111000;
    LogicCell40 \POWERLED.count_clk_RNILKND2_14_LC_12_7_6  (
            .in0(N__28697),
            .in1(N__29074),
            .in2(N__28685),
            .in3(N__28682),
            .lcout(),
            .ltout(\POWERLED.un2_count_clk_17_0_o2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNISLCE7_10_LC_12_7_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNISLCE7_10_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNISLCE7_10_LC_12_7_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNISLCE7_10_LC_12_7_7  (
            .in0(N__28673),
            .in1(N__28931),
            .in2(N__28661),
            .in3(N__28658),
            .lcout(\POWERLED.count_clk_RNISLCE7Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5SKJ1_0_1_LC_12_8_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5SKJ1_0_1_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5SKJ1_0_1_LC_12_8_0 .LUT_INIT=16'b0000000011101100;
    LogicCell40 \POWERLED.func_state_RNI5SKJ1_0_1_LC_12_8_0  (
            .in0(N__30740),
            .in1(N__29608),
            .in2(N__28637),
            .in3(N__28892),
            .lcout(),
            .ltout(\POWERLED.count_clk_en_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI6GV92_1_LC_12_8_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI6GV92_1_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI6GV92_1_LC_12_8_1 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \POWERLED.func_state_RNI6GV92_1_LC_12_8_1  (
            .in0(N__28623),
            .in1(N__32644),
            .in2(N__28601),
            .in3(N__28598),
            .lcout(\POWERLED.count_clk_en ),
            .ltout(\POWERLED.count_clk_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIPK3G2_0_12_LC_12_8_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIPK3G2_0_12_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIPK3G2_0_12_LC_12_8_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \POWERLED.count_clk_RNIPK3G2_0_12_LC_12_8_2  (
            .in0(N__29134),
            .in1(_gnd_net_),
            .in2(N__28574),
            .in3(N__28939),
            .lcout(\POWERLED.un1_count_clk_2_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_12_LC_12_8_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_12_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_12_LC_12_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_12_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29133),
            .lcout(\POWERLED.count_clkZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32407),
            .ce(N__29069),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_13_LC_12_8_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_13_LC_12_8_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_13_LC_12_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_13_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29161),
            .lcout(\POWERLED.count_clk_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32407),
            .ce(N__29069),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIRN4G2_13_LC_12_8_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIRN4G2_13_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIRN4G2_13_LC_12_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_clk_RNIRN4G2_13_LC_12_8_5  (
            .in0(N__29162),
            .in1(N__29150),
            .in2(_gnd_net_),
            .in3(N__29070),
            .lcout(\POWERLED.count_clkZ0Z_13 ),
            .ltout(\POWERLED.count_clkZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIPK3G2_12_LC_12_8_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIPK3G2_12_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIPK3G2_12_LC_12_8_6 .LUT_INIT=16'b1111101111111000;
    LogicCell40 \POWERLED.count_clk_RNIPK3G2_12_LC_12_8_6  (
            .in0(N__29135),
            .in1(N__29037),
            .in2(N__28943),
            .in3(N__28940),
            .lcout(\POWERLED.un2_count_clk_17_0_o2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_4_0_LC_12_8_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_4_0_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_4_0_LC_12_8_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.func_state_RNI_4_0_LC_12_8_7  (
            .in0(N__31588),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28908),
            .lcout(\POWERLED.N_492 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_5_LC_12_9_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_5_LC_12_9_1 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_5_LC_12_9_1 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \POWERLED.dutycycle_5_LC_12_9_1  (
            .in0(N__28874),
            .in1(N__28885),
            .in2(N__32836),
            .in3(N__30434),
            .lcout(\POWERLED.dutycycle_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32465),
            .ce(),
            .sr(N__31756));
    defparam \POWERLED.dutycycle_RNIKVDEF_5_LC_12_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKVDEF_5_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKVDEF_5_LC_12_9_2 .LUT_INIT=16'b0111011111110000;
    LogicCell40 \POWERLED.dutycycle_RNIKVDEF_5_LC_12_9_2  (
            .in0(N__30433),
            .in1(N__32821),
            .in2(N__28886),
            .in3(N__28873),
            .lcout(\POWERLED.dutycycleZ1Z_5 ),
            .ltout(\POWERLED.dutycycleZ1Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_5_LC_12_9_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_5_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_5_LC_12_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_5_LC_12_9_3  (
            .in0(N__29369),
            .in1(N__31105),
            .in2(N__28859),
            .in3(N__28845),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_5 ),
            .ltout(\POWERLED.dutycycle_RNI_3Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_5_LC_12_9_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_5_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_5_LC_12_9_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_5_LC_12_9_4  (
            .in0(N__30785),
            .in1(_gnd_net_),
            .in2(N__28856),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.dutycycle_0_sqmuxa_i_i_a3_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_5_LC_12_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_5_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_5_LC_12_9_5 .LUT_INIT=16'b1100111011011111;
    LogicCell40 \POWERLED.dutycycle_RNI_8_5_LC_12_9_5  (
            .in0(N__29173),
            .in1(N__31591),
            .in2(N__28853),
            .in3(N__28846),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_8Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOGRS_1_LC_12_9_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOGRS_1_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOGRS_1_LC_12_9_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \POWERLED.func_state_RNIOGRS_1_LC_12_9_6  (
            .in0(N__28739),
            .in1(N__30835),
            .in2(N__29762),
            .in3(N__29293),
            .lcout(),
            .ltout(\POWERLED.func_state_RNIOGRSZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNITCGG2_1_LC_12_9_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNITCGG2_1_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNITCGG2_1_LC_12_9_7 .LUT_INIT=16'b0000111111101110;
    LogicCell40 \POWERLED.func_state_RNITCGG2_1_LC_12_9_7  (
            .in0(N__29725),
            .in1(N__29669),
            .in2(N__29633),
            .in3(N__29600),
            .lcout(\POWERLED.N_413_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_6_LC_12_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_6_LC_12_10_0 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_6_LC_12_10_0 .LUT_INIT=16'b0101110011111100;
    LogicCell40 \POWERLED.dutycycle_6_LC_12_10_0  (
            .in0(N__30812),
            .in1(N__29470),
            .in2(N__32492),
            .in3(N__32815),
            .lcout(\POWERLED.dutycycle_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32461),
            .ce(),
            .sr(N__31755));
    defparam \POWERLED.dutycycle_RNIQCMNB_6_LC_12_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQCMNB_6_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQCMNB_6_LC_12_10_1 .LUT_INIT=16'b0111011111110000;
    LogicCell40 \POWERLED.dutycycle_RNIQCMNB_6_LC_12_10_1  (
            .in0(N__32814),
            .in1(N__30811),
            .in2(N__29471),
            .in3(N__32488),
            .lcout(\POWERLED.dutycycleZ0Z_6 ),
            .ltout(\POWERLED.dutycycleZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_6_LC_12_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_6_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_6_LC_12_10_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_6_LC_12_10_2  (
            .in0(N__29364),
            .in1(_gnd_net_),
            .in2(N__29459),
            .in3(N__29455),
            .lcout(\POWERLED.N_672 ),
            .ltout(\POWERLED.N_672_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_6_LC_12_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_6_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_6_LC_12_10_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \POWERLED.dutycycle_RNI_5_6_LC_12_10_3  (
            .in0(N__29389),
            .in1(_gnd_net_),
            .in2(N__29411),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_dutycycle_168_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_1_6_LC_12_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_1_6_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_1_6_LC_12_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.count_clk_RNI_1_6_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29388),
            .lcout(\POWERLED.N_412_i ),
            .ltout(\POWERLED.N_412_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_3_LC_12_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_12_10_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_3_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(N__29365),
            .in2(N__29339),
            .in3(N__29336),
            .lcout(\POWERLED.dutycycle_RNI_6Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_5_1_LC_12_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_5_1_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_5_1_LC_12_10_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \POWERLED.func_state_RNI_5_1_LC_12_10_6  (
            .in0(N__29291),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29209),
            .lcout(\POWERLED.func_state_RNI_5Z0Z_1 ),
            .ltout(\POWERLED.func_state_RNI_5Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_9_1_LC_12_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_9_1_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_9_1_LC_12_10_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.func_state_RNI_9_1_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30842),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_23_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIJM2T1_LC_12_11_0 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIJM2T1_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIJM2T1_LC_12_11_0 .LUT_INIT=16'b1111111110100011;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNIJM2T1_LC_12_11_0  (
            .in0(N__30469),
            .in1(N__30824),
            .in2(N__30316),
            .in3(N__30442),
            .lcout(\POWERLED.N_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI12AS_1_LC_12_11_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI12AS_1_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI12AS_1_LC_12_11_1 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \POWERLED.func_state_RNI12AS_1_LC_12_11_1  (
            .in0(N__30598),
            .in1(N__29896),
            .in2(_gnd_net_),
            .in3(N__30124),
            .lcout(\POWERLED.func_state_RNI12ASZ0Z_1 ),
            .ltout(\POWERLED.func_state_RNI12ASZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI12AS_5_LC_12_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI12AS_5_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI12AS_5_LC_12_11_2 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \POWERLED.dutycycle_RNI12AS_5_LC_12_11_2  (
            .in0(N__30803),
            .in1(_gnd_net_),
            .in2(N__30788),
            .in3(N__30769),
            .lcout(\POWERLED.dutycycle_eena_13_c_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI12AS_6_LC_12_11_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI12AS_6_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI12AS_6_LC_12_11_3 .LUT_INIT=16'b0100010101010101;
    LogicCell40 \POWERLED.dutycycle_RNI12AS_6_LC_12_11_3  (
            .in0(N__31088),
            .in1(N__30125),
            .in2(N__30664),
            .in3(N__29895),
            .lcout(\POWERLED.N_530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIIK1T1_LC_12_11_4 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIIK1T1_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIIK1T1_LC_12_11_4 .LUT_INIT=16'b1111111110100011;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNIIK1T1_LC_12_11_4  (
            .in0(N__30470),
            .in1(N__30455),
            .in2(N__30315),
            .in3(N__30443),
            .lcout(\POWERLED.N_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI01AS_6_LC_12_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI01AS_6_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI01AS_6_LC_12_11_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.dutycycle_RNI01AS_6_LC_12_11_5  (
            .in0(N__31087),
            .in1(N__30289),
            .in2(N__30148),
            .in3(N__29897),
            .lcout(),
            .ltout(\POWERLED.N_532_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIBD845_6_LC_12_11_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIBD845_6_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIBD845_6_LC_12_11_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.dutycycle_RNIBD845_6_LC_12_11_6  (
            .in0(N__29813),
            .in1(N__29789),
            .in2(N__29771),
            .in3(N__29768),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_51_and_i_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI0DF58_5_LC_12_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI0DF58_5_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI0DF58_5_LC_12_11_7 .LUT_INIT=16'b0011101100000000;
    LogicCell40 \POWERLED.dutycycle_RNI0DF58_5_LC_12_11_7  (
            .in0(N__32849),
            .in1(N__32825),
            .in2(N__32678),
            .in3(N__32637),
            .lcout(\POWERLED.dutycycle_RNI0DF58Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_3_LC_12_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_3_LC_12_12_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_3_LC_12_12_0 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \POWERLED.dutycycle_3_LC_12_12_0  (
            .in0(N__31498),
            .in1(N__31603),
            .in2(N__31637),
            .in3(N__31622),
            .lcout(\POWERLED.dutycycleZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32464),
            .ce(),
            .sr(N__31773));
    defparam \POWERLED.dutycycle_RNIH92L6_3_LC_12_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIH92L6_3_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIH92L6_3_LC_12_12_1 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \POWERLED.dutycycle_RNIH92L6_3_LC_12_12_1  (
            .in0(N__31633),
            .in1(N__31621),
            .in2(N__31604),
            .in3(N__31497),
            .lcout(\POWERLED.dutycycleZ0Z_8 ),
            .ltout(\POWERLED.dutycycleZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_2_LC_12_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_12_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_2_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__31103),
            .in2(N__31442),
            .in3(N__32944),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_5_LC_12_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_5_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_5_LC_12_12_3 .LUT_INIT=16'b0001111011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_5_LC_12_12_3  (
            .in0(N__31263),
            .in1(N__31426),
            .in2(N__31439),
            .in3(N__30917),
            .lcout(\POWERLED.un1_dutycycle_53_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_3_LC_12_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_12_12_5 .LUT_INIT=16'b0000011000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_3_LC_12_12_5  (
            .in0(N__31104),
            .in1(N__30982),
            .in2(N__31436),
            .in3(N__30918),
            .lcout(),
            .ltout(\POWERLED.un1_i3_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_5_LC_12_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_5_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_5_LC_12_12_6 .LUT_INIT=16'b1010001110100011;
    LogicCell40 \POWERLED.dutycycle_RNI_1_5_LC_12_12_6  (
            .in0(N__31264),
            .in1(N__30848),
            .in2(N__31190),
            .in3(N__31187),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_3_LC_12_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_12_12_7 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_3_LC_12_12_7  (
            .in0(N__31102),
            .in1(N__30981),
            .in2(_gnd_net_),
            .in3(N__30916),
            .lcout(\POWERLED.d_i3_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNISQ2V_LC_12_13_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNISQ2V_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNISQ2V_LC_12_13_1 .LUT_INIT=16'b1011101110111011;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNISQ2V_LC_12_13_1  (
            .in0(N__33161),
            .in1(N__33123),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vpp_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_LC_12_13_5 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_LC_12_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_LC_12_13_5  (
            .in0(N__33020),
            .in1(N__33002),
            .in2(N__32987),
            .in3(N__32975),
            .lcout(vccin_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_2_LC_12_13_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_2_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_2_LC_12_13_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_2_2_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__32948),
            .in2(_gnd_net_),
            .in3(N__32864),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TOP
