// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Aug 16 2022 15:17:42

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VR_READY_VCCINAUX,
    V33A_ENn,
    V1P8A_EN,
    VDDQ_EN,
    VCCST_OVERRIDE_3V3,
    V5S_OK,
    SLP_S3n,
    SLP_S0n,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    GPIO_FPGA_SoC_2,
    VCCIN_VR_PROCHOT_FPGA,
    SLP_SUSn,
    CPU_C10_GATE_N,
    VCCST_EN,
    V33DSW_OK,
    TPM_GPIO,
    SUSWARN_N,
    PLTRSTn,
    GPIO_FPGA_SoC_4,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    FPGA_OSC,
    VCCST_PWRGD,
    SYS_PWROK,
    SPI_FP_IO2,
    SATAXPCIE1_FPGA,
    GPIO_FPGA_EXP_1,
    VCCINAUX_VR_PROCHOT_FPGA,
    VCCINAUX_VR_PE,
    HDA_SDO_ATP,
    GPIO_FPGA_EXP_2,
    VPP_EN,
    VDDQ_OK,
    SUSACK_N,
    SLP_S4n,
    VCCST_CPU_OK,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    GPIO_FPGA_SoC_1,
    DSW_PWROK,
    V5A_EN,
    GPIO_FPGA_SoC_3,
    VR_PROCHOT_FPGA_OUT_N,
    VPP_OK,
    VCCIN_VR_PE,
    VCCIN_EN,
    SOC_SPKR,
    SLP_S5n,
    V12_MAIN_MON,
    SPI_FP_IO3,
    SATAXPCIE0_FPGA,
    V33A_OK,
    PCH_PWROK,
    FPGA_SLP_WLAN_N);

    input VR_READY_VCCINAUX;
    output V33A_ENn;
    output V1P8A_EN;
    output VDDQ_EN;
    input VCCST_OVERRIDE_3V3;
    input V5S_OK;
    input SLP_S3n;
    input SLP_S0n;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input GPIO_FPGA_SoC_2;
    input VCCIN_VR_PROCHOT_FPGA;
    input SLP_SUSn;
    input CPU_C10_GATE_N;
    output VCCST_EN;
    input V33DSW_OK;
    input TPM_GPIO;
    output SUSWARN_N;
    input PLTRSTn;
    input GPIO_FPGA_SoC_4;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output SYS_PWROK;
    input SPI_FP_IO2;
    input SATAXPCIE1_FPGA;
    input GPIO_FPGA_EXP_1;
    input VCCINAUX_VR_PROCHOT_FPGA;
    output VCCINAUX_VR_PE;
    output HDA_SDO_ATP;
    input GPIO_FPGA_EXP_2;
    output VPP_EN;
    input VDDQ_OK;
    input SUSACK_N;
    input SLP_S4n;
    input VCCST_CPU_OK;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input GPIO_FPGA_SoC_1;
    output DSW_PWROK;
    output V5A_EN;
    input GPIO_FPGA_SoC_3;
    input VR_PROCHOT_FPGA_OUT_N;
    input VPP_OK;
    output VCCIN_VR_PE;
    output VCCIN_EN;
    input SOC_SPKR;
    input SLP_S5n;
    input V12_MAIN_MON;
    input SPI_FP_IO3;
    input SATAXPCIE0_FPGA;
    input V33A_OK;
    output PCH_PWROK;
    input FPGA_SLP_WLAN_N;

    wire N__19975;
    wire N__19974;
    wire N__19973;
    wire N__19966;
    wire N__19965;
    wire N__19964;
    wire N__19957;
    wire N__19956;
    wire N__19955;
    wire N__19948;
    wire N__19947;
    wire N__19946;
    wire N__19939;
    wire N__19938;
    wire N__19937;
    wire N__19930;
    wire N__19929;
    wire N__19928;
    wire N__19921;
    wire N__19920;
    wire N__19919;
    wire N__19912;
    wire N__19911;
    wire N__19910;
    wire N__19903;
    wire N__19902;
    wire N__19901;
    wire N__19894;
    wire N__19893;
    wire N__19892;
    wire N__19885;
    wire N__19884;
    wire N__19883;
    wire N__19876;
    wire N__19875;
    wire N__19874;
    wire N__19867;
    wire N__19866;
    wire N__19865;
    wire N__19858;
    wire N__19857;
    wire N__19856;
    wire N__19849;
    wire N__19848;
    wire N__19847;
    wire N__19840;
    wire N__19839;
    wire N__19838;
    wire N__19831;
    wire N__19830;
    wire N__19829;
    wire N__19822;
    wire N__19821;
    wire N__19820;
    wire N__19813;
    wire N__19812;
    wire N__19811;
    wire N__19804;
    wire N__19803;
    wire N__19802;
    wire N__19795;
    wire N__19794;
    wire N__19793;
    wire N__19786;
    wire N__19785;
    wire N__19784;
    wire N__19777;
    wire N__19776;
    wire N__19775;
    wire N__19768;
    wire N__19767;
    wire N__19766;
    wire N__19759;
    wire N__19758;
    wire N__19757;
    wire N__19750;
    wire N__19749;
    wire N__19748;
    wire N__19741;
    wire N__19740;
    wire N__19739;
    wire N__19732;
    wire N__19731;
    wire N__19730;
    wire N__19723;
    wire N__19722;
    wire N__19721;
    wire N__19714;
    wire N__19713;
    wire N__19712;
    wire N__19705;
    wire N__19704;
    wire N__19703;
    wire N__19696;
    wire N__19695;
    wire N__19694;
    wire N__19687;
    wire N__19686;
    wire N__19685;
    wire N__19678;
    wire N__19677;
    wire N__19676;
    wire N__19669;
    wire N__19668;
    wire N__19667;
    wire N__19660;
    wire N__19659;
    wire N__19658;
    wire N__19651;
    wire N__19650;
    wire N__19649;
    wire N__19642;
    wire N__19641;
    wire N__19640;
    wire N__19633;
    wire N__19632;
    wire N__19631;
    wire N__19624;
    wire N__19623;
    wire N__19622;
    wire N__19615;
    wire N__19614;
    wire N__19613;
    wire N__19606;
    wire N__19605;
    wire N__19604;
    wire N__19597;
    wire N__19596;
    wire N__19595;
    wire N__19588;
    wire N__19587;
    wire N__19586;
    wire N__19579;
    wire N__19578;
    wire N__19577;
    wire N__19570;
    wire N__19569;
    wire N__19568;
    wire N__19561;
    wire N__19560;
    wire N__19559;
    wire N__19552;
    wire N__19551;
    wire N__19550;
    wire N__19543;
    wire N__19542;
    wire N__19541;
    wire N__19534;
    wire N__19533;
    wire N__19532;
    wire N__19525;
    wire N__19524;
    wire N__19523;
    wire N__19516;
    wire N__19515;
    wire N__19514;
    wire N__19507;
    wire N__19506;
    wire N__19505;
    wire N__19498;
    wire N__19497;
    wire N__19496;
    wire N__19489;
    wire N__19488;
    wire N__19487;
    wire N__19480;
    wire N__19479;
    wire N__19478;
    wire N__19471;
    wire N__19470;
    wire N__19469;
    wire N__19462;
    wire N__19461;
    wire N__19460;
    wire N__19453;
    wire N__19452;
    wire N__19451;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19427;
    wire N__19424;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19397;
    wire N__19394;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19374;
    wire N__19371;
    wire N__19370;
    wire N__19369;
    wire N__19368;
    wire N__19367;
    wire N__19366;
    wire N__19365;
    wire N__19364;
    wire N__19363;
    wire N__19362;
    wire N__19361;
    wire N__19360;
    wire N__19359;
    wire N__19358;
    wire N__19357;
    wire N__19356;
    wire N__19353;
    wire N__19344;
    wire N__19337;
    wire N__19330;
    wire N__19319;
    wire N__19316;
    wire N__19309;
    wire N__19302;
    wire N__19299;
    wire N__19298;
    wire N__19297;
    wire N__19296;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19271;
    wire N__19268;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19258;
    wire N__19255;
    wire N__19248;
    wire N__19245;
    wire N__19244;
    wire N__19243;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19232;
    wire N__19231;
    wire N__19230;
    wire N__19229;
    wire N__19226;
    wire N__19225;
    wire N__19224;
    wire N__19223;
    wire N__19222;
    wire N__19215;
    wire N__19214;
    wire N__19213;
    wire N__19212;
    wire N__19211;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19201;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19185;
    wire N__19182;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19174;
    wire N__19171;
    wire N__19170;
    wire N__19167;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19159;
    wire N__19156;
    wire N__19155;
    wire N__19154;
    wire N__19151;
    wire N__19146;
    wire N__19139;
    wire N__19138;
    wire N__19137;
    wire N__19134;
    wire N__19131;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19119;
    wire N__19116;
    wire N__19115;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19097;
    wire N__19094;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19086;
    wire N__19085;
    wire N__19082;
    wire N__19081;
    wire N__19074;
    wire N__19071;
    wire N__19068;
    wire N__19067;
    wire N__19066;
    wire N__19061;
    wire N__19058;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19042;
    wire N__19037;
    wire N__19032;
    wire N__19027;
    wire N__19024;
    wire N__19023;
    wire N__19022;
    wire N__19017;
    wire N__19014;
    wire N__19013;
    wire N__19012;
    wire N__19009;
    wire N__19008;
    wire N__19005;
    wire N__19002;
    wire N__19001;
    wire N__18996;
    wire N__18993;
    wire N__18990;
    wire N__18987;
    wire N__18982;
    wire N__18975;
    wire N__18972;
    wire N__18969;
    wire N__18962;
    wire N__18959;
    wire N__18958;
    wire N__18955;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18937;
    wire N__18932;
    wire N__18929;
    wire N__18920;
    wire N__18913;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18895;
    wire N__18894;
    wire N__18891;
    wire N__18886;
    wire N__18883;
    wire N__18878;
    wire N__18873;
    wire N__18868;
    wire N__18863;
    wire N__18860;
    wire N__18851;
    wire N__18840;
    wire N__18839;
    wire N__18838;
    wire N__18837;
    wire N__18836;
    wire N__18835;
    wire N__18834;
    wire N__18833;
    wire N__18832;
    wire N__18831;
    wire N__18830;
    wire N__18829;
    wire N__18828;
    wire N__18827;
    wire N__18826;
    wire N__18825;
    wire N__18824;
    wire N__18823;
    wire N__18822;
    wire N__18821;
    wire N__18820;
    wire N__18819;
    wire N__18818;
    wire N__18817;
    wire N__18816;
    wire N__18815;
    wire N__18814;
    wire N__18813;
    wire N__18812;
    wire N__18811;
    wire N__18810;
    wire N__18809;
    wire N__18808;
    wire N__18807;
    wire N__18806;
    wire N__18805;
    wire N__18804;
    wire N__18803;
    wire N__18802;
    wire N__18801;
    wire N__18800;
    wire N__18799;
    wire N__18798;
    wire N__18797;
    wire N__18796;
    wire N__18795;
    wire N__18794;
    wire N__18793;
    wire N__18792;
    wire N__18791;
    wire N__18790;
    wire N__18789;
    wire N__18788;
    wire N__18787;
    wire N__18786;
    wire N__18785;
    wire N__18784;
    wire N__18783;
    wire N__18782;
    wire N__18781;
    wire N__18780;
    wire N__18779;
    wire N__18778;
    wire N__18777;
    wire N__18776;
    wire N__18775;
    wire N__18774;
    wire N__18773;
    wire N__18772;
    wire N__18771;
    wire N__18770;
    wire N__18769;
    wire N__18768;
    wire N__18767;
    wire N__18766;
    wire N__18765;
    wire N__18764;
    wire N__18763;
    wire N__18762;
    wire N__18761;
    wire N__18760;
    wire N__18759;
    wire N__18758;
    wire N__18757;
    wire N__18756;
    wire N__18755;
    wire N__18754;
    wire N__18753;
    wire N__18752;
    wire N__18751;
    wire N__18750;
    wire N__18749;
    wire N__18748;
    wire N__18747;
    wire N__18746;
    wire N__18745;
    wire N__18744;
    wire N__18743;
    wire N__18742;
    wire N__18741;
    wire N__18740;
    wire N__18739;
    wire N__18738;
    wire N__18737;
    wire N__18728;
    wire N__18719;
    wire N__18710;
    wire N__18701;
    wire N__18692;
    wire N__18683;
    wire N__18674;
    wire N__18667;
    wire N__18658;
    wire N__18651;
    wire N__18642;
    wire N__18635;
    wire N__18626;
    wire N__18619;
    wire N__18610;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18585;
    wire N__18578;
    wire N__18569;
    wire N__18562;
    wire N__18559;
    wire N__18550;
    wire N__18543;
    wire N__18538;
    wire N__18529;
    wire N__18520;
    wire N__18517;
    wire N__18510;
    wire N__18507;
    wire N__18504;
    wire N__18501;
    wire N__18498;
    wire N__18495;
    wire N__18492;
    wire N__18491;
    wire N__18490;
    wire N__18489;
    wire N__18488;
    wire N__18487;
    wire N__18486;
    wire N__18485;
    wire N__18482;
    wire N__18481;
    wire N__18478;
    wire N__18477;
    wire N__18476;
    wire N__18475;
    wire N__18474;
    wire N__18473;
    wire N__18472;
    wire N__18469;
    wire N__18468;
    wire N__18465;
    wire N__18462;
    wire N__18459;
    wire N__18456;
    wire N__18453;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18409;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18397;
    wire N__18394;
    wire N__18391;
    wire N__18388;
    wire N__18385;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18373;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18255;
    wire N__18252;
    wire N__18249;
    wire N__18246;
    wire N__18243;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18231;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18219;
    wire N__18218;
    wire N__18215;
    wire N__18212;
    wire N__18207;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18192;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18180;
    wire N__18177;
    wire N__18174;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18162;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18150;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18135;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18093;
    wire N__18090;
    wire N__18087;
    wire N__18084;
    wire N__18081;
    wire N__18078;
    wire N__18075;
    wire N__18072;
    wire N__18071;
    wire N__18070;
    wire N__18069;
    wire N__18066;
    wire N__18061;
    wire N__18058;
    wire N__18055;
    wire N__18052;
    wire N__18049;
    wire N__18042;
    wire N__18039;
    wire N__18036;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18024;
    wire N__18023;
    wire N__18020;
    wire N__18019;
    wire N__18016;
    wire N__18015;
    wire N__18012;
    wire N__18009;
    wire N__18006;
    wire N__18003;
    wire N__17994;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17982;
    wire N__17981;
    wire N__17978;
    wire N__17975;
    wire N__17970;
    wire N__17969;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17955;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17943;
    wire N__17940;
    wire N__17937;
    wire N__17934;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17926;
    wire N__17925;
    wire N__17922;
    wire N__17919;
    wire N__17916;
    wire N__17913;
    wire N__17910;
    wire N__17905;
    wire N__17902;
    wire N__17895;
    wire N__17892;
    wire N__17889;
    wire N__17886;
    wire N__17883;
    wire N__17880;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17868;
    wire N__17865;
    wire N__17862;
    wire N__17861;
    wire N__17860;
    wire N__17857;
    wire N__17854;
    wire N__17851;
    wire N__17848;
    wire N__17845;
    wire N__17842;
    wire N__17835;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17823;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17813;
    wire N__17808;
    wire N__17805;
    wire N__17802;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17790;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17775;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17765;
    wire N__17760;
    wire N__17757;
    wire N__17754;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17742;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17730;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17715;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17700;
    wire N__17697;
    wire N__17694;
    wire N__17691;
    wire N__17688;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17676;
    wire N__17675;
    wire N__17674;
    wire N__17671;
    wire N__17670;
    wire N__17667;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17653;
    wire N__17650;
    wire N__17649;
    wire N__17646;
    wire N__17641;
    wire N__17638;
    wire N__17635;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17617;
    wire N__17610;
    wire N__17607;
    wire N__17604;
    wire N__17601;
    wire N__17598;
    wire N__17595;
    wire N__17594;
    wire N__17593;
    wire N__17592;
    wire N__17591;
    wire N__17590;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17562;
    wire N__17561;
    wire N__17558;
    wire N__17557;
    wire N__17556;
    wire N__17555;
    wire N__17554;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17538;
    wire N__17529;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17514;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17502;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17490;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17480;
    wire N__17475;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17463;
    wire N__17460;
    wire N__17457;
    wire N__17454;
    wire N__17451;
    wire N__17448;
    wire N__17445;
    wire N__17442;
    wire N__17441;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17427;
    wire N__17424;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17409;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17394;
    wire N__17391;
    wire N__17390;
    wire N__17389;
    wire N__17388;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17374;
    wire N__17373;
    wire N__17372;
    wire N__17371;
    wire N__17370;
    wire N__17363;
    wire N__17354;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17328;
    wire N__17325;
    wire N__17322;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17307;
    wire N__17304;
    wire N__17301;
    wire N__17300;
    wire N__17299;
    wire N__17298;
    wire N__17297;
    wire N__17294;
    wire N__17293;
    wire N__17292;
    wire N__17289;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17278;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17266;
    wire N__17261;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17236;
    wire N__17233;
    wire N__17232;
    wire N__17227;
    wire N__17224;
    wire N__17219;
    wire N__17214;
    wire N__17209;
    wire N__17206;
    wire N__17201;
    wire N__17192;
    wire N__17187;
    wire N__17184;
    wire N__17183;
    wire N__17180;
    wire N__17177;
    wire N__17172;
    wire N__17169;
    wire N__17166;
    wire N__17163;
    wire N__17160;
    wire N__17157;
    wire N__17154;
    wire N__17151;
    wire N__17148;
    wire N__17145;
    wire N__17142;
    wire N__17139;
    wire N__17136;
    wire N__17133;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17121;
    wire N__17120;
    wire N__17117;
    wire N__17114;
    wire N__17109;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17094;
    wire N__17093;
    wire N__17090;
    wire N__17087;
    wire N__17082;
    wire N__17081;
    wire N__17078;
    wire N__17075;
    wire N__17072;
    wire N__17067;
    wire N__17066;
    wire N__17063;
    wire N__17060;
    wire N__17055;
    wire N__17052;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17040;
    wire N__17037;
    wire N__17036;
    wire N__17035;
    wire N__17032;
    wire N__17027;
    wire N__17022;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17014;
    wire N__17011;
    wire N__17008;
    wire N__17005;
    wire N__17004;
    wire N__17001;
    wire N__16996;
    wire N__16993;
    wire N__16986;
    wire N__16983;
    wire N__16980;
    wire N__16977;
    wire N__16974;
    wire N__16971;
    wire N__16970;
    wire N__16969;
    wire N__16968;
    wire N__16965;
    wire N__16962;
    wire N__16957;
    wire N__16954;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16932;
    wire N__16929;
    wire N__16926;
    wire N__16923;
    wire N__16920;
    wire N__16917;
    wire N__16914;
    wire N__16911;
    wire N__16910;
    wire N__16909;
    wire N__16908;
    wire N__16907;
    wire N__16906;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16896;
    wire N__16895;
    wire N__16894;
    wire N__16891;
    wire N__16884;
    wire N__16881;
    wire N__16878;
    wire N__16873;
    wire N__16868;
    wire N__16865;
    wire N__16864;
    wire N__16861;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16833;
    wire N__16826;
    wire N__16823;
    wire N__16818;
    wire N__16815;
    wire N__16812;
    wire N__16809;
    wire N__16808;
    wire N__16807;
    wire N__16804;
    wire N__16801;
    wire N__16798;
    wire N__16795;
    wire N__16788;
    wire N__16787;
    wire N__16784;
    wire N__16783;
    wire N__16782;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16764;
    wire N__16761;
    wire N__16758;
    wire N__16755;
    wire N__16752;
    wire N__16749;
    wire N__16742;
    wire N__16737;
    wire N__16734;
    wire N__16731;
    wire N__16728;
    wire N__16725;
    wire N__16722;
    wire N__16721;
    wire N__16718;
    wire N__16715;
    wire N__16712;
    wire N__16707;
    wire N__16706;
    wire N__16705;
    wire N__16704;
    wire N__16703;
    wire N__16702;
    wire N__16701;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16693;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16681;
    wire N__16676;
    wire N__16671;
    wire N__16664;
    wire N__16653;
    wire N__16650;
    wire N__16647;
    wire N__16646;
    wire N__16645;
    wire N__16644;
    wire N__16641;
    wire N__16634;
    wire N__16629;
    wire N__16628;
    wire N__16627;
    wire N__16624;
    wire N__16623;
    wire N__16620;
    wire N__16613;
    wire N__16608;
    wire N__16607;
    wire N__16606;
    wire N__16605;
    wire N__16602;
    wire N__16599;
    wire N__16596;
    wire N__16591;
    wire N__16584;
    wire N__16583;
    wire N__16582;
    wire N__16581;
    wire N__16578;
    wire N__16575;
    wire N__16570;
    wire N__16563;
    wire N__16562;
    wire N__16559;
    wire N__16558;
    wire N__16557;
    wire N__16556;
    wire N__16551;
    wire N__16544;
    wire N__16539;
    wire N__16536;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16528;
    wire N__16527;
    wire N__16526;
    wire N__16525;
    wire N__16524;
    wire N__16521;
    wire N__16518;
    wire N__16515;
    wire N__16512;
    wire N__16505;
    wire N__16502;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16471;
    wire N__16464;
    wire N__16461;
    wire N__16460;
    wire N__16459;
    wire N__16458;
    wire N__16457;
    wire N__16456;
    wire N__16453;
    wire N__16448;
    wire N__16441;
    wire N__16436;
    wire N__16435;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16410;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16397;
    wire N__16396;
    wire N__16395;
    wire N__16392;
    wire N__16389;
    wire N__16386;
    wire N__16383;
    wire N__16378;
    wire N__16371;
    wire N__16368;
    wire N__16367;
    wire N__16362;
    wire N__16359;
    wire N__16356;
    wire N__16355;
    wire N__16354;
    wire N__16351;
    wire N__16346;
    wire N__16345;
    wire N__16344;
    wire N__16343;
    wire N__16338;
    wire N__16333;
    wire N__16330;
    wire N__16323;
    wire N__16322;
    wire N__16319;
    wire N__16316;
    wire N__16311;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16299;
    wire N__16298;
    wire N__16297;
    wire N__16294;
    wire N__16289;
    wire N__16288;
    wire N__16287;
    wire N__16286;
    wire N__16285;
    wire N__16284;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16254;
    wire N__16245;
    wire N__16242;
    wire N__16239;
    wire N__16236;
    wire N__16233;
    wire N__16232;
    wire N__16231;
    wire N__16230;
    wire N__16229;
    wire N__16228;
    wire N__16227;
    wire N__16224;
    wire N__16219;
    wire N__16210;
    wire N__16207;
    wire N__16202;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16190;
    wire N__16189;
    wire N__16184;
    wire N__16181;
    wire N__16178;
    wire N__16175;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16154;
    wire N__16153;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16141;
    wire N__16138;
    wire N__16131;
    wire N__16128;
    wire N__16125;
    wire N__16124;
    wire N__16123;
    wire N__16122;
    wire N__16119;
    wire N__16116;
    wire N__16113;
    wire N__16110;
    wire N__16101;
    wire N__16098;
    wire N__16095;
    wire N__16092;
    wire N__16089;
    wire N__16086;
    wire N__16085;
    wire N__16084;
    wire N__16083;
    wire N__16080;
    wire N__16077;
    wire N__16074;
    wire N__16071;
    wire N__16070;
    wire N__16067;
    wire N__16064;
    wire N__16063;
    wire N__16062;
    wire N__16061;
    wire N__16058;
    wire N__16057;
    wire N__16056;
    wire N__16051;
    wire N__16048;
    wire N__16045;
    wire N__16038;
    wire N__16035;
    wire N__16030;
    wire N__16025;
    wire N__16014;
    wire N__16011;
    wire N__16008;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15987;
    wire N__15984;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15972;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15960;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15945;
    wire N__15944;
    wire N__15941;
    wire N__15938;
    wire N__15933;
    wire N__15930;
    wire N__15927;
    wire N__15924;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15912;
    wire N__15911;
    wire N__15908;
    wire N__15905;
    wire N__15900;
    wire N__15899;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15885;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15873;
    wire N__15870;
    wire N__15867;
    wire N__15864;
    wire N__15863;
    wire N__15862;
    wire N__15861;
    wire N__15860;
    wire N__15857;
    wire N__15856;
    wire N__15853;
    wire N__15850;
    wire N__15845;
    wire N__15842;
    wire N__15839;
    wire N__15836;
    wire N__15825;
    wire N__15824;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15810;
    wire N__15807;
    wire N__15804;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15792;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15780;
    wire N__15779;
    wire N__15778;
    wire N__15777;
    wire N__15776;
    wire N__15775;
    wire N__15774;
    wire N__15773;
    wire N__15768;
    wire N__15761;
    wire N__15754;
    wire N__15751;
    wire N__15744;
    wire N__15743;
    wire N__15742;
    wire N__15739;
    wire N__15738;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15720;
    wire N__15719;
    wire N__15718;
    wire N__15715;
    wire N__15710;
    wire N__15705;
    wire N__15704;
    wire N__15703;
    wire N__15700;
    wire N__15695;
    wire N__15690;
    wire N__15689;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15675;
    wire N__15674;
    wire N__15673;
    wire N__15670;
    wire N__15665;
    wire N__15660;
    wire N__15657;
    wire N__15654;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15642;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15630;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15615;
    wire N__15614;
    wire N__15611;
    wire N__15608;
    wire N__15603;
    wire N__15600;
    wire N__15597;
    wire N__15594;
    wire N__15593;
    wire N__15590;
    wire N__15587;
    wire N__15582;
    wire N__15581;
    wire N__15578;
    wire N__15575;
    wire N__15570;
    wire N__15569;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15555;
    wire N__15554;
    wire N__15551;
    wire N__15548;
    wire N__15543;
    wire N__15540;
    wire N__15537;
    wire N__15534;
    wire N__15533;
    wire N__15530;
    wire N__15527;
    wire N__15522;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15510;
    wire N__15509;
    wire N__15506;
    wire N__15503;
    wire N__15500;
    wire N__15495;
    wire N__15494;
    wire N__15491;
    wire N__15488;
    wire N__15483;
    wire N__15480;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15465;
    wire N__15462;
    wire N__15459;
    wire N__15456;
    wire N__15453;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15441;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15429;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15414;
    wire N__15413;
    wire N__15410;
    wire N__15407;
    wire N__15402;
    wire N__15399;
    wire N__15398;
    wire N__15395;
    wire N__15392;
    wire N__15389;
    wire N__15386;
    wire N__15385;
    wire N__15380;
    wire N__15377;
    wire N__15372;
    wire N__15369;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15357;
    wire N__15356;
    wire N__15353;
    wire N__15350;
    wire N__15345;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15330;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15300;
    wire N__15299;
    wire N__15296;
    wire N__15293;
    wire N__15288;
    wire N__15287;
    wire N__15284;
    wire N__15281;
    wire N__15278;
    wire N__15273;
    wire N__15272;
    wire N__15269;
    wire N__15266;
    wire N__15261;
    wire N__15258;
    wire N__15255;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15243;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15231;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15216;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15204;
    wire N__15201;
    wire N__15198;
    wire N__15195;
    wire N__15192;
    wire N__15191;
    wire N__15190;
    wire N__15189;
    wire N__15186;
    wire N__15179;
    wire N__15174;
    wire N__15171;
    wire N__15168;
    wire N__15165;
    wire N__15164;
    wire N__15163;
    wire N__15158;
    wire N__15155;
    wire N__15152;
    wire N__15147;
    wire N__15144;
    wire N__15141;
    wire N__15138;
    wire N__15135;
    wire N__15132;
    wire N__15129;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15119;
    wire N__15116;
    wire N__15113;
    wire N__15110;
    wire N__15105;
    wire N__15102;
    wire N__15099;
    wire N__15098;
    wire N__15097;
    wire N__15094;
    wire N__15089;
    wire N__15084;
    wire N__15081;
    wire N__15080;
    wire N__15079;
    wire N__15076;
    wire N__15073;
    wire N__15070;
    wire N__15063;
    wire N__15060;
    wire N__15059;
    wire N__15058;
    wire N__15055;
    wire N__15050;
    wire N__15045;
    wire N__15042;
    wire N__15039;
    wire N__15038;
    wire N__15037;
    wire N__15036;
    wire N__15035;
    wire N__15034;
    wire N__15033;
    wire N__15030;
    wire N__15029;
    wire N__15028;
    wire N__15025;
    wire N__15022;
    wire N__15019;
    wire N__15014;
    wire N__15011;
    wire N__15002;
    wire N__14991;
    wire N__14990;
    wire N__14987;
    wire N__14986;
    wire N__14985;
    wire N__14984;
    wire N__14983;
    wire N__14982;
    wire N__14981;
    wire N__14980;
    wire N__14977;
    wire N__14974;
    wire N__14971;
    wire N__14962;
    wire N__14955;
    wire N__14946;
    wire N__14945;
    wire N__14944;
    wire N__14943;
    wire N__14942;
    wire N__14939;
    wire N__14936;
    wire N__14935;
    wire N__14934;
    wire N__14931;
    wire N__14930;
    wire N__14925;
    wire N__14922;
    wire N__14917;
    wire N__14910;
    wire N__14907;
    wire N__14898;
    wire N__14897;
    wire N__14896;
    wire N__14895;
    wire N__14894;
    wire N__14893;
    wire N__14892;
    wire N__14887;
    wire N__14886;
    wire N__14885;
    wire N__14882;
    wire N__14877;
    wire N__14872;
    wire N__14869;
    wire N__14864;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14844;
    wire N__14841;
    wire N__14838;
    wire N__14835;
    wire N__14834;
    wire N__14833;
    wire N__14830;
    wire N__14825;
    wire N__14820;
    wire N__14817;
    wire N__14814;
    wire N__14811;
    wire N__14808;
    wire N__14805;
    wire N__14802;
    wire N__14801;
    wire N__14800;
    wire N__14799;
    wire N__14798;
    wire N__14797;
    wire N__14796;
    wire N__14795;
    wire N__14792;
    wire N__14791;
    wire N__14788;
    wire N__14787;
    wire N__14784;
    wire N__14783;
    wire N__14780;
    wire N__14779;
    wire N__14778;
    wire N__14775;
    wire N__14774;
    wire N__14771;
    wire N__14770;
    wire N__14769;
    wire N__14766;
    wire N__14763;
    wire N__14746;
    wire N__14735;
    wire N__14730;
    wire N__14721;
    wire N__14718;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14710;
    wire N__14709;
    wire N__14706;
    wire N__14703;
    wire N__14700;
    wire N__14697;
    wire N__14696;
    wire N__14687;
    wire N__14684;
    wire N__14683;
    wire N__14682;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14667;
    wire N__14658;
    wire N__14655;
    wire N__14652;
    wire N__14651;
    wire N__14648;
    wire N__14647;
    wire N__14646;
    wire N__14645;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14634;
    wire N__14633;
    wire N__14630;
    wire N__14625;
    wire N__14622;
    wire N__14619;
    wire N__14616;
    wire N__14615;
    wire N__14612;
    wire N__14609;
    wire N__14606;
    wire N__14603;
    wire N__14600;
    wire N__14595;
    wire N__14588;
    wire N__14577;
    wire N__14574;
    wire N__14571;
    wire N__14568;
    wire N__14565;
    wire N__14564;
    wire N__14559;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14544;
    wire N__14543;
    wire N__14540;
    wire N__14539;
    wire N__14536;
    wire N__14535;
    wire N__14534;
    wire N__14531;
    wire N__14526;
    wire N__14523;
    wire N__14522;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14504;
    wire N__14493;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14478;
    wire N__14477;
    wire N__14476;
    wire N__14475;
    wire N__14474;
    wire N__14473;
    wire N__14470;
    wire N__14467;
    wire N__14466;
    wire N__14459;
    wire N__14458;
    wire N__14457;
    wire N__14454;
    wire N__14447;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14436;
    wire N__14435;
    wire N__14434;
    wire N__14433;
    wire N__14432;
    wire N__14431;
    wire N__14430;
    wire N__14429;
    wire N__14426;
    wire N__14423;
    wire N__14420;
    wire N__14413;
    wire N__14404;
    wire N__14395;
    wire N__14382;
    wire N__14381;
    wire N__14376;
    wire N__14375;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14359;
    wire N__14356;
    wire N__14349;
    wire N__14348;
    wire N__14345;
    wire N__14344;
    wire N__14341;
    wire N__14334;
    wire N__14331;
    wire N__14328;
    wire N__14325;
    wire N__14324;
    wire N__14323;
    wire N__14322;
    wire N__14321;
    wire N__14320;
    wire N__14319;
    wire N__14318;
    wire N__14315;
    wire N__14312;
    wire N__14309;
    wire N__14302;
    wire N__14297;
    wire N__14286;
    wire N__14285;
    wire N__14284;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14274;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14264;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14256;
    wire N__14253;
    wire N__14248;
    wire N__14245;
    wire N__14242;
    wire N__14237;
    wire N__14226;
    wire N__14225;
    wire N__14224;
    wire N__14223;
    wire N__14220;
    wire N__14219;
    wire N__14218;
    wire N__14215;
    wire N__14212;
    wire N__14211;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14199;
    wire N__14198;
    wire N__14197;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14174;
    wire N__14163;
    wire N__14162;
    wire N__14159;
    wire N__14156;
    wire N__14153;
    wire N__14152;
    wire N__14151;
    wire N__14150;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14140;
    wire N__14139;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14124;
    wire N__14121;
    wire N__14116;
    wire N__14103;
    wire N__14102;
    wire N__14099;
    wire N__14096;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14088;
    wire N__14087;
    wire N__14084;
    wire N__14083;
    wire N__14078;
    wire N__14077;
    wire N__14074;
    wire N__14071;
    wire N__14070;
    wire N__14067;
    wire N__14064;
    wire N__14061;
    wire N__14058;
    wire N__14053;
    wire N__14050;
    wire N__14037;
    wire N__14036;
    wire N__14035;
    wire N__14034;
    wire N__14033;
    wire N__14030;
    wire N__14029;
    wire N__14028;
    wire N__14025;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14017;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__13997;
    wire N__13992;
    wire N__13977;
    wire N__13976;
    wire N__13975;
    wire N__13974;
    wire N__13971;
    wire N__13970;
    wire N__13967;
    wire N__13966;
    wire N__13965;
    wire N__13964;
    wire N__13961;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13953;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13935;
    wire N__13930;
    wire N__13927;
    wire N__13922;
    wire N__13905;
    wire N__13904;
    wire N__13903;
    wire N__13902;
    wire N__13901;
    wire N__13900;
    wire N__13897;
    wire N__13896;
    wire N__13895;
    wire N__13894;
    wire N__13893;
    wire N__13890;
    wire N__13887;
    wire N__13882;
    wire N__13879;
    wire N__13874;
    wire N__13865;
    wire N__13854;
    wire N__13851;
    wire N__13848;
    wire N__13845;
    wire N__13842;
    wire N__13839;
    wire N__13836;
    wire N__13833;
    wire N__13832;
    wire N__13827;
    wire N__13824;
    wire N__13821;
    wire N__13820;
    wire N__13815;
    wire N__13812;
    wire N__13811;
    wire N__13808;
    wire N__13803;
    wire N__13800;
    wire N__13799;
    wire N__13794;
    wire N__13791;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13779;
    wire N__13776;
    wire N__13775;
    wire N__13770;
    wire N__13767;
    wire N__13764;
    wire N__13761;
    wire N__13758;
    wire N__13757;
    wire N__13756;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13748;
    wire N__13745;
    wire N__13742;
    wire N__13741;
    wire N__13738;
    wire N__13733;
    wire N__13728;
    wire N__13725;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13707;
    wire N__13704;
    wire N__13701;
    wire N__13698;
    wire N__13695;
    wire N__13692;
    wire N__13689;
    wire N__13686;
    wire N__13683;
    wire N__13680;
    wire N__13677;
    wire N__13674;
    wire N__13671;
    wire N__13668;
    wire N__13665;
    wire N__13662;
    wire N__13659;
    wire N__13656;
    wire N__13653;
    wire N__13650;
    wire N__13647;
    wire N__13646;
    wire N__13645;
    wire N__13642;
    wire N__13639;
    wire N__13634;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13617;
    wire N__13614;
    wire N__13611;
    wire N__13608;
    wire N__13605;
    wire N__13602;
    wire N__13599;
    wire N__13596;
    wire N__13593;
    wire N__13590;
    wire N__13587;
    wire N__13584;
    wire N__13581;
    wire N__13580;
    wire N__13577;
    wire N__13576;
    wire N__13575;
    wire N__13572;
    wire N__13569;
    wire N__13566;
    wire N__13563;
    wire N__13560;
    wire N__13557;
    wire N__13554;
    wire N__13551;
    wire N__13542;
    wire N__13541;
    wire N__13540;
    wire N__13537;
    wire N__13532;
    wire N__13527;
    wire N__13524;
    wire N__13521;
    wire N__13518;
    wire N__13517;
    wire N__13516;
    wire N__13513;
    wire N__13508;
    wire N__13503;
    wire N__13500;
    wire N__13497;
    wire N__13494;
    wire N__13491;
    wire N__13488;
    wire N__13485;
    wire N__13482;
    wire N__13479;
    wire N__13476;
    wire N__13473;
    wire N__13470;
    wire N__13467;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13455;
    wire N__13452;
    wire N__13451;
    wire N__13450;
    wire N__13449;
    wire N__13448;
    wire N__13447;
    wire N__13442;
    wire N__13433;
    wire N__13428;
    wire N__13427;
    wire N__13426;
    wire N__13425;
    wire N__13424;
    wire N__13423;
    wire N__13420;
    wire N__13413;
    wire N__13408;
    wire N__13401;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13391;
    wire N__13388;
    wire N__13383;
    wire N__13380;
    wire N__13377;
    wire N__13374;
    wire N__13371;
    wire N__13368;
    wire N__13365;
    wire N__13362;
    wire N__13359;
    wire N__13356;
    wire N__13353;
    wire N__13350;
    wire N__13347;
    wire N__13344;
    wire N__13341;
    wire N__13340;
    wire N__13339;
    wire N__13336;
    wire N__13331;
    wire N__13326;
    wire N__13323;
    wire N__13322;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13308;
    wire N__13305;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13293;
    wire N__13290;
    wire N__13287;
    wire N__13284;
    wire N__13281;
    wire N__13278;
    wire N__13275;
    wire N__13272;
    wire N__13269;
    wire N__13266;
    wire N__13263;
    wire N__13262;
    wire N__13261;
    wire N__13258;
    wire N__13253;
    wire N__13252;
    wire N__13251;
    wire N__13250;
    wire N__13249;
    wire N__13246;
    wire N__13243;
    wire N__13238;
    wire N__13233;
    wire N__13224;
    wire N__13223;
    wire N__13218;
    wire N__13215;
    wire N__13212;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13188;
    wire N__13185;
    wire N__13182;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13167;
    wire N__13164;
    wire N__13161;
    wire N__13158;
    wire N__13157;
    wire N__13154;
    wire N__13151;
    wire N__13148;
    wire N__13145;
    wire N__13140;
    wire N__13137;
    wire N__13134;
    wire N__13131;
    wire N__13128;
    wire N__13127;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13113;
    wire N__13112;
    wire N__13111;
    wire N__13110;
    wire N__13109;
    wire N__13102;
    wire N__13097;
    wire N__13092;
    wire N__13091;
    wire N__13090;
    wire N__13087;
    wire N__13082;
    wire N__13077;
    wire N__13076;
    wire N__13075;
    wire N__13074;
    wire N__13073;
    wire N__13070;
    wire N__13063;
    wire N__13060;
    wire N__13057;
    wire N__13050;
    wire N__13047;
    wire N__13044;
    wire N__13041;
    wire N__13038;
    wire N__13037;
    wire N__13034;
    wire N__13031;
    wire N__13026;
    wire N__13023;
    wire N__13020;
    wire N__13019;
    wire N__13016;
    wire N__13013;
    wire N__13010;
    wire N__13007;
    wire N__13002;
    wire N__12999;
    wire N__12996;
    wire N__12993;
    wire N__12990;
    wire N__12989;
    wire N__12986;
    wire N__12983;
    wire N__12978;
    wire N__12975;
    wire N__12972;
    wire N__12969;
    wire N__12966;
    wire N__12963;
    wire N__12960;
    wire N__12957;
    wire N__12954;
    wire N__12951;
    wire N__12948;
    wire N__12945;
    wire N__12942;
    wire N__12939;
    wire N__12936;
    wire N__12935;
    wire N__12934;
    wire N__12933;
    wire N__12930;
    wire N__12927;
    wire N__12924;
    wire N__12921;
    wire N__12912;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12896;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12876;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12861;
    wire N__12858;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12840;
    wire N__12837;
    wire N__12834;
    wire N__12831;
    wire N__12828;
    wire N__12825;
    wire N__12822;
    wire N__12819;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12801;
    wire N__12798;
    wire N__12797;
    wire N__12794;
    wire N__12791;
    wire N__12788;
    wire N__12783;
    wire N__12780;
    wire N__12777;
    wire N__12774;
    wire N__12771;
    wire N__12768;
    wire N__12765;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12723;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12708;
    wire N__12705;
    wire N__12702;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12690;
    wire N__12687;
    wire N__12684;
    wire N__12681;
    wire N__12678;
    wire N__12675;
    wire N__12672;
    wire N__12669;
    wire N__12666;
    wire N__12663;
    wire N__12662;
    wire N__12659;
    wire N__12658;
    wire N__12655;
    wire N__12654;
    wire N__12651;
    wire N__12646;
    wire N__12643;
    wire N__12636;
    wire N__12633;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12618;
    wire N__12615;
    wire N__12612;
    wire N__12611;
    wire N__12608;
    wire N__12607;
    wire N__12604;
    wire N__12597;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12585;
    wire N__12582;
    wire N__12579;
    wire N__12576;
    wire N__12573;
    wire N__12570;
    wire N__12567;
    wire N__12566;
    wire N__12563;
    wire N__12562;
    wire N__12559;
    wire N__12558;
    wire N__12555;
    wire N__12550;
    wire N__12547;
    wire N__12540;
    wire N__12537;
    wire N__12536;
    wire N__12533;
    wire N__12532;
    wire N__12529;
    wire N__12522;
    wire N__12519;
    wire N__12516;
    wire N__12513;
    wire N__12510;
    wire N__12507;
    wire N__12504;
    wire N__12501;
    wire N__12498;
    wire N__12495;
    wire N__12492;
    wire N__12489;
    wire N__12486;
    wire N__12483;
    wire N__12480;
    wire N__12477;
    wire N__12474;
    wire N__12471;
    wire N__12468;
    wire N__12465;
    wire N__12462;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12452;
    wire N__12449;
    wire N__12448;
    wire N__12445;
    wire N__12444;
    wire N__12441;
    wire N__12436;
    wire N__12433;
    wire N__12426;
    wire N__12423;
    wire N__12422;
    wire N__12419;
    wire N__12418;
    wire N__12415;
    wire N__12408;
    wire N__12405;
    wire N__12402;
    wire N__12401;
    wire N__12398;
    wire N__12395;
    wire N__12392;
    wire N__12389;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12363;
    wire N__12360;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12348;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12299;
    wire N__12296;
    wire N__12295;
    wire N__12292;
    wire N__12291;
    wire N__12288;
    wire N__12283;
    wire N__12280;
    wire N__12273;
    wire N__12270;
    wire N__12269;
    wire N__12266;
    wire N__12265;
    wire N__12262;
    wire N__12255;
    wire N__12252;
    wire N__12249;
    wire N__12246;
    wire N__12243;
    wire N__12240;
    wire N__12237;
    wire N__12234;
    wire N__12231;
    wire N__12228;
    wire N__12225;
    wire N__12222;
    wire N__12219;
    wire N__12216;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12204;
    wire N__12201;
    wire N__12200;
    wire N__12199;
    wire N__12196;
    wire N__12195;
    wire N__12192;
    wire N__12187;
    wire N__12184;
    wire N__12177;
    wire N__12174;
    wire N__12171;
    wire N__12168;
    wire N__12165;
    wire N__12162;
    wire N__12159;
    wire N__12156;
    wire N__12153;
    wire N__12152;
    wire N__12149;
    wire N__12148;
    wire N__12145;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12123;
    wire N__12120;
    wire N__12117;
    wire N__12114;
    wire N__12113;
    wire N__12110;
    wire N__12109;
    wire N__12106;
    wire N__12105;
    wire N__12102;
    wire N__12097;
    wire N__12094;
    wire N__12087;
    wire N__12084;
    wire N__12083;
    wire N__12080;
    wire N__12079;
    wire N__12076;
    wire N__12069;
    wire N__12066;
    wire N__12063;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12051;
    wire N__12048;
    wire N__12045;
    wire N__12044;
    wire N__12041;
    wire N__12040;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12022;
    wire N__12015;
    wire N__12012;
    wire N__12011;
    wire N__12008;
    wire N__12007;
    wire N__12004;
    wire N__12003;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11991;
    wire N__11988;
    wire N__11979;
    wire N__11976;
    wire N__11973;
    wire N__11972;
    wire N__11969;
    wire N__11968;
    wire N__11965;
    wire N__11964;
    wire N__11961;
    wire N__11958;
    wire N__11955;
    wire N__11952;
    wire N__11949;
    wire N__11940;
    wire N__11937;
    wire N__11934;
    wire N__11933;
    wire N__11932;
    wire N__11929;
    wire N__11926;
    wire N__11925;
    wire N__11922;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11908;
    wire N__11905;
    wire N__11900;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11885;
    wire N__11882;
    wire N__11879;
    wire N__11878;
    wire N__11875;
    wire N__11872;
    wire N__11871;
    wire N__11868;
    wire N__11867;
    wire N__11866;
    wire N__11863;
    wire N__11860;
    wire N__11857;
    wire N__11854;
    wire N__11851;
    wire N__11848;
    wire N__11835;
    wire N__11834;
    wire N__11831;
    wire N__11828;
    wire N__11825;
    wire N__11822;
    wire N__11817;
    wire N__11814;
    wire N__11811;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11783;
    wire N__11780;
    wire N__11777;
    wire N__11776;
    wire N__11773;
    wire N__11770;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11757;
    wire N__11748;
    wire N__11745;
    wire N__11744;
    wire N__11741;
    wire N__11738;
    wire N__11737;
    wire N__11734;
    wire N__11733;
    wire N__11730;
    wire N__11727;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11709;
    wire N__11706;
    wire N__11705;
    wire N__11702;
    wire N__11699;
    wire N__11696;
    wire N__11695;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11667;
    wire N__11664;
    wire N__11663;
    wire N__11660;
    wire N__11657;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11628;
    wire N__11625;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11617;
    wire N__11614;
    wire N__11611;
    wire N__11610;
    wire N__11607;
    wire N__11604;
    wire N__11601;
    wire N__11598;
    wire N__11589;
    wire N__11586;
    wire N__11585;
    wire N__11582;
    wire N__11581;
    wire N__11578;
    wire N__11575;
    wire N__11574;
    wire N__11571;
    wire N__11568;
    wire N__11565;
    wire N__11562;
    wire N__11553;
    wire N__11550;
    wire N__11547;
    wire N__11546;
    wire N__11543;
    wire N__11542;
    wire N__11541;
    wire N__11538;
    wire N__11535;
    wire N__11532;
    wire N__11529;
    wire N__11526;
    wire N__11523;
    wire N__11520;
    wire N__11511;
    wire N__11508;
    wire N__11507;
    wire N__11504;
    wire N__11503;
    wire N__11502;
    wire N__11499;
    wire N__11496;
    wire N__11493;
    wire N__11490;
    wire N__11485;
    wire N__11478;
    wire N__11475;
    wire N__11474;
    wire N__11471;
    wire N__11468;
    wire N__11463;
    wire N__11460;
    wire N__11459;
    wire N__11456;
    wire N__11453;
    wire N__11448;
    wire N__11445;
    wire N__11444;
    wire N__11441;
    wire N__11438;
    wire N__11433;
    wire N__11430;
    wire N__11427;
    wire N__11426;
    wire N__11423;
    wire N__11420;
    wire N__11417;
    wire N__11412;
    wire N__11409;
    wire N__11406;
    wire N__11405;
    wire N__11404;
    wire N__11401;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11385;
    wire N__11384;
    wire N__11383;
    wire N__11382;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11357;
    wire N__11354;
    wire N__11349;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11341;
    wire N__11338;
    wire N__11335;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11313;
    wire N__11310;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11295;
    wire N__11292;
    wire N__11289;
    wire N__11286;
    wire N__11283;
    wire N__11274;
    wire N__11271;
    wire N__11270;
    wire N__11267;
    wire N__11264;
    wire N__11259;
    wire N__11256;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11244;
    wire N__11241;
    wire N__11240;
    wire N__11237;
    wire N__11234;
    wire N__11229;
    wire N__11226;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11214;
    wire N__11211;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11196;
    wire N__11193;
    wire N__11192;
    wire N__11189;
    wire N__11186;
    wire N__11181;
    wire N__11178;
    wire N__11177;
    wire N__11174;
    wire N__11171;
    wire N__11166;
    wire N__11163;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11148;
    wire N__11145;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11130;
    wire N__11127;
    wire N__11124;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11111;
    wire N__11110;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11098;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11084;
    wire N__11083;
    wire N__11080;
    wire N__11077;
    wire N__11074;
    wire N__11071;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11043;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11031;
    wire N__11028;
    wire N__11027;
    wire N__11024;
    wire N__11021;
    wire N__11016;
    wire N__11013;
    wire N__11010;
    wire N__11007;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10994;
    wire N__10991;
    wire N__10988;
    wire N__10985;
    wire N__10980;
    wire N__10977;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10967;
    wire N__10962;
    wire N__10959;
    wire N__10956;
    wire N__10953;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10938;
    wire N__10935;
    wire N__10932;
    wire N__10929;
    wire N__10926;
    wire N__10923;
    wire N__10920;
    wire N__10917;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10907;
    wire N__10902;
    wire N__10899;
    wire N__10896;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10875;
    wire N__10872;
    wire N__10869;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10839;
    wire N__10836;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10806;
    wire N__10803;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10773;
    wire N__10770;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10758;
    wire N__10755;
    wire N__10752;
    wire N__10749;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10734;
    wire N__10733;
    wire N__10732;
    wire N__10729;
    wire N__10722;
    wire N__10719;
    wire N__10716;
    wire N__10713;
    wire N__10710;
    wire N__10707;
    wire N__10704;
    wire N__10701;
    wire N__10698;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10686;
    wire N__10683;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10670;
    wire N__10669;
    wire N__10666;
    wire N__10665;
    wire N__10662;
    wire N__10657;
    wire N__10654;
    wire N__10647;
    wire N__10644;
    wire N__10641;
    wire N__10638;
    wire N__10635;
    wire N__10632;
    wire N__10629;
    wire N__10628;
    wire N__10625;
    wire N__10624;
    wire N__10621;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10605;
    wire N__10602;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10587;
    wire N__10584;
    wire N__10581;
    wire N__10578;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10563;
    wire N__10560;
    wire N__10557;
    wire N__10554;
    wire N__10551;
    wire N__10550;
    wire N__10547;
    wire N__10546;
    wire N__10543;
    wire N__10536;
    wire N__10533;
    wire N__10530;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10515;
    wire N__10512;
    wire N__10509;
    wire N__10508;
    wire N__10505;
    wire N__10504;
    wire N__10503;
    wire N__10502;
    wire N__10497;
    wire N__10494;
    wire N__10489;
    wire N__10482;
    wire N__10479;
    wire N__10476;
    wire N__10473;
    wire N__10470;
    wire N__10467;
    wire N__10464;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10452;
    wire N__10449;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10419;
    wire N__10418;
    wire N__10413;
    wire N__10410;
    wire N__10407;
    wire N__10404;
    wire N__10401;
    wire N__10398;
    wire N__10395;
    wire N__10392;
    wire N__10389;
    wire N__10386;
    wire N__10383;
    wire N__10380;
    wire N__10377;
    wire N__10374;
    wire N__10371;
    wire N__10368;
    wire N__10365;
    wire N__10362;
    wire N__10359;
    wire N__10356;
    wire N__10353;
    wire N__10350;
    wire N__10347;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10335;
    wire N__10332;
    wire N__10329;
    wire N__10326;
    wire N__10323;
    wire N__10320;
    wire N__10317;
    wire N__10314;
    wire N__10311;
    wire N__10308;
    wire N__10305;
    wire N__10302;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10290;
    wire N__10287;
    wire N__10284;
    wire N__10281;
    wire N__10278;
    wire N__10277;
    wire N__10276;
    wire N__10275;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10248;
    wire N__10239;
    wire N__10238;
    wire N__10235;
    wire N__10234;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10222;
    wire N__10217;
    wire N__10212;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10200;
    wire N__10197;
    wire N__10194;
    wire N__10191;
    wire N__10188;
    wire N__10185;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10170;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10152;
    wire N__10149;
    wire N__10146;
    wire N__10143;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10135;
    wire N__10130;
    wire N__10129;
    wire N__10126;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10114;
    wire N__10107;
    wire N__10104;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10086;
    wire N__10083;
    wire N__10080;
    wire N__10077;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10062;
    wire N__10059;
    wire N__10056;
    wire N__10055;
    wire N__10052;
    wire N__10051;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10039;
    wire N__10036;
    wire N__10033;
    wire N__10030;
    wire N__10027;
    wire N__10020;
    wire N__10017;
    wire N__10014;
    wire N__10011;
    wire N__10008;
    wire N__10005;
    wire N__10002;
    wire N__9999;
    wire N__9996;
    wire N__9993;
    wire N__9990;
    wire N__9987;
    wire N__9984;
    wire N__9981;
    wire N__9980;
    wire N__9977;
    wire N__9976;
    wire N__9973;
    wire N__9966;
    wire N__9963;
    wire N__9960;
    wire N__9957;
    wire N__9954;
    wire N__9951;
    wire N__9948;
    wire N__9945;
    wire N__9942;
    wire N__9939;
    wire N__9936;
    wire N__9933;
    wire N__9930;
    wire N__9927;
    wire N__9924;
    wire N__9921;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9909;
    wire N__9906;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9882;
    wire N__9879;
    wire N__9876;
    wire N__9873;
    wire N__9870;
    wire N__9867;
    wire N__9864;
    wire N__9861;
    wire N__9858;
    wire N__9855;
    wire N__9852;
    wire N__9849;
    wire N__9846;
    wire N__9843;
    wire N__9840;
    wire N__9837;
    wire N__9834;
    wire N__9831;
    wire N__9828;
    wire N__9825;
    wire N__9822;
    wire N__9819;
    wire N__9816;
    wire N__9813;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9805;
    wire N__9802;
    wire N__9799;
    wire N__9796;
    wire N__9793;
    wire N__9790;
    wire N__9787;
    wire N__9780;
    wire N__9777;
    wire N__9774;
    wire N__9771;
    wire N__9768;
    wire N__9765;
    wire N__9762;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9744;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9736;
    wire N__9733;
    wire N__9730;
    wire N__9727;
    wire N__9720;
    wire N__9717;
    wire N__9714;
    wire N__9711;
    wire N__9708;
    wire N__9705;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9690;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9678;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9666;
    wire N__9665;
    wire N__9662;
    wire N__9661;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9647;
    wire N__9642;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9630;
    wire N__9629;
    wire N__9626;
    wire N__9623;
    wire N__9618;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9608;
    wire N__9603;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9591;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9579;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9567;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9552;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9540;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9528;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9516;
    wire N__9513;
    wire N__9510;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9498;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9486;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9471;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9459;
    wire N__9456;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9444;
    wire N__9441;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9429;
    wire N__9426;
    wire N__9423;
    wire N__9420;
    wire N__9419;
    wire N__9416;
    wire N__9415;
    wire N__9414;
    wire N__9411;
    wire N__9404;
    wire N__9399;
    wire N__9396;
    wire N__9393;
    wire N__9392;
    wire N__9389;
    wire N__9388;
    wire N__9385;
    wire N__9378;
    wire N__9375;
    wire N__9372;
    wire N__9369;
    wire N__9366;
    wire N__9363;
    wire N__9360;
    wire N__9357;
    wire N__9354;
    wire N__9351;
    wire N__9348;
    wire N__9345;
    wire N__9342;
    wire N__9339;
    wire N__9336;
    wire N__9333;
    wire N__9330;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9311;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9292;
    wire N__9289;
    wire N__9286;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9270;
    wire N__9267;
    wire N__9264;
    wire N__9261;
    wire N__9258;
    wire N__9255;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9200;
    wire N__9199;
    wire N__9196;
    wire N__9195;
    wire N__9192;
    wire N__9187;
    wire N__9184;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9159;
    wire N__9156;
    wire N__9153;
    wire N__9150;
    wire N__9147;
    wire N__9144;
    wire N__9141;
    wire N__9138;
    wire N__9135;
    wire N__9132;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9114;
    wire N__9111;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9093;
    wire N__9090;
    wire N__9087;
    wire N__9084;
    wire N__9081;
    wire N__9078;
    wire N__9075;
    wire N__9072;
    wire N__9071;
    wire N__9068;
    wire N__9067;
    wire N__9064;
    wire N__9063;
    wire N__9062;
    wire N__9059;
    wire N__9054;
    wire N__9051;
    wire N__9048;
    wire N__9039;
    wire N__9038;
    wire N__9035;
    wire N__9034;
    wire N__9029;
    wire N__9028;
    wire N__9027;
    wire N__9026;
    wire N__9025;
    wire N__9022;
    wire N__9019;
    wire N__9016;
    wire N__9009;
    wire N__9000;
    wire N__8999;
    wire N__8998;
    wire N__8995;
    wire N__8994;
    wire N__8993;
    wire N__8990;
    wire N__8985;
    wire N__8982;
    wire N__8979;
    wire N__8970;
    wire N__8967;
    wire N__8964;
    wire N__8961;
    wire N__8958;
    wire N__8955;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8943;
    wire N__8940;
    wire N__8937;
    wire N__8934;
    wire N__8931;
    wire N__8928;
    wire N__8925;
    wire N__8922;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8910;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8898;
    wire N__8895;
    wire N__8892;
    wire N__8889;
    wire N__8886;
    wire N__8883;
    wire N__8880;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8864;
    wire N__8861;
    wire N__8860;
    wire N__8857;
    wire N__8850;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8838;
    wire N__8835;
    wire N__8834;
    wire N__8831;
    wire N__8830;
    wire N__8827;
    wire N__8820;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8808;
    wire N__8805;
    wire N__8802;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8781;
    wire N__8778;
    wire N__8775;
    wire N__8772;
    wire N__8769;
    wire N__8766;
    wire N__8763;
    wire N__8760;
    wire N__8757;
    wire N__8754;
    wire N__8751;
    wire N__8748;
    wire N__8745;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8717;
    wire N__8714;
    wire N__8713;
    wire N__8710;
    wire N__8703;
    wire N__8700;
    wire N__8697;
    wire N__8694;
    wire N__8691;
    wire N__8688;
    wire N__8685;
    wire N__8682;
    wire N__8679;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8648;
    wire N__8645;
    wire N__8644;
    wire N__8641;
    wire N__8634;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8622;
    wire N__8619;
    wire N__8616;
    wire N__8613;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8595;
    wire N__8592;
    wire N__8589;
    wire N__8586;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8574;
    wire N__8571;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8547;
    wire N__8544;
    wire N__8541;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8529;
    wire N__8526;
    wire N__8523;
    wire N__8520;
    wire N__8517;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8489;
    wire N__8486;
    wire N__8485;
    wire N__8482;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8466;
    wire N__8463;
    wire N__8460;
    wire N__8457;
    wire N__8456;
    wire N__8453;
    wire N__8452;
    wire N__8449;
    wire N__8448;
    wire N__8445;
    wire N__8440;
    wire N__8437;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8421;
    wire N__8418;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8388;
    wire N__8385;
    wire N__8382;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8355;
    wire N__8352;
    wire N__8349;
    wire N__8346;
    wire N__8343;
    wire N__8340;
    wire N__8337;
    wire VCCG0;
    wire bfn_1_2_0_;
    wire \POWERLED.mult1_un131_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_cry_3 ;
    wire \POWERLED.mult1_un131_sum_cry_4 ;
    wire \POWERLED.mult1_un131_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_cry_6 ;
    wire \POWERLED.mult1_un131_sum_cry_7 ;
    wire \POWERLED.mult1_un131_sum_s_8_cascade_ ;
    wire bfn_1_3_0_;
    wire \POWERLED.mult1_un138_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_cry_3_s ;
    wire \POWERLED.mult1_un138_sum_cry_3 ;
    wire \POWERLED.mult1_un131_sum_cry_4_s ;
    wire \POWERLED.mult1_un138_sum_cry_4 ;
    wire \POWERLED.mult1_un131_sum_cry_5_s ;
    wire \POWERLED.mult1_un138_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_cry_6_s ;
    wire \POWERLED.mult1_un131_sum_i_0_8 ;
    wire \POWERLED.mult1_un138_sum_cry_6 ;
    wire \POWERLED.mult1_un138_sum_axb_8 ;
    wire \POWERLED.mult1_un138_sum_cry_7 ;
    wire \POWERLED.mult1_un131_sum_s_8 ;
    wire bfn_1_5_0_;
    wire \POWERLED.mult1_un138_sum_i_0_8 ;
    wire \POWERLED.mult1_un145_sum_cry_2 ;
    wire \POWERLED.mult1_un138_sum_cry_3_s ;
    wire \POWERLED.mult1_un145_sum_axb_4_l_fx ;
    wire \POWERLED.mult1_un145_sum_cry_3 ;
    wire \POWERLED.mult1_un138_sum_cry_4_s ;
    wire \POWERLED.mult1_un145_sum_cry_4 ;
    wire \POWERLED.mult1_un138_sum_cry_5_s ;
    wire \POWERLED.mult1_un145_sum_cry_5 ;
    wire \POWERLED.mult1_un138_sum_cry_6_s ;
    wire \POWERLED.mult1_un145_sum_axb_7_l_fx ;
    wire \POWERLED.mult1_un145_sum_cry_6 ;
    wire \POWERLED.mult1_un145_sum_axb_8 ;
    wire \POWERLED.mult1_un145_sum_cry_7 ;
    wire bfn_1_6_0_;
    wire \POWERLED.mult1_un152_sum_cry_2 ;
    wire \POWERLED.mult1_un145_sum_cry_3_s ;
    wire \POWERLED.mult1_un152_sum_cry_3 ;
    wire \POWERLED.mult1_un145_sum_cry_4_s ;
    wire \POWERLED.mult1_un152_sum_cry_4 ;
    wire \POWERLED.mult1_un145_sum_cry_5_s ;
    wire \POWERLED.mult1_un152_sum_cry_5 ;
    wire \POWERLED.mult1_un145_sum_cry_6_s ;
    wire \POWERLED.mult1_un145_sum_i_0_8 ;
    wire \POWERLED.mult1_un152_sum_cry_6 ;
    wire \POWERLED.mult1_un152_sum_axb_8 ;
    wire \POWERLED.mult1_un152_sum_cry_7 ;
    wire \POWERLED.mult1_un152_sum_s_8_cascade_ ;
    wire bfn_1_7_0_;
    wire \POWERLED.mult1_un159_sum_cry_1 ;
    wire \POWERLED.mult1_un152_sum_cry_3_s ;
    wire \POWERLED.mult1_un159_sum_cry_2 ;
    wire \POWERLED.mult1_un152_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_cry_3 ;
    wire \POWERLED.mult1_un152_sum_cry_5_s ;
    wire \POWERLED.mult1_un159_sum_cry_4 ;
    wire \POWERLED.mult1_un152_sum_cry_6_s ;
    wire \POWERLED.mult1_un152_sum_i_0_8 ;
    wire \POWERLED.mult1_un159_sum_cry_5 ;
    wire \POWERLED.mult1_un159_sum_axb_7 ;
    wire \POWERLED.mult1_un159_sum_cry_6 ;
    wire \POWERLED.mult1_un159_sum_s_7_cascade_ ;
    wire \POWERLED.mult1_un145_sum_i ;
    wire bfn_1_10_0_;
    wire \RSMRST_PWRGD.un1_count_1_cry_0 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_1 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_2 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_3 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_4 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_5 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_6 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_7 ;
    wire bfn_1_11_0_;
    wire \RSMRST_PWRGD.un1_count_1_cry_8 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_9 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_10 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_11 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_12 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_13 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_1_12_0_;
    wire vpp_ok;
    wire vddq_en;
    wire bfn_2_2_0_;
    wire \POWERLED.mult1_un124_sum_cry_3_s ;
    wire \POWERLED.mult1_un124_sum_cry_2 ;
    wire \POWERLED.mult1_un124_sum_cry_4_s ;
    wire \POWERLED.mult1_un124_sum_cry_3 ;
    wire \POWERLED.mult1_un124_sum_cry_5_s ;
    wire \POWERLED.mult1_un124_sum_cry_4 ;
    wire \POWERLED.mult1_un124_sum_cry_6_s ;
    wire \POWERLED.mult1_un124_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_axb_8 ;
    wire \POWERLED.mult1_un124_sum_cry_6 ;
    wire \POWERLED.mult1_un124_sum_cry_7 ;
    wire \POWERLED.mult1_un124_sum_i_0_8 ;
    wire \POWERLED.mult1_un131_sum_i ;
    wire \POWERLED.mult1_un124_sum_i ;
    wire \POWERLED.mult1_un117_sum_i_0_8 ;
    wire \POWERLED.mult1_un117_sum_i ;
    wire \POWERLED.mult1_un124_sum_s_8 ;
    wire \POWERLED.mult1_un138_sum_s_8 ;
    wire \POWERLED.mult1_un145_sum_s_8 ;
    wire \POWERLED.count_i_0_0 ;
    wire bfn_2_5_0_;
    wire \POWERLED.un1_count_2_1 ;
    wire \POWERLED.count_i_1 ;
    wire \POWERLED.un1_count_2_cry_0 ;
    wire \POWERLED.count_i_2 ;
    wire \POWERLED.un1_count_2_cry_1 ;
    wire \POWERLED.un1_count_2_3 ;
    wire \POWERLED.count_i_3 ;
    wire \POWERLED.un1_count_2_cry_2 ;
    wire \POWERLED.un1_count_2_4 ;
    wire \POWERLED.count_i_4 ;
    wire \POWERLED.un1_count_2_cry_3 ;
    wire \POWERLED.un1_count_2_5 ;
    wire \POWERLED.count_i_5 ;
    wire \POWERLED.un1_count_2_cry_4 ;
    wire \POWERLED.un1_count_2_6 ;
    wire \POWERLED.count_i_6 ;
    wire \POWERLED.un1_count_2_cry_5 ;
    wire \POWERLED.count_i_7 ;
    wire \POWERLED.un1_count_2_cry_6 ;
    wire \POWERLED.un1_count_2_cry_7 ;
    wire \POWERLED.count_i_8 ;
    wire bfn_2_6_0_;
    wire \POWERLED.count_i_9 ;
    wire \POWERLED.un1_count_2_cry_8 ;
    wire \POWERLED.count_i_10 ;
    wire \POWERLED.un1_count_2_cry_9 ;
    wire \POWERLED.count_i_11 ;
    wire \POWERLED.un1_count_2_cry_10 ;
    wire \POWERLED.count_i_12 ;
    wire \POWERLED.un1_count_2_cry_11 ;
    wire \POWERLED.count_i_13 ;
    wire \POWERLED.un1_count_2_cry_12 ;
    wire \POWERLED.count_i_14 ;
    wire \POWERLED.un1_count_2_cry_13 ;
    wire \POWERLED.count_i_15 ;
    wire \POWERLED.un1_count_2_cry_14 ;
    wire \POWERLED.un1_count_2_cry_15 ;
    wire bfn_2_7_0_;
    wire \POWERLED.mult1_un138_sum_i ;
    wire slp_susn;
    wire v5a_ok;
    wire v33a_ok;
    wire v1p8a_ok;
    wire \POWERLED.mult1_un152_sum_i ;
    wire \POWERLED.mult1_un152_sum_s_8 ;
    wire \POWERLED.un1_count_2_2 ;
    wire \POWERLED.un1_count_2_12 ;
    wire \POWERLED.un1_count_2_cry_15_THRU_CO ;
    wire bfn_2_8_0_;
    wire \POWERLED.mult1_un166_sum_cry_0 ;
    wire \POWERLED.mult1_un159_sum_cry_2_s ;
    wire \POWERLED.mult1_un166_sum_cry_1 ;
    wire \POWERLED.mult1_un159_sum_cry_3_s ;
    wire \POWERLED.mult1_un166_sum_cry_2 ;
    wire \POWERLED.mult1_un159_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_s_7 ;
    wire \POWERLED.mult1_un166_sum_cry_3 ;
    wire \POWERLED.mult1_un159_sum_cry_5_s ;
    wire G_385;
    wire \POWERLED.mult1_un166_sum_cry_4 ;
    wire \POWERLED.mult1_un166_sum_axb_6 ;
    wire \POWERLED.mult1_un166_sum_cry_5 ;
    wire \POWERLED.un1_count_2_0 ;
    wire \POWERLED.mult1_un159_sum_i ;
    wire \RSMRST_PWRGD.N_37 ;
    wire \RSMRST_PWRGD.countZ0Z_7 ;
    wire \RSMRST_PWRGD.countZ0Z_3 ;
    wire \RSMRST_PWRGD.curr_stateZ0Z_1 ;
    wire \RSMRST_PWRGD.countZ0Z_4 ;
    wire \RSMRST_PWRGD.countZ0Z_1 ;
    wire \RSMRST_PWRGD.countZ0Z_5 ;
    wire \RSMRST_PWRGD.countZ0Z_2 ;
    wire \RSMRST_PWRGD.countZ0Z_10 ;
    wire \RSMRST_PWRGD.countZ0Z_11 ;
    wire \RSMRST_PWRGD.countZ0Z_13 ;
    wire \RSMRST_PWRGD.countZ0Z_6 ;
    wire \RSMRST_PWRGD.countZ0Z_15 ;
    wire \RSMRST_PWRGD.countZ0Z_14 ;
    wire \RSMRST_PWRGD.m4_i_i_a2_0_7 ;
    wire \RSMRST_PWRGD.countZ0Z_9 ;
    wire \RSMRST_PWRGD.countZ0Z_8 ;
    wire \RSMRST_PWRGD.countZ0Z_12 ;
    wire \RSMRST_PWRGD.countZ0Z_0 ;
    wire \RSMRST_PWRGD.m4_i_i_a2_0_10 ;
    wire \RSMRST_PWRGD.m4_i_i_a2_0_11 ;
    wire \RSMRST_PWRGD.m4_i_i_a2_0_9_cascade_ ;
    wire \RSMRST_PWRGD.m4_i_i_a2_0_12 ;
    wire \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0 ;
    wire \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0_cascade_ ;
    wire \RSMRST_PWRGD.N_49_2 ;
    wire v5s_enn;
    wire \RSMRST_PWRGD.N_241 ;
    wire \POWERLED.g0_0_4_cascade_ ;
    wire \POWERLED.un1_count_0 ;
    wire \POWERLED.un1_countlt6_0 ;
    wire \POWERLED.g0_0_5_cascade_ ;
    wire \POWERLED.g0_0_7 ;
    wire bfn_4_5_0_;
    wire \POWERLED.mult1_un117_sum_cry_3_s ;
    wire \POWERLED.mult1_un117_sum_cry_2 ;
    wire \POWERLED.mult1_un117_sum_cry_4_s ;
    wire \POWERLED.mult1_un117_sum_cry_3 ;
    wire \POWERLED.mult1_un117_sum_cry_5_s ;
    wire \POWERLED.mult1_un117_sum_cry_4 ;
    wire \POWERLED.mult1_un117_sum_cry_6_s ;
    wire \POWERLED.mult1_un117_sum_cry_5 ;
    wire \POWERLED.mult1_un124_sum_axb_8 ;
    wire \POWERLED.mult1_un117_sum_cry_6 ;
    wire \POWERLED.mult1_un117_sum_cry_7 ;
    wire \POWERLED.mult1_un117_sum_s_8 ;
    wire \POWERLED.mult1_un117_sum_s_8_cascade_ ;
    wire \POWERLED.un1_count_2_7 ;
    wire \POWERLED.un1_count_2_14 ;
    wire \POWERLED.un1_count_2_9 ;
    wire \POWERLED.un1_count_2_8 ;
    wire \POWERLED.mult1_un110_sum_i_0_8 ;
    wire \POWERLED.un1_count_2_13 ;
    wire \POWERLED.un1_count_2_10 ;
    wire \POWERLED.un1_count_2_11 ;
    wire \POWERLED.curr_state_0_0 ;
    wire pwrbtn_led;
    wire \POWERLED.pwm_out_RNOZ0 ;
    wire bfn_4_8_0_;
    wire \POWERLED.mult1_un54_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6 ;
    wire \POWERLED.mult1_un54_sum_cry_7 ;
    wire \POWERLED.un1_count_2_15 ;
    wire bfn_4_9_0_;
    wire \POWERLED.mult1_un47_sum_cry_3_s ;
    wire \POWERLED.mult1_un47_sum_cry_2 ;
    wire \POWERLED.mult1_un47_sum_cry_4_s ;
    wire \POWERLED.mult1_un47_sum_cry_3 ;
    wire \POWERLED.mult1_un47_sum_cry_5_s ;
    wire \POWERLED.mult1_un47_sum_cry_4 ;
    wire \POWERLED.mult1_un47_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_7_THRU_CO ;
    wire \POWERLED.mult1_un47_sum_cry_6 ;
    wire \POWERLED.mult1_un54_sum_s_8_cascade_ ;
    wire \POWERLED.un1_dutycycle_1_i_29 ;
    wire \POWERLED.un1_dutycycle_1_i_28 ;
    wire \POWERLED.mult1_un47_sum_axb_4 ;
    wire vccst_en_cascade_;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_5 ;
    wire \RSMRST_PWRGD.curr_stateZ0Z_0 ;
    wire \RSMRST_PWRGD.N_240 ;
    wire \VPP_VDDQ.un6_count_10 ;
    wire \VPP_VDDQ.un6_count_9_cascade_ ;
    wire \VPP_VDDQ.un6_count_8 ;
    wire \VPP_VDDQ.un6_count_11 ;
    wire \POWERLED.count_RNIOVT24Z0Z_11 ;
    wire \POWERLED.un1_countlto15_4 ;
    wire \POWERLED.un1_countlt6_cascade_ ;
    wire \POWERLED.un1_countlto15_5 ;
    wire \POWERLED.un1_countlto15_7 ;
    wire tmp_RNIRH3P;
    wire \POWERLED.mult1_un110_sum_i ;
    wire \COUNTER.tmp_i ;
    wire bfn_5_6_0_;
    wire \POWERLED.mult1_un110_sum_cry_3_s ;
    wire \POWERLED.mult1_un110_sum_cry_2 ;
    wire \POWERLED.mult1_un110_sum_cry_4_s ;
    wire \POWERLED.mult1_un110_sum_cry_3 ;
    wire \POWERLED.mult1_un110_sum_cry_5_s ;
    wire \POWERLED.mult1_un110_sum_cry_4 ;
    wire \POWERLED.mult1_un110_sum_cry_6_s ;
    wire \POWERLED.mult1_un110_sum_cry_5 ;
    wire \POWERLED.mult1_un117_sum_axb_8 ;
    wire \POWERLED.mult1_un110_sum_cry_6 ;
    wire \POWERLED.mult1_un110_sum_cry_7 ;
    wire \POWERLED.mult1_un110_sum_s_8 ;
    wire \POWERLED.mult1_un103_sum_i ;
    wire bfn_5_7_0_;
    wire \POWERLED.mult1_un96_sum_cry_2 ;
    wire \POWERLED.mult1_un96_sum_cry_3 ;
    wire \POWERLED.mult1_un96_sum_cry_4 ;
    wire \POWERLED.mult1_un96_sum_cry_5 ;
    wire \POWERLED.mult1_un96_sum_cry_6 ;
    wire \POWERLED.mult1_un96_sum_cry_7 ;
    wire \POWERLED.mult1_un96_sum_s_8_cascade_ ;
    wire bfn_5_8_0_;
    wire \POWERLED.mult1_un54_sum_i ;
    wire \POWERLED.mult1_un61_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3_s ;
    wire \POWERLED.mult1_un61_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4_s ;
    wire \POWERLED.mult1_un61_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_cry_5_s ;
    wire \POWERLED.mult1_un61_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6_s ;
    wire \POWERLED.mult1_un54_sum_i_8 ;
    wire \POWERLED.mult1_un61_sum_cry_6 ;
    wire \POWERLED.mult1_un47_sum_cry_6_s ;
    wire \POWERLED.mult1_un54_sum_s_8 ;
    wire \POWERLED.mult1_un54_sum_cry_6_THRU_CO ;
    wire \POWERLED.mult1_un61_sum_cry_7 ;
    wire \POWERLED.mult1_un61_sum_s_8_cascade_ ;
    wire bfn_5_9_0_;
    wire \POWERLED.mult1_un61_sum_i ;
    wire \POWERLED.mult1_un68_sum_cry_2 ;
    wire \POWERLED.mult1_un61_sum_cry_3_s ;
    wire \POWERLED.mult1_un68_sum_cry_3 ;
    wire \POWERLED.mult1_un61_sum_cry_4_s ;
    wire \POWERLED.mult1_un68_sum_cry_4 ;
    wire \POWERLED.mult1_un61_sum_s_8 ;
    wire \POWERLED.mult1_un61_sum_cry_5_s ;
    wire \POWERLED.mult1_un68_sum_cry_5 ;
    wire \POWERLED.mult1_un61_sum_cry_6_s ;
    wire \POWERLED.mult1_un61_sum_i_0_8 ;
    wire \POWERLED.mult1_un68_sum_cry_6 ;
    wire \POWERLED.mult1_un68_sum_axb_8 ;
    wire \POWERLED.mult1_un68_sum_cry_7 ;
    wire \POWERLED.mult1_un68_sum_s_8_cascade_ ;
    wire \POWERLED.un1_dutycycle_1_axb_0 ;
    wire bfn_5_10_0_;
    wire \POWERLED.mult1_un138_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_0 ;
    wire \POWERLED.mult1_un131_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_1 ;
    wire \POWERLED.mult1_un124_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_2 ;
    wire \POWERLED.mult1_un117_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_3 ;
    wire \POWERLED.mult1_un110_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_4 ;
    wire \POWERLED.un1_dutycycle_1_cry_5 ;
    wire \POWERLED.un1_dutycycle_1_cry_6 ;
    wire \POWERLED.un1_dutycycle_1_cry_7 ;
    wire bfn_5_11_0_;
    wire \POWERLED.un1_dutycycle_1_cry_8 ;
    wire \POWERLED.un1_dutycycle_1_cry_9 ;
    wire \POWERLED.un1_dutycycle_1_cry_10 ;
    wire \POWERLED.mult1_un61_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_11 ;
    wire \POWERLED.mult1_un54_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_12 ;
    wire \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1 ;
    wire \POWERLED.un1_dutycycle_1_cry_13 ;
    wire \POWERLED.un1_dutycycle_1_cry_14 ;
    wire \POWERLED.un1_dutycycle_1_cry_15 ;
    wire bfn_5_12_0_;
    wire \POWERLED.CO2 ;
    wire \POWERLED.CO2_THRU_CO ;
    wire \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1 ;
    wire \POWERLED.CO2_THRU_CO_cascade_ ;
    wire \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_4 ;
    wire \VPP_VDDQ.countZ0Z_0 ;
    wire bfn_5_13_0_;
    wire \VPP_VDDQ.countZ0Z_1 ;
    wire \VPP_VDDQ.un1_count_1_cry_0 ;
    wire \VPP_VDDQ.countZ0Z_2 ;
    wire \VPP_VDDQ.un1_count_1_cry_1 ;
    wire \VPP_VDDQ.countZ0Z_3 ;
    wire \VPP_VDDQ.un1_count_1_cry_2 ;
    wire \VPP_VDDQ.countZ0Z_4 ;
    wire \VPP_VDDQ.un1_count_1_cry_3 ;
    wire \VPP_VDDQ.countZ0Z_5 ;
    wire \VPP_VDDQ.un1_count_1_cry_4 ;
    wire \VPP_VDDQ.countZ0Z_6 ;
    wire \VPP_VDDQ.un1_count_1_cry_5 ;
    wire \VPP_VDDQ.countZ0Z_7 ;
    wire \VPP_VDDQ.un1_count_1_cry_6 ;
    wire \VPP_VDDQ.un1_count_1_cry_7 ;
    wire \VPP_VDDQ.countZ0Z_8 ;
    wire bfn_5_14_0_;
    wire \VPP_VDDQ.countZ0Z_9 ;
    wire \VPP_VDDQ.un1_count_1_cry_8 ;
    wire \VPP_VDDQ.countZ0Z_10 ;
    wire \VPP_VDDQ.un1_count_1_cry_9 ;
    wire \VPP_VDDQ.countZ0Z_11 ;
    wire \VPP_VDDQ.un1_count_1_cry_10 ;
    wire \VPP_VDDQ.countZ0Z_12 ;
    wire \VPP_VDDQ.un1_count_1_cry_11 ;
    wire \VPP_VDDQ.countZ0Z_13 ;
    wire \VPP_VDDQ.un1_count_1_cry_12 ;
    wire \VPP_VDDQ.countZ0Z_14 ;
    wire \VPP_VDDQ.un1_count_1_cry_13 ;
    wire \VPP_VDDQ.un1_count_1_cry_14 ;
    wire \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_5_15_0_;
    wire \VPP_VDDQ.countZ0Z_15 ;
    wire \POWERLED.countZ0Z_1 ;
    wire \POWERLED.countZ0Z_0 ;
    wire bfn_6_3_0_;
    wire \POWERLED.countZ0Z_2 ;
    wire \POWERLED.un1_count_1_cry_1 ;
    wire \POWERLED.countZ0Z_3 ;
    wire \POWERLED.un1_count_1_cry_2 ;
    wire \POWERLED.countZ0Z_4 ;
    wire \POWERLED.un1_count_1_cry_3 ;
    wire \POWERLED.countZ0Z_5 ;
    wire \POWERLED.un1_count_1_cry_4 ;
    wire \POWERLED.countZ0Z_6 ;
    wire \POWERLED.un1_count_1_cry_5 ;
    wire \POWERLED.countZ0Z_7 ;
    wire \POWERLED.un1_count_1_cry_6 ;
    wire \POWERLED.countZ0Z_8 ;
    wire \POWERLED.un1_count_1_cry_7 ;
    wire \POWERLED.un1_count_1_cry_8 ;
    wire \POWERLED.countZ0Z_9 ;
    wire bfn_6_4_0_;
    wire \POWERLED.countZ0Z_10 ;
    wire \POWERLED.un1_count_1_cry_9 ;
    wire \POWERLED.countZ0Z_11 ;
    wire \POWERLED.un1_count_1_cry_10 ;
    wire \POWERLED.countZ0Z_12 ;
    wire \POWERLED.un1_count_1_cry_11 ;
    wire \POWERLED.countZ0Z_13 ;
    wire \POWERLED.un1_count_1_cry_12 ;
    wire \POWERLED.countZ0Z_14 ;
    wire \POWERLED.un1_count_1_cry_13 ;
    wire \POWERLED.un1_count_1_cry_14 ;
    wire \POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire \POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO ;
    wire bfn_6_5_0_;
    wire \POWERLED.countZ0Z_15 ;
    wire \POWERLED.N_49_5 ;
    wire \POWERLED.curr_state_RNI75RB5Z0Z_0 ;
    wire \POWERLED.mult1_un103_sum ;
    wire bfn_6_6_0_;
    wire \POWERLED.mult1_un103_sum_cry_3_s ;
    wire \POWERLED.mult1_un103_sum_cry_2 ;
    wire \POWERLED.mult1_un96_sum_cry_3_s ;
    wire \POWERLED.mult1_un103_sum_cry_4_s ;
    wire \POWERLED.mult1_un103_sum_cry_3 ;
    wire \POWERLED.mult1_un96_sum_cry_4_s ;
    wire \POWERLED.mult1_un103_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_cry_4 ;
    wire \POWERLED.mult1_un96_sum_s_8 ;
    wire \POWERLED.mult1_un96_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_cry_6_s ;
    wire \POWERLED.mult1_un103_sum_cry_5 ;
    wire \POWERLED.mult1_un96_sum_cry_6_s ;
    wire \POWERLED.mult1_un96_sum_i_0_8 ;
    wire \POWERLED.mult1_un110_sum_axb_8 ;
    wire \POWERLED.mult1_un103_sum_cry_6 ;
    wire \POWERLED.mult1_un103_sum_axb_8 ;
    wire \POWERLED.mult1_un103_sum_cry_7 ;
    wire \POWERLED.mult1_un103_sum_s_8 ;
    wire \POWERLED.mult1_un103_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un103_sum_i_0_8 ;
    wire bfn_6_7_0_;
    wire \POWERLED.mult1_un89_sum_cry_3_s ;
    wire \POWERLED.mult1_un89_sum_cry_2 ;
    wire \POWERLED.mult1_un89_sum_cry_4_s ;
    wire \POWERLED.mult1_un89_sum_cry_3 ;
    wire \POWERLED.mult1_un89_sum_cry_5_s ;
    wire \POWERLED.mult1_un89_sum_cry_4 ;
    wire \POWERLED.mult1_un89_sum_cry_6_s ;
    wire \POWERLED.mult1_un89_sum_cry_5 ;
    wire \POWERLED.mult1_un96_sum_axb_8 ;
    wire \POWERLED.mult1_un89_sum_cry_6 ;
    wire \POWERLED.mult1_un89_sum_cry_7 ;
    wire \POWERLED.mult1_un89_sum_s_8 ;
    wire \POWERLED.mult1_un89_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un89_sum_i_0_8 ;
    wire bfn_6_8_0_;
    wire \POWERLED.mult1_un75_sum_i ;
    wire \POWERLED.mult1_un82_sum_cry_3_s ;
    wire \POWERLED.mult1_un82_sum_cry_2 ;
    wire \POWERLED.mult1_un82_sum_cry_4_s ;
    wire \POWERLED.mult1_un82_sum_cry_3 ;
    wire \POWERLED.mult1_un82_sum_cry_5_s ;
    wire \POWERLED.mult1_un82_sum_cry_4 ;
    wire \POWERLED.mult1_un82_sum_cry_6_s ;
    wire \POWERLED.mult1_un82_sum_cry_5 ;
    wire \POWERLED.mult1_un89_sum_axb_8 ;
    wire \POWERLED.mult1_un82_sum_cry_6 ;
    wire \POWERLED.mult1_un82_sum_cry_7 ;
    wire \POWERLED.mult1_un82_sum_s_8 ;
    wire \POWERLED.mult1_un82_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un82_sum_i_0_8 ;
    wire \POWERLED.mult1_un75_sum ;
    wire bfn_6_9_0_;
    wire \POWERLED.mult1_un75_sum_cry_3_s ;
    wire \POWERLED.mult1_un75_sum_cry_2 ;
    wire \POWERLED.mult1_un68_sum_cry_3_s ;
    wire \POWERLED.mult1_un75_sum_cry_4_s ;
    wire \POWERLED.mult1_un75_sum_cry_3 ;
    wire \POWERLED.mult1_un68_sum_cry_4_s ;
    wire \POWERLED.mult1_un75_sum_cry_5_s ;
    wire \POWERLED.mult1_un75_sum_cry_4 ;
    wire \POWERLED.mult1_un68_sum_s_8 ;
    wire \POWERLED.mult1_un68_sum_cry_5_s ;
    wire \POWERLED.mult1_un75_sum_cry_6_s ;
    wire \POWERLED.mult1_un75_sum_cry_5 ;
    wire \POWERLED.mult1_un68_sum_cry_6_s ;
    wire \POWERLED.mult1_un68_sum_i_0_8 ;
    wire \POWERLED.mult1_un82_sum_axb_8 ;
    wire \POWERLED.mult1_un75_sum_cry_6 ;
    wire \POWERLED.mult1_un75_sum_axb_8 ;
    wire \POWERLED.mult1_un75_sum_cry_7 ;
    wire \POWERLED.mult1_un75_sum_s_8 ;
    wire \POWERLED.mult1_un75_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un75_sum_i_0_8 ;
    wire \POWERLED.dutycycle_RNIJL1R1Z0Z_6 ;
    wire \POWERLED.un1_dutycycle_1_19_0_cascade_ ;
    wire \POWERLED.dutycycle_RNIEJ021Z0Z_4 ;
    wire \POWERLED.dutycycle_RNIQAI81Z0Z_4 ;
    wire \POWERLED.mult1_un68_sum ;
    wire \POWERLED.mult1_un68_sum_i ;
    wire \POWERLED.dutycycle_RNI53MGZ0Z_14 ;
    wire \POWERLED.dutycycle_RNIJNBA1Z0Z_6 ;
    wire \POWERLED.dutycycle_RNIOQLJZ0Z_4 ;
    wire \POWERLED.un1_dutycycle_1_34_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_1_axb_8 ;
    wire \POWERLED.dutycycle_RNIB1FLZ0Z_8 ;
    wire \POWERLED.dutycycle_fast_RNILMLMZ0Z_6 ;
    wire \POWERLED.dutycycle_RNI84C11Z0Z_14 ;
    wire \POWERLED.dutycycle_RNIQ09G1Z0Z_10 ;
    wire \POWERLED.un1_dutycycle_1_39_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI34C41Z0Z_8 ;
    wire \POWERLED.dutycycle_RNI73C11Z0Z_15 ;
    wire \POWERLED.dutycycle_RNIE4FLZ0Z_9 ;
    wire \POWERLED.dutycycle_RNI2V0PZ0Z_10 ;
    wire \POWERLED.dutycycle_RNI2V0PZ0Z_10_cascade_ ;
    wire \POWERLED.dutycycle_RNI712I1Z0Z_15 ;
    wire \POWERLED.dutycycle_RNIO18NZ0Z_9 ;
    wire \POWERLED.dutycycle_RNIC8C11Z0Z_15 ;
    wire \POWERLED.dutycycle_RNI31MGZ0Z_12 ;
    wire \POWERLED.dutycycle_RNI31MG_0Z0Z_12 ;
    wire \POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI75MGZ0Z_15 ;
    wire \VPP_VDDQ.N_108_i ;
    wire \VPP_VDDQ.N_242_cascade_ ;
    wire N_154_cascade_;
    wire N_128;
    wire N_128_cascade_;
    wire \VPP_VDDQ.delayed_vddq_pwrgd_0 ;
    wire G_111;
    wire \VPP_VDDQ.N_49_1 ;
    wire \PCH_PWRGD.N_3_i_cascade_ ;
    wire \PCH_PWRGD.un1_curr_state_0_sqmuxa_0_cascade_ ;
    wire vr_ready_vccin;
    wire \PCH_PWRGD.curr_stateZ0Z_1 ;
    wire \PCH_PWRGD.N_3_i ;
    wire \PCH_PWRGD.curr_stateZ0Z_0 ;
    wire pch_pwrok;
    wire \POWERLED.mult1_un96_sum ;
    wire \POWERLED.mult1_un96_sum_i ;
    wire \POWERLED.mult1_un89_sum ;
    wire \POWERLED.mult1_un89_sum_i ;
    wire \POWERLED.N_117 ;
    wire \POWERLED.N_117_cascade_ ;
    wire \POWERLED.mult1_un82_sum ;
    wire \POWERLED.mult1_un82_sum_i ;
    wire \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5 ;
    wire \POWERLED.dutycycle_RNI6NI81Z0Z_5 ;
    wire \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5 ;
    wire \POWERLED.dutycycle_RNIK4I81Z0Z_6 ;
    wire \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6 ;
    wire \POWERLED.dutycycle_fastZ0Z_6 ;
    wire \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6 ;
    wire \POWERLED.dutycycle ;
    wire bfn_7_11_0_;
    wire \POWERLED.dutycycle_cry_c_0_THRU_CO ;
    wire \POWERLED.dutycycle_cry_0 ;
    wire \POWERLED.dutycycle_s_2 ;
    wire \POWERLED.dutycycle_cry_1 ;
    wire \POWERLED.dutycycle_cry_2 ;
    wire \POWERLED.dutycycle_cry_3 ;
    wire \POWERLED.dutycycle_cry_4 ;
    wire \POWERLED.dutycycleZ0Z_6 ;
    wire \POWERLED.dutycycle_s_6 ;
    wire \POWERLED.dutycycle_cry_5 ;
    wire \POWERLED.dutycycle_cry_6 ;
    wire bfn_7_12_0_;
    wire \POWERLED.dutycycle_cry_7 ;
    wire \POWERLED.dutycycle_cry_8 ;
    wire \POWERLED.dutycycle_cry_9 ;
    wire \POWERLED.dutycycle_cry_10 ;
    wire \POWERLED.dutycycle_cry_11 ;
    wire \POWERLED.dutycycle_cry_12 ;
    wire \POWERLED.dutycycle_cry_13 ;
    wire \POWERLED.dutycycle_cry_14 ;
    wire bfn_7_13_0_;
    wire \VPP_VDDQ.count_esr_RNIRFM64Z0Z_15 ;
    wire \VPP_VDDQ.curr_stateZ0Z_1 ;
    wire VPP_VDDQ_curr_state_0;
    wire \PCH_PWRGD.un1_curr_state10_0 ;
    wire bfn_8_1_0_;
    wire \PCH_PWRGD.un1_count_1_cry_0 ;
    wire \PCH_PWRGD.un1_count_1_cry_1 ;
    wire \PCH_PWRGD.un1_count_1_cry_2 ;
    wire \PCH_PWRGD.un1_count_1_cry_3 ;
    wire \PCH_PWRGD.un1_count_1_cry_4 ;
    wire \PCH_PWRGD.un1_count_1_cry_5 ;
    wire \PCH_PWRGD.un1_count_1_cry_6 ;
    wire \PCH_PWRGD.un1_count_1_cry_7 ;
    wire bfn_8_2_0_;
    wire \PCH_PWRGD.un1_count_1_cry_8 ;
    wire \PCH_PWRGD.un1_count_1_cry_9 ;
    wire \PCH_PWRGD.un1_count_1_cry_10 ;
    wire \PCH_PWRGD.un1_count_1_cry_11 ;
    wire \PCH_PWRGD.un1_count_1_cry_12 ;
    wire \PCH_PWRGD.un1_count_1_cry_13 ;
    wire \PCH_PWRGD.un1_count_1_cry_14 ;
    wire \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_8_3_0_;
    wire \PCH_PWRGD.N_49_3 ;
    wire \PCH_PWRGD.curr_state_RNI7N705Z0Z_0 ;
    wire bfn_8_5_0_;
    wire \COUNTER.counterZ0Z_2 ;
    wire \COUNTER.counter_1_cry_1_THRU_CO ;
    wire \COUNTER.counter_1_cry_1 ;
    wire \COUNTER.counterZ0Z_3 ;
    wire \COUNTER.counter_1_cry_2_THRU_CO ;
    wire \COUNTER.counter_1_cry_2 ;
    wire \COUNTER.counterZ0Z_4 ;
    wire \COUNTER.counter_1_cry_3_THRU_CO ;
    wire \COUNTER.counter_1_cry_3 ;
    wire \COUNTER.counter_1_cry_4 ;
    wire \COUNTER.counter_1_cry_5 ;
    wire \COUNTER.counter_1_cry_6 ;
    wire \COUNTER.counter_1_cry_7 ;
    wire \COUNTER.counter_1_cry_8 ;
    wire bfn_8_6_0_;
    wire \COUNTER.counter_1_cry_9 ;
    wire \COUNTER.counter_1_cry_10 ;
    wire \COUNTER.counter_1_cry_11 ;
    wire \COUNTER.counter_1_cry_12 ;
    wire \COUNTER.counter_1_cry_13 ;
    wire \COUNTER.counter_1_cry_14 ;
    wire \COUNTER.counter_1_cry_15 ;
    wire \COUNTER.counter_1_cry_16 ;
    wire bfn_8_7_0_;
    wire \COUNTER.counter_1_cry_17 ;
    wire \COUNTER.counter_1_cry_18 ;
    wire \COUNTER.counter_1_cry_19 ;
    wire \COUNTER.counter_1_cry_20 ;
    wire \COUNTER.counter_1_cry_21 ;
    wire \COUNTER.counter_1_cry_22 ;
    wire \COUNTER.counter_1_cry_23 ;
    wire \COUNTER.counter_1_cry_24 ;
    wire bfn_8_8_0_;
    wire \COUNTER.counter_1_cry_25 ;
    wire \COUNTER.counter_1_cry_26 ;
    wire \COUNTER.counter_1_cry_27 ;
    wire \COUNTER.counter_1_cry_28 ;
    wire \COUNTER.counter_1_cry_29 ;
    wire \COUNTER.counter_1_cry_30 ;
    wire \COUNTER.counterZ0Z_30 ;
    wire \COUNTER.counterZ0Z_29 ;
    wire \COUNTER.counterZ0Z_31 ;
    wire \COUNTER.counterZ0Z_28 ;
    wire \POWERLED.N_234 ;
    wire \POWERLED.N_248_cascade_ ;
    wire \POWERLED.N_118 ;
    wire \POWERLED.dutycycle_RNIFHLJZ0Z_0 ;
    wire \POWERLED.dutycycleZ0Z_5 ;
    wire \POWERLED.dutycycle_RNIFHLJZ0Z_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI16B71Z0Z_5 ;
    wire \POWERLED.dutycycle_s_1 ;
    wire \POWERLED.dutycycleZ0Z_1 ;
    wire \POWERLED.un1_dutycycle_1_axb_1 ;
    wire \POWERLED.N_53 ;
    wire \POWERLED.dutycycle_s_0 ;
    wire \POWERLED.dutycycleZ0Z_0 ;
    wire \POWERLED.dutycycle_s_5 ;
    wire \POWERLED.un1_dutycycle_4_sqmuxa_0 ;
    wire \POWERLED.N_213 ;
    wire \POWERLED.dutycycle_fastZ0Z_5 ;
    wire \POWERLED.dutycycleZ0Z_4 ;
    wire \POWERLED.dutycycleZ0Z_15 ;
    wire \POWERLED.dutycycleZ0Z_7 ;
    wire \POWERLED.dutycycleZ0Z_3 ;
    wire \POWERLED.dutycycleZ0Z_2 ;
    wire \POWERLED.dutycycleZ0Z_14 ;
    wire \POWERLED.dutycycleZ0Z_13 ;
    wire \POWERLED.dutycycleZ0Z_12 ;
    wire \POWERLED.un1_dutycycle_1_44_0_cascade_ ;
    wire \POWERLED.dutycycle_RNIF3561Z0Z_9 ;
    wire \POWERLED.dutycycleZ0Z_10 ;
    wire \POWERLED.dutycycleZ0Z_11 ;
    wire \POWERLED.dutycycleZ0Z_9 ;
    wire \POWERLED.dutycycleZ0Z_8 ;
    wire \POWERLED.un2_slp_s3n_2_0_o2_3_7 ;
    wire \POWERLED.un2_slp_s3n_2_0_o2_3_8_cascade_ ;
    wire \POWERLED.un2_slp_s3n_2_0_o2_3_6 ;
    wire \POWERLED.N_112 ;
    wire \POWERLED.N_177_5_cascade_ ;
    wire \POWERLED.N_177_5 ;
    wire \POWERLED.N_368_0_i_i_a6_0_cascade_ ;
    wire \POWERLED.N_177 ;
    wire rsmrstn;
    wire \POWERLED.count_clk_0_sqmuxa_5_0_o2_0_0_cascade_ ;
    wire \POWERLED.N_141_cascade_ ;
    wire \POWERLED.count_clk_1_sqmuxa_5_i ;
    wire bfn_8_13_0_;
    wire \POWERLED.un1_count_clk_1_cry_0 ;
    wire \POWERLED.count_clkZ0Z_2 ;
    wire \POWERLED.un1_count_clk_1_cry_1 ;
    wire \POWERLED.count_clkZ0Z_3 ;
    wire \POWERLED.un1_count_clk_1_cry_2 ;
    wire \POWERLED.count_clkZ0Z_4 ;
    wire \POWERLED.un1_count_clk_1_cry_3 ;
    wire \POWERLED.un1_count_clk_1_cry_4 ;
    wire \POWERLED.count_clkZ0Z_6 ;
    wire \POWERLED.un1_count_clk_1_cry_5 ;
    wire \POWERLED.un1_count_clk_1_cry_6 ;
    wire \POWERLED.un1_count_clk_1_cry_7 ;
    wire \POWERLED.count_clkZ0Z_8 ;
    wire bfn_8_14_0_;
    wire \POWERLED.un1_count_clk_1_cry_8 ;
    wire \POWERLED.un1_count_clk_1_cry_9 ;
    wire \POWERLED.un1_count_clk_1_cry_10 ;
    wire \POWERLED.un1_count_clk_1_cry_11 ;
    wire \POWERLED.un1_count_clk_1_cry_12 ;
    wire \POWERLED.un1_count_clk_1_cry_13 ;
    wire \POWERLED.un1_count_clk_1_cry_14 ;
    wire \POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_8_15_0_;
    wire \PCH_PWRGD.countZ0Z_6 ;
    wire \PCH_PWRGD.countZ0Z_1 ;
    wire \PCH_PWRGD.countZ0Z_10 ;
    wire \PCH_PWRGD.countZ0Z_2 ;
    wire \PCH_PWRGD.un4_count_9_cascade_ ;
    wire \PCH_PWRGD.N_1_i ;
    wire \PCH_PWRGD.countZ0Z_5 ;
    wire \PCH_PWRGD.countZ0Z_4 ;
    wire \PCH_PWRGD.countZ0Z_7 ;
    wire \PCH_PWRGD.countZ0Z_3 ;
    wire \PCH_PWRGD.un4_count_11 ;
    wire \PCH_PWRGD.countZ0Z_9 ;
    wire \PCH_PWRGD.countZ0Z_8 ;
    wire \PCH_PWRGD.countZ0Z_11 ;
    wire \PCH_PWRGD.countZ0Z_0 ;
    wire \PCH_PWRGD.un4_count_10 ;
    wire \PCH_PWRGD.countZ0Z_14 ;
    wire \PCH_PWRGD.countZ0Z_13 ;
    wire \PCH_PWRGD.countZ0Z_12 ;
    wire \PCH_PWRGD.countZ0Z_15 ;
    wire \PCH_PWRGD.un4_count_8 ;
    wire \COUNTER.un4_counter_0_and ;
    wire bfn_9_4_0_;
    wire \COUNTER.un4_counter_0 ;
    wire \COUNTER.un4_counter_1 ;
    wire \COUNTER.un4_counter_2 ;
    wire \COUNTER.un4_counter_3 ;
    wire \COUNTER.un4_counter_4 ;
    wire \COUNTER.un4_counter_5 ;
    wire \COUNTER.un4_counter_7_and ;
    wire \COUNTER.un4_counter_6 ;
    wire \COUNTER.un4_counter_7 ;
    wire bfn_9_5_0_;
    wire \COUNTER.un4_counter_7_THRU_CO_cascade_ ;
    wire \COUNTER.counter_1_cry_5_THRU_CO ;
    wire \COUNTER.counter_1_cry_4_THRU_CO ;
    wire \COUNTER.un4_counter_7_THRU_CO ;
    wire \COUNTER.counterZ0Z_0 ;
    wire \COUNTER.counterZ0Z_6 ;
    wire \COUNTER.counterZ0Z_5 ;
    wire \COUNTER.counterZ0Z_7 ;
    wire \COUNTER.counterZ0Z_1 ;
    wire \COUNTER.un4_counter_1_and ;
    wire \COUNTER.counterZ0Z_18 ;
    wire \COUNTER.counterZ0Z_17 ;
    wire \COUNTER.counterZ0Z_19 ;
    wire \COUNTER.counterZ0Z_16 ;
    wire \COUNTER.un4_counter_4_and ;
    wire \COUNTER.counterZ0Z_10 ;
    wire \COUNTER.counterZ0Z_9 ;
    wire \COUNTER.counterZ0Z_11 ;
    wire \COUNTER.counterZ0Z_8 ;
    wire \COUNTER.un4_counter_2_and ;
    wire \COUNTER.counterZ0Z_14 ;
    wire \COUNTER.counterZ0Z_13 ;
    wire \COUNTER.counterZ0Z_15 ;
    wire \COUNTER.counterZ0Z_12 ;
    wire \COUNTER.un4_counter_3_and ;
    wire \COUNTER.counterZ0Z_26 ;
    wire \COUNTER.counterZ0Z_25 ;
    wire \COUNTER.counterZ0Z_27 ;
    wire \COUNTER.counterZ0Z_24 ;
    wire \COUNTER.un4_counter_6_and ;
    wire \COUNTER.counterZ0Z_22 ;
    wire \COUNTER.counterZ0Z_21 ;
    wire \COUNTER.counterZ0Z_23 ;
    wire \COUNTER.counterZ0Z_20 ;
    wire \COUNTER.un4_counter_5_and ;
    wire \POWERLED.N_214 ;
    wire \POWERLED.N_250 ;
    wire \POWERLED.N_178 ;
    wire \POWERLED.N_148_cascade_ ;
    wire \POWERLED.N_208_cascade_ ;
    wire \POWERLED.func_state_ns_i_0_1_1 ;
    wire \POWERLED.N_228 ;
    wire \POWERLED.func_state_ns_i_0_0_1 ;
    wire \POWERLED.N_248 ;
    wire \POWERLED.N_127 ;
    wire \POWERLED.N_179 ;
    wire \POWERLED.N_211 ;
    wire \POWERLED.func_stateZ0Z_0 ;
    wire \POWERLED.N_88_cascade_ ;
    wire \POWERLED.dutycycle_3_sqmuxa_1_i_0_1_1_cascade_ ;
    wire \POWERLED.N_366_1 ;
    wire \POWERLED.count_clk_1_sqmuxa_5_0_2 ;
    wire slp_s3n;
    wire slp_s4n;
    wire \POWERLED.dutycycle_lm_0_1_2 ;
    wire \POWERLED.N_88 ;
    wire \POWERLED.N_205_cascade_ ;
    wire \POWERLED.N_203_4 ;
    wire \POWERLED.count_clk_0_sqmuxa_5_0_a6_3_cascade_ ;
    wire \POWERLED.N_226 ;
    wire \POWERLED.N_200_2 ;
    wire \POWERLED.N_217 ;
    wire \POWERLED.func_stateZ0Z_1 ;
    wire \POWERLED.N_141 ;
    wire \POWERLED.N_149 ;
    wire \POWERLED.N_222 ;
    wire \POWERLED.N_149_cascade_ ;
    wire \POWERLED.N_207 ;
    wire \POWERLED.count_off_1_sqmuxa_i_a6_0_3 ;
    wire gpio_fpga_soc_4;
    wire \POWERLED.count_off_1_sqmuxa_i_a6_0_1 ;
    wire \POWERLED.N_243 ;
    wire vccst_en;
    wire \POWERLED.un2_slp_s3n_2_0_a6_3_0_cascade_ ;
    wire \POWERLED.un2_slp_s3n_2_0_1_0 ;
    wire \POWERLED.un2_slp_s3n_2_0_1_cascade_ ;
    wire \POWERLED.N_251 ;
    wire \POWERLED.count_clkZ0Z_7 ;
    wire \POWERLED.count_clk_0_sqmuxa_5_0_a6_1 ;
    wire \POWERLED.count_clkZ0Z_5 ;
    wire \POWERLED.count_clkZ0Z_9 ;
    wire \POWERLED.count_clkZ0Z_1 ;
    wire \POWERLED.N_146 ;
    wire \VPP_VDDQ.N_238 ;
    wire \POWERLED.count_clk_137_tz_0 ;
    wire \POWERLED.un2_slp_s3n_2_0 ;
    wire \POWERLED.count_clkZ0Z_11 ;
    wire \POWERLED.count_clkZ0Z_10 ;
    wire \POWERLED.count_clkZ0Z_12 ;
    wire \POWERLED.count_clkZ0Z_0 ;
    wire \POWERLED.count_clkZ0Z_15 ;
    wire \POWERLED.count_clkZ0Z_14 ;
    wire \POWERLED.count_clk_0_sqmuxa_5_0_o2_4_cascade_ ;
    wire \POWERLED.count_clkZ0Z_13 ;
    wire \POWERLED.N_136 ;
    wire \POWERLED.count_clk_RNIOH1J11Z0Z_7 ;
    wire \POWERLED.N_49_0 ;
    wire vccst_pwrgd;
    wire \ALL_SYS_PWRGD.N_186 ;
    wire \ALL_SYS_PWRGD.N_247 ;
    wire \ALL_SYS_PWRGD.N_186_cascade_ ;
    wire bfn_11_7_0_;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_0 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_1 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_2 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_3 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_4 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_5 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_6 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_7 ;
    wire bfn_11_8_0_;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_8 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_9 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_10 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_11 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_12 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_13 ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_14 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_11_9_0_;
    wire bfn_11_10_0_;
    wire \POWERLED.un1_count_off_1_cry_0 ;
    wire \POWERLED.un1_count_off_1_cry_1 ;
    wire \POWERLED.un1_count_off_1_cry_2 ;
    wire \POWERLED.un1_count_off_1_cry_3 ;
    wire \POWERLED.un1_count_off_1_cry_4 ;
    wire \POWERLED.un1_count_off_1_cry_5 ;
    wire \POWERLED.un1_count_off_1_cry_6 ;
    wire \POWERLED.un1_count_off_1_cry_7 ;
    wire bfn_11_11_0_;
    wire \POWERLED.un1_count_off_1_cry_8 ;
    wire \POWERLED.un1_count_off_1_cry_9 ;
    wire \POWERLED.un1_count_off_1_cry_10 ;
    wire \POWERLED.un1_count_off_1_cry_11 ;
    wire \POWERLED.un1_count_off_1_cry_12 ;
    wire \POWERLED.un1_count_off_1_cry_13 ;
    wire \POWERLED.un1_count_off_1_cry_14 ;
    wire \POWERLED.count_offZ0Z_4 ;
    wire \POWERLED.count_offZ0Z_7 ;
    wire \POWERLED.count_offZ0Z_3 ;
    wire \POWERLED.func_state_ns_0_a2_8_0_cascade_ ;
    wire \POWERLED.count_off_RNIIKVR3Z0Z_10 ;
    wire \POWERLED.count_offZ0Z_9 ;
    wire \POWERLED.count_offZ0Z_8 ;
    wire \POWERLED.func_state_ns_0_a2_9_0 ;
    wire \POWERLED.count_offZ0Z_10 ;
    wire \POWERLED.count_offZ0Z_14 ;
    wire \POWERLED.count_offZ0Z_11 ;
    wire \POWERLED.func_state_ns_0_a2_10_0 ;
    wire \POWERLED.count_offZ0Z_13 ;
    wire \POWERLED.count_offZ0Z_12 ;
    wire \POWERLED.count_offZ0Z_15 ;
    wire \POWERLED.count_offZ0Z_1 ;
    wire \POWERLED.func_state_ns_0_a2_11_0 ;
    wire \VPP_VDDQ.delayed_vddq_pwrgdZ0 ;
    wire N_55;
    wire vpp_en;
    wire \ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa ;
    wire \ALL_SYS_PWRGD.curr_stateZ0Z_1 ;
    wire \ALL_SYS_PWRGD.curr_stateZ0Z_0 ;
    wire \ALL_SYS_PWRGD.un1_curr_state10_0 ;
    wire \ALL_SYS_PWRGD.countZ0Z_9 ;
    wire \ALL_SYS_PWRGD.countZ0Z_1 ;
    wire \ALL_SYS_PWRGD.countZ0Z_10 ;
    wire \ALL_SYS_PWRGD.countZ0Z_0 ;
    wire \ALL_SYS_PWRGD.un4_count_9_cascade_ ;
    wire \ALL_SYS_PWRGD.N_1_i ;
    wire \ALL_SYS_PWRGD.countZ0Z_7 ;
    wire \ALL_SYS_PWRGD.countZ0Z_6 ;
    wire \ALL_SYS_PWRGD.countZ0Z_8 ;
    wire \ALL_SYS_PWRGD.countZ0Z_4 ;
    wire \ALL_SYS_PWRGD.un4_count_8 ;
    wire \ALL_SYS_PWRGD.countZ0Z_3 ;
    wire \ALL_SYS_PWRGD.countZ0Z_11 ;
    wire \ALL_SYS_PWRGD.countZ0Z_5 ;
    wire \ALL_SYS_PWRGD.countZ0Z_2 ;
    wire \ALL_SYS_PWRGD.un4_count_10 ;
    wire vddq_ok;
    wire v5s_ok;
    wire vccst_cpu_ok;
    wire rsmrst_pwrgd_signal;
    wire \ALL_SYS_PWRGD.m4_0_0_a2_1_cascade_ ;
    wire v33s_ok;
    wire \ALL_SYS_PWRGD.N_245 ;
    wire \ALL_SYS_PWRGD.countZ0Z_14 ;
    wire \ALL_SYS_PWRGD.countZ0Z_13 ;
    wire \ALL_SYS_PWRGD.countZ0Z_15 ;
    wire \ALL_SYS_PWRGD.countZ0Z_12 ;
    wire \ALL_SYS_PWRGD.un4_count_11 ;
    wire \ALL_SYS_PWRGD.curr_state_RNIDP9H7Z0Z_1 ;
    wire \ALL_SYS_PWRGD.N_49_4 ;
    wire \POWERLED.N_48 ;
    wire \POWERLED.count_offZ0Z_0 ;
    wire \POWERLED.un1_count_off_1_cry_1_THRU_CO ;
    wire \POWERLED.count_offZ0Z_2 ;
    wire \POWERLED.un1_count_off_1_cry_4_THRU_CO ;
    wire \POWERLED.count_offZ0Z_5 ;
    wire \POWERLED.count_off_0_sqmuxa ;
    wire \POWERLED.N_205 ;
    wire \POWERLED.un1_count_off_1_cry_5_THRU_CO ;
    wire \POWERLED.count_offZ0Z_6 ;
    wire fpga_osc;
    wire N_49_g;
    wire _gnd_net_;

    defparam ipInertedIOPad_VR_READY_VCCINAUX_iopad.PULLUP=1'b0;
    IO_PAD ipInertedIOPad_VR_READY_VCCINAUX_iopad (
            .OE(N__19975),
            .DIN(N__19974),
            .DOUT(N__19973),
            .PACKAGEPIN(VR_READY_VCCINAUX));
    defparam ipInertedIOPad_VR_READY_VCCINAUX_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCINAUX_preio (
            .PADOEN(N__19975),
            .PADOUT(N__19974),
            .PADIN(N__19973),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_ENn_iopad (
            .OE(N__19966),
            .DIN(N__19965),
            .DOUT(N__19964),
            .PACKAGEPIN(V33A_ENn));
    defparam ipInertedIOPad_V33A_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33A_ENn_preio (
            .PADOEN(N__19966),
            .PADOUT(N__19965),
            .PADIN(N__19964),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V1P8A_EN_iopad (
            .OE(N__19957),
            .DIN(N__19956),
            .DOUT(N__19955),
            .PACKAGEPIN(V1P8A_EN));
    defparam ipInertedIOPad_V1P8A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V1P8A_EN_preio (
            .PADOEN(N__19957),
            .PADOUT(N__19956),
            .PADIN(N__19955),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__9311),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDDQ_EN_iopad (
            .OE(N__19948),
            .DIN(N__19947),
            .DOUT(N__19946),
            .PACKAGEPIN(VDDQ_EN));
    defparam ipInertedIOPad_VDDQ_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDDQ_EN_preio (
            .PADOEN(N__19948),
            .PADOUT(N__19947),
            .PADIN(N__19946),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__8793),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad (
            .OE(N__19939),
            .DIN(N__19938),
            .DOUT(N__19937),
            .PACKAGEPIN(VCCST_OVERRIDE_3V3));
    defparam ipInertedIOPad_VCCST_OVERRIDE_3V3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_OVERRIDE_3V3_preio (
            .PADOEN(N__19939),
            .PADOUT(N__19938),
            .PADIN(N__19937),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_OK_iopad (
            .OE(N__19930),
            .DIN(N__19929),
            .DOUT(N__19928),
            .PACKAGEPIN(V5S_OK));
    defparam ipInertedIOPad_V5S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5S_OK_preio (
            .PADOEN(N__19930),
            .PADOUT(N__19929),
            .PADIN(N__19928),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S3n_iopad (
            .OE(N__19921),
            .DIN(N__19920),
            .DOUT(N__19919),
            .PACKAGEPIN(SLP_S3n));
    defparam ipInertedIOPad_SLP_S3n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S3n_preio (
            .PADOEN(N__19921),
            .PADOUT(N__19920),
            .PADIN(N__19919),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s3n),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S0n_iopad (
            .OE(N__19912),
            .DIN(N__19911),
            .DOUT(N__19910),
            .PACKAGEPIN(SLP_S0n));
    defparam ipInertedIOPad_SLP_S0n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S0n_preio (
            .PADOEN(N__19912),
            .PADOUT(N__19911),
            .PADIN(N__19910),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_ENn_iopad (
            .OE(N__19903),
            .DIN(N__19902),
            .DOUT(N__19901),
            .PACKAGEPIN(V5S_ENn));
    defparam ipInertedIOPad_V5S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5S_ENn_preio (
            .PADOEN(N__19903),
            .PADOUT(N__19902),
            .PADIN(N__19901),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__9765),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V1P8A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V1P8A_OK_iopad (
            .OE(N__19894),
            .DIN(N__19893),
            .DOUT(N__19892),
            .PACKAGEPIN(V1P8A_OK));
    defparam ipInertedIOPad_V1P8A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V1P8A_OK_preio (
            .PADOEN(N__19894),
            .PADOUT(N__19893),
            .PADIN(N__19892),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v1p8a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTNn_iopad (
            .OE(N__19885),
            .DIN(N__19884),
            .DOUT(N__19883),
            .PACKAGEPIN(PWRBTNn));
    defparam ipInertedIOPad_PWRBTNn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PWRBTNn_preio (
            .PADOEN(N__19885),
            .PADOUT(N__19884),
            .PADIN(N__19883),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTN_LED_iopad (
            .OE(N__19876),
            .DIN(N__19875),
            .DOUT(N__19874),
            .PACKAGEPIN(PWRBTN_LED));
    defparam ipInertedIOPad_PWRBTN_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PWRBTN_LED_preio (
            .PADOEN(N__19876),
            .PADOUT(N__19875),
            .PADIN(N__19874),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__10107),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_2_iopad (
            .OE(N__19867),
            .DIN(N__19866),
            .DOUT(N__19865),
            .PACKAGEPIN(GPIO_FPGA_SoC_2));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_2_preio (
            .PADOEN(N__19867),
            .PADOUT(N__19866),
            .PADIN(N__19865),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad (
            .OE(N__19858),
            .DIN(N__19857),
            .DOUT(N__19856),
            .PACKAGEPIN(VCCIN_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__19858),
            .PADOUT(N__19857),
            .PADIN(N__19856),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_SLP_SUSn_iopad.PULLUP=1'b0;
    IO_PAD ipInertedIOPad_SLP_SUSn_iopad (
            .OE(N__19849),
            .DIN(N__19848),
            .DOUT(N__19847),
            .PACKAGEPIN(SLP_SUSn));
    defparam ipInertedIOPad_SLP_SUSn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_SUSn_preio (
            .PADOEN(N__19849),
            .PADOUT(N__19848),
            .PADIN(N__19847),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_susn),
            .DIN1());
    IO_PAD ipInertedIOPad_CPU_C10_GATE_N_iopad (
            .OE(N__19840),
            .DIN(N__19839),
            .DOUT(N__19838),
            .PACKAGEPIN(CPU_C10_GATE_N));
    defparam ipInertedIOPad_CPU_C10_GATE_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_CPU_C10_GATE_N_preio (
            .PADOEN(N__19840),
            .PADOUT(N__19839),
            .PADIN(N__19838),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_EN_iopad (
            .OE(N__19831),
            .DIN(N__19830),
            .DOUT(N__19829),
            .PACKAGEPIN(VCCST_EN));
    defparam ipInertedIOPad_VCCST_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_EN_preio (
            .PADOEN(N__19831),
            .PADOUT(N__19830),
            .PADIN(N__19829),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16783),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V33DSW_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V33DSW_OK_iopad (
            .OE(N__19822),
            .DIN(N__19821),
            .DOUT(N__19820),
            .PACKAGEPIN(V33DSW_OK));
    defparam ipInertedIOPad_V33DSW_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33DSW_OK_preio (
            .PADOEN(N__19822),
            .PADOUT(N__19821),
            .PADIN(N__19820),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_TPM_GPIO_iopad (
            .OE(N__19813),
            .DIN(N__19812),
            .DOUT(N__19811),
            .PACKAGEPIN(TPM_GPIO));
    defparam ipInertedIOPad_TPM_GPIO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_TPM_GPIO_preio (
            .PADOEN(N__19813),
            .PADOUT(N__19812),
            .PADIN(N__19811),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSWARN_N_iopad (
            .OE(N__19804),
            .DIN(N__19803),
            .DOUT(N__19802),
            .PACKAGEPIN(SUSWARN_N));
    defparam ipInertedIOPad_SUSWARN_N_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SUSWARN_N_preio (
            .PADOEN(N__19804),
            .PADOUT(N__19803),
            .PADIN(N__19802),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16914),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PLTRSTn_iopad (
            .OE(N__19795),
            .DIN(N__19794),
            .DOUT(N__19793),
            .PACKAGEPIN(PLTRSTn));
    defparam ipInertedIOPad_PLTRSTn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PLTRSTn_preio (
            .PADOEN(N__19795),
            .PADOUT(N__19794),
            .PADIN(N__19793),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_4_iopad (
            .OE(N__19786),
            .DIN(N__19785),
            .DOUT(N__19784),
            .PACKAGEPIN(GPIO_FPGA_SoC_4));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_4_preio (
            .PADOEN(N__19786),
            .PADOUT(N__19785),
            .PADIN(N__19784),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_4),
            .DIN1());
    defparam ipInertedIOPad_VR_READY_VCCIN_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VR_READY_VCCIN_iopad (
            .OE(N__19777),
            .DIN(N__19776),
            .DOUT(N__19775),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam ipInertedIOPad_VR_READY_VCCIN_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCIN_preio (
            .PADOEN(N__19777),
            .PADOUT(N__19776),
            .PADIN(N__19775),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccin),
            .DIN1());
    defparam ipInertedIOPad_V5A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V5A_OK_iopad (
            .OE(N__19768),
            .DIN(N__19767),
            .DOUT(N__19766),
            .PACKAGEPIN(V5A_OK));
    defparam ipInertedIOPad_V5A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5A_OK_preio (
            .PADOEN(N__19768),
            .PADOUT(N__19767),
            .PADIN(N__19766),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_RSMRSTn_iopad (
            .OE(N__19759),
            .DIN(N__19758),
            .DOUT(N__19757),
            .PACKAGEPIN(RSMRSTn));
    defparam ipInertedIOPad_RSMRSTn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RSMRSTn_preio (
            .PADOEN(N__19759),
            .PADOUT(N__19758),
            .PADIN(N__19757),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__14721),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_OSC_iopad (
            .OE(N__19750),
            .DIN(N__19749),
            .DOUT(N__19748),
            .PACKAGEPIN(FPGA_OSC));
    defparam ipInertedIOPad_FPGA_OSC_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_OSC_preio (
            .PADOEN(N__19750),
            .PADOUT(N__19749),
            .PADIN(N__19748),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(fpga_osc),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_PWRGD_iopad (
            .OE(N__19741),
            .DIN(N__19740),
            .DOUT(N__19739),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam ipInertedIOPad_VCCST_PWRGD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_PWRGD_preio (
            .PADOEN(N__19741),
            .PADOUT(N__19740),
            .PADIN(N__19739),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16970),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SYS_PWROK_iopad (
            .OE(N__19732),
            .DIN(N__19731),
            .DOUT(N__19730),
            .PACKAGEPIN(SYS_PWROK));
    defparam ipInertedIOPad_SYS_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SYS_PWROK_preio (
            .PADOEN(N__19732),
            .PADOUT(N__19731),
            .PADIN(N__19730),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__13050),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO2_iopad (
            .OE(N__19723),
            .DIN(N__19722),
            .DOUT(N__19721),
            .PACKAGEPIN(SPI_FP_IO2));
    defparam ipInertedIOPad_SPI_FP_IO2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO2_preio (
            .PADOEN(N__19723),
            .PADOUT(N__19722),
            .PADIN(N__19721),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE1_FPGA_iopad (
            .OE(N__19714),
            .DIN(N__19713),
            .DOUT(N__19712),
            .PACKAGEPIN(SATAXPCIE1_FPGA));
    defparam ipInertedIOPad_SATAXPCIE1_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE1_FPGA_preio (
            .PADOEN(N__19714),
            .PADOUT(N__19713),
            .PADIN(N__19712),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_1_iopad (
            .OE(N__19705),
            .DIN(N__19704),
            .DOUT(N__19703),
            .PACKAGEPIN(GPIO_FPGA_EXP_1));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_1_preio (
            .PADOEN(N__19705),
            .PADOUT(N__19704),
            .PADIN(N__19703),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad (
            .OE(N__19696),
            .DIN(N__19695),
            .DOUT(N__19694),
            .PACKAGEPIN(VCCINAUX_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__19696),
            .PADOUT(N__19695),
            .PADIN(N__19694),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PE_iopad (
            .OE(N__19687),
            .DIN(N__19686),
            .DOUT(N__19685),
            .PACKAGEPIN(VCCINAUX_VR_PE));
    defparam ipInertedIOPad_VCCINAUX_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PE_preio (
            .PADOEN(N__19687),
            .PADOUT(N__19686),
            .PADIN(N__19685),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_HDA_SDO_ATP_iopad (
            .OE(N__19678),
            .DIN(N__19677),
            .DOUT(N__19676),
            .PACKAGEPIN(HDA_SDO_ATP));
    defparam ipInertedIOPad_HDA_SDO_ATP_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_HDA_SDO_ATP_preio (
            .PADOEN(N__19678),
            .PADOUT(N__19677),
            .PADIN(N__19676),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_2_iopad (
            .OE(N__19669),
            .DIN(N__19668),
            .DOUT(N__19667),
            .PACKAGEPIN(GPIO_FPGA_EXP_2));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_2_preio (
            .PADOEN(N__19669),
            .PADOUT(N__19668),
            .PADIN(N__19667),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VPP_EN_iopad (
            .OE(N__19660),
            .DIN(N__19659),
            .DOUT(N__19658),
            .PACKAGEPIN(VPP_EN));
    defparam ipInertedIOPad_VPP_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VPP_EN_preio (
            .PADOEN(N__19660),
            .PADOUT(N__19659),
            .PADIN(N__19658),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17610),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VDDQ_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VDDQ_OK_iopad (
            .OE(N__19651),
            .DIN(N__19650),
            .DOUT(N__19649),
            .PACKAGEPIN(VDDQ_OK));
    defparam ipInertedIOPad_VDDQ_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDDQ_OK_preio (
            .PADOEN(N__19651),
            .PADOUT(N__19650),
            .PADIN(N__19649),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vddq_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSACK_N_iopad (
            .OE(N__19642),
            .DIN(N__19641),
            .DOUT(N__19640),
            .PACKAGEPIN(SUSACK_N));
    defparam ipInertedIOPad_SUSACK_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSACK_N_preio (
            .PADOEN(N__19642),
            .PADOUT(N__19641),
            .PADIN(N__19640),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S4n_iopad (
            .OE(N__19633),
            .DIN(N__19632),
            .DOUT(N__19631),
            .PACKAGEPIN(SLP_S4n));
    defparam ipInertedIOPad_SLP_S4n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S4n_preio (
            .PADOEN(N__19633),
            .PADOUT(N__19632),
            .PADIN(N__19631),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s4n),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_CPU_OK_iopad (
            .OE(N__19624),
            .DIN(N__19623),
            .DOUT(N__19622),
            .PACKAGEPIN(VCCST_CPU_OK));
    defparam ipInertedIOPad_VCCST_CPU_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_CPU_OK_preio (
            .PADOEN(N__19624),
            .PADOUT(N__19623),
            .PADIN(N__19622),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vccst_cpu_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_EN_iopad (
            .OE(N__19615),
            .DIN(N__19614),
            .DOUT(N__19613),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam ipInertedIOPad_VCCINAUX_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_EN_preio (
            .PADOEN(N__19615),
            .PADOUT(N__19614),
            .PADIN(N__19613),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__9237),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_OK_iopad (
            .OE(N__19606),
            .DIN(N__19605),
            .DOUT(N__19604),
            .PACKAGEPIN(V33S_OK));
    defparam ipInertedIOPad_V33S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33S_OK_preio (
            .PADOEN(N__19606),
            .PADOUT(N__19605),
            .PADIN(N__19604),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_ENn_iopad (
            .OE(N__19597),
            .DIN(N__19596),
            .DOUT(N__19595),
            .PACKAGEPIN(V33S_ENn));
    defparam ipInertedIOPad_V33S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33S_ENn_preio (
            .PADOEN(N__19597),
            .PADOUT(N__19596),
            .PADIN(N__19595),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__9761),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_1_iopad (
            .OE(N__19588),
            .DIN(N__19587),
            .DOUT(N__19586),
            .PACKAGEPIN(GPIO_FPGA_SoC_1));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_1_preio (
            .PADOEN(N__19588),
            .PADOUT(N__19587),
            .PADIN(N__19586),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_DSW_PWROK_iopad.PULLUP=1'b0;
    IO_PAD ipInertedIOPad_DSW_PWROK_iopad (
            .OE(N__19579),
            .DIN(N__19578),
            .DOUT(N__19577),
            .PACKAGEPIN(DSW_PWROK));
    defparam ipInertedIOPad_DSW_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DSW_PWROK_preio (
            .PADOEN(N__19579),
            .PADOUT(N__19578),
            .PADIN(N__19577),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17300),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5A_EN_iopad (
            .OE(N__19570),
            .DIN(N__19569),
            .DOUT(N__19568),
            .PACKAGEPIN(V5A_EN));
    defparam ipInertedIOPad_V5A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5A_EN_preio (
            .PADOEN(N__19570),
            .PADOUT(N__19569),
            .PADIN(N__19568),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__9310),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_3_iopad (
            .OE(N__19561),
            .DIN(N__19560),
            .DOUT(N__19559),
            .PACKAGEPIN(GPIO_FPGA_SoC_3));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_3_preio (
            .PADOEN(N__19561),
            .PADOUT(N__19560),
            .PADIN(N__19559),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad (
            .OE(N__19552),
            .DIN(N__19551),
            .DOUT(N__19550),
            .PACKAGEPIN(VR_PROCHOT_FPGA_OUT_N));
    defparam ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio (
            .PADOEN(N__19552),
            .PADOUT(N__19551),
            .PADIN(N__19550),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VPP_OK_iopad.PULLUP=1'b0;
    IO_PAD ipInertedIOPad_VPP_OK_iopad (
            .OE(N__19543),
            .DIN(N__19542),
            .DOUT(N__19541),
            .PACKAGEPIN(VPP_OK));
    defparam ipInertedIOPad_VPP_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VPP_OK_preio (
            .PADOEN(N__19543),
            .PADOUT(N__19542),
            .PADIN(N__19541),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vpp_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PE_iopad (
            .OE(N__19534),
            .DIN(N__19533),
            .DOUT(N__19532),
            .PACKAGEPIN(VCCIN_VR_PE));
    defparam ipInertedIOPad_VCCIN_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PE_preio (
            .PADOEN(N__19534),
            .PADOUT(N__19533),
            .PADIN(N__19532),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_EN_iopad (
            .OE(N__19525),
            .DIN(N__19524),
            .DOUT(N__19523),
            .PACKAGEPIN(VCCIN_EN));
    defparam ipInertedIOPad_VCCIN_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_EN_preio (
            .PADOEN(N__19525),
            .PADOUT(N__19524),
            .PADIN(N__19523),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16977),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SOC_SPKR_iopad (
            .OE(N__19516),
            .DIN(N__19515),
            .DOUT(N__19514),
            .PACKAGEPIN(SOC_SPKR));
    defparam ipInertedIOPad_SOC_SPKR_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SOC_SPKR_preio (
            .PADOEN(N__19516),
            .PADOUT(N__19515),
            .PADIN(N__19514),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S5n_iopad (
            .OE(N__19507),
            .DIN(N__19506),
            .DOUT(N__19505),
            .PACKAGEPIN(SLP_S5n));
    defparam ipInertedIOPad_SLP_S5n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S5n_preio (
            .PADOEN(N__19507),
            .PADOUT(N__19506),
            .PADIN(N__19505),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V12_MAIN_MON_iopad (
            .OE(N__19498),
            .DIN(N__19497),
            .DOUT(N__19496),
            .PACKAGEPIN(V12_MAIN_MON));
    defparam ipInertedIOPad_V12_MAIN_MON_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V12_MAIN_MON_preio (
            .PADOEN(N__19498),
            .PADOUT(N__19497),
            .PADIN(N__19496),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO3_iopad (
            .OE(N__19489),
            .DIN(N__19488),
            .DOUT(N__19487),
            .PACKAGEPIN(SPI_FP_IO3));
    defparam ipInertedIOPad_SPI_FP_IO3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO3_preio (
            .PADOEN(N__19489),
            .PADOUT(N__19488),
            .PADIN(N__19487),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE0_FPGA_iopad (
            .OE(N__19480),
            .DIN(N__19479),
            .DOUT(N__19478),
            .PACKAGEPIN(SATAXPCIE0_FPGA));
    defparam ipInertedIOPad_SATAXPCIE0_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE0_FPGA_preio (
            .PADOEN(N__19480),
            .PADOUT(N__19479),
            .PADIN(N__19478),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_OK_iopad (
            .OE(N__19471),
            .DIN(N__19470),
            .DOUT(N__19469),
            .PACKAGEPIN(V33A_OK));
    defparam ipInertedIOPad_V33A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33A_OK_preio (
            .PADOEN(N__19471),
            .PADOUT(N__19470),
            .PADIN(N__19469),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PCH_PWROK_iopad (
            .OE(N__19462),
            .DIN(N__19461),
            .DOUT(N__19460),
            .PACKAGEPIN(PCH_PWROK));
    defparam ipInertedIOPad_PCH_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PCH_PWROK_preio (
            .PADOEN(N__19462),
            .PADOUT(N__19461),
            .PADIN(N__19460),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__13037),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_SLP_WLAN_N_iopad (
            .OE(N__19453),
            .DIN(N__19452),
            .DOUT(N__19451),
            .PACKAGEPIN(FPGA_SLP_WLAN_N));
    defparam ipInertedIOPad_FPGA_SLP_WLAN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_SLP_WLAN_N_preio (
            .PADOEN(N__19453),
            .PADOUT(N__19452),
            .PADIN(N__19451),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    InMux I__4416 (
            .O(N__19434),
            .I(N__19431));
    LocalMux I__4415 (
            .O(N__19431),
            .I(\POWERLED.un1_count_off_1_cry_1_THRU_CO ));
    CascadeMux I__4414 (
            .O(N__19428),
            .I(N__19424));
    InMux I__4413 (
            .O(N__19427),
            .I(N__19420));
    InMux I__4412 (
            .O(N__19424),
            .I(N__19417));
    InMux I__4411 (
            .O(N__19423),
            .I(N__19414));
    LocalMux I__4410 (
            .O(N__19420),
            .I(N__19411));
    LocalMux I__4409 (
            .O(N__19417),
            .I(\POWERLED.count_offZ0Z_2 ));
    LocalMux I__4408 (
            .O(N__19414),
            .I(\POWERLED.count_offZ0Z_2 ));
    Odrv4 I__4407 (
            .O(N__19411),
            .I(\POWERLED.count_offZ0Z_2 ));
    InMux I__4406 (
            .O(N__19404),
            .I(N__19401));
    LocalMux I__4405 (
            .O(N__19401),
            .I(\POWERLED.un1_count_off_1_cry_4_THRU_CO ));
    CascadeMux I__4404 (
            .O(N__19398),
            .I(N__19394));
    InMux I__4403 (
            .O(N__19397),
            .I(N__19390));
    InMux I__4402 (
            .O(N__19394),
            .I(N__19387));
    InMux I__4401 (
            .O(N__19393),
            .I(N__19384));
    LocalMux I__4400 (
            .O(N__19390),
            .I(N__19381));
    LocalMux I__4399 (
            .O(N__19387),
            .I(\POWERLED.count_offZ0Z_5 ));
    LocalMux I__4398 (
            .O(N__19384),
            .I(\POWERLED.count_offZ0Z_5 ));
    Odrv4 I__4397 (
            .O(N__19381),
            .I(\POWERLED.count_offZ0Z_5 ));
    InMux I__4396 (
            .O(N__19374),
            .I(N__19371));
    LocalMux I__4395 (
            .O(N__19371),
            .I(N__19353));
    InMux I__4394 (
            .O(N__19370),
            .I(N__19344));
    InMux I__4393 (
            .O(N__19369),
            .I(N__19344));
    InMux I__4392 (
            .O(N__19368),
            .I(N__19344));
    InMux I__4391 (
            .O(N__19367),
            .I(N__19344));
    InMux I__4390 (
            .O(N__19366),
            .I(N__19337));
    InMux I__4389 (
            .O(N__19365),
            .I(N__19337));
    InMux I__4388 (
            .O(N__19364),
            .I(N__19337));
    InMux I__4387 (
            .O(N__19363),
            .I(N__19330));
    InMux I__4386 (
            .O(N__19362),
            .I(N__19330));
    InMux I__4385 (
            .O(N__19361),
            .I(N__19330));
    InMux I__4384 (
            .O(N__19360),
            .I(N__19319));
    InMux I__4383 (
            .O(N__19359),
            .I(N__19319));
    InMux I__4382 (
            .O(N__19358),
            .I(N__19319));
    InMux I__4381 (
            .O(N__19357),
            .I(N__19319));
    InMux I__4380 (
            .O(N__19356),
            .I(N__19319));
    Span4Mux_v I__4379 (
            .O(N__19353),
            .I(N__19316));
    LocalMux I__4378 (
            .O(N__19344),
            .I(N__19309));
    LocalMux I__4377 (
            .O(N__19337),
            .I(N__19309));
    LocalMux I__4376 (
            .O(N__19330),
            .I(N__19309));
    LocalMux I__4375 (
            .O(N__19319),
            .I(N__19302));
    Span4Mux_s0_h I__4374 (
            .O(N__19316),
            .I(N__19302));
    Span4Mux_v I__4373 (
            .O(N__19309),
            .I(N__19302));
    Odrv4 I__4372 (
            .O(N__19302),
            .I(\POWERLED.count_off_0_sqmuxa ));
    InMux I__4371 (
            .O(N__19299),
            .I(N__19287));
    InMux I__4370 (
            .O(N__19298),
            .I(N__19287));
    InMux I__4369 (
            .O(N__19297),
            .I(N__19287));
    InMux I__4368 (
            .O(N__19296),
            .I(N__19287));
    LocalMux I__4367 (
            .O(N__19287),
            .I(N__19284));
    Span4Mux_s2_h I__4366 (
            .O(N__19284),
            .I(N__19281));
    Odrv4 I__4365 (
            .O(N__19281),
            .I(\POWERLED.N_205 ));
    InMux I__4364 (
            .O(N__19278),
            .I(N__19275));
    LocalMux I__4363 (
            .O(N__19275),
            .I(\POWERLED.un1_count_off_1_cry_5_THRU_CO ));
    CascadeMux I__4362 (
            .O(N__19272),
            .I(N__19268));
    InMux I__4361 (
            .O(N__19271),
            .I(N__19264));
    InMux I__4360 (
            .O(N__19268),
            .I(N__19261));
    InMux I__4359 (
            .O(N__19267),
            .I(N__19258));
    LocalMux I__4358 (
            .O(N__19264),
            .I(N__19255));
    LocalMux I__4357 (
            .O(N__19261),
            .I(\POWERLED.count_offZ0Z_6 ));
    LocalMux I__4356 (
            .O(N__19258),
            .I(\POWERLED.count_offZ0Z_6 ));
    Odrv4 I__4355 (
            .O(N__19255),
            .I(\POWERLED.count_offZ0Z_6 ));
    ClkMux I__4354 (
            .O(N__19248),
            .I(N__19245));
    LocalMux I__4353 (
            .O(N__19245),
            .I(N__19239));
    ClkMux I__4352 (
            .O(N__19244),
            .I(N__19236));
    ClkMux I__4351 (
            .O(N__19243),
            .I(N__19233));
    ClkMux I__4350 (
            .O(N__19242),
            .I(N__19226));
    Span4Mux_v I__4349 (
            .O(N__19239),
            .I(N__19215));
    LocalMux I__4348 (
            .O(N__19236),
            .I(N__19215));
    LocalMux I__4347 (
            .O(N__19233),
            .I(N__19215));
    ClkMux I__4346 (
            .O(N__19232),
            .I(N__19207));
    ClkMux I__4345 (
            .O(N__19231),
            .I(N__19204));
    ClkMux I__4344 (
            .O(N__19230),
            .I(N__19201));
    ClkMux I__4343 (
            .O(N__19229),
            .I(N__19198));
    LocalMux I__4342 (
            .O(N__19226),
            .I(N__19195));
    ClkMux I__4341 (
            .O(N__19225),
            .I(N__19192));
    ClkMux I__4340 (
            .O(N__19224),
            .I(N__19189));
    ClkMux I__4339 (
            .O(N__19223),
            .I(N__19186));
    ClkMux I__4338 (
            .O(N__19222),
            .I(N__19182));
    Span4Mux_v I__4337 (
            .O(N__19215),
            .I(N__19178));
    ClkMux I__4336 (
            .O(N__19214),
            .I(N__19175));
    ClkMux I__4335 (
            .O(N__19213),
            .I(N__19171));
    ClkMux I__4334 (
            .O(N__19212),
            .I(N__19167));
    ClkMux I__4333 (
            .O(N__19211),
            .I(N__19163));
    ClkMux I__4332 (
            .O(N__19210),
            .I(N__19160));
    LocalMux I__4331 (
            .O(N__19207),
            .I(N__19156));
    LocalMux I__4330 (
            .O(N__19204),
            .I(N__19151));
    LocalMux I__4329 (
            .O(N__19201),
            .I(N__19146));
    LocalMux I__4328 (
            .O(N__19198),
            .I(N__19146));
    Span4Mux_h I__4327 (
            .O(N__19195),
            .I(N__19139));
    LocalMux I__4326 (
            .O(N__19192),
            .I(N__19139));
    LocalMux I__4325 (
            .O(N__19189),
            .I(N__19139));
    LocalMux I__4324 (
            .O(N__19186),
            .I(N__19134));
    ClkMux I__4323 (
            .O(N__19185),
            .I(N__19131));
    LocalMux I__4322 (
            .O(N__19182),
            .I(N__19127));
    ClkMux I__4321 (
            .O(N__19181),
            .I(N__19124));
    Span4Mux_h I__4320 (
            .O(N__19178),
            .I(N__19119));
    LocalMux I__4319 (
            .O(N__19175),
            .I(N__19119));
    ClkMux I__4318 (
            .O(N__19174),
            .I(N__19116));
    LocalMux I__4317 (
            .O(N__19171),
            .I(N__19111));
    ClkMux I__4316 (
            .O(N__19170),
            .I(N__19108));
    LocalMux I__4315 (
            .O(N__19167),
            .I(N__19105));
    ClkMux I__4314 (
            .O(N__19166),
            .I(N__19102));
    LocalMux I__4313 (
            .O(N__19163),
            .I(N__19097));
    LocalMux I__4312 (
            .O(N__19160),
            .I(N__19097));
    ClkMux I__4311 (
            .O(N__19159),
            .I(N__19094));
    Span4Mux_s1_h I__4310 (
            .O(N__19156),
            .I(N__19090));
    ClkMux I__4309 (
            .O(N__19155),
            .I(N__19087));
    ClkMux I__4308 (
            .O(N__19154),
            .I(N__19082));
    Span4Mux_h I__4307 (
            .O(N__19151),
            .I(N__19074));
    Span4Mux_v I__4306 (
            .O(N__19146),
            .I(N__19074));
    Span4Mux_v I__4305 (
            .O(N__19139),
            .I(N__19074));
    ClkMux I__4304 (
            .O(N__19138),
            .I(N__19071));
    ClkMux I__4303 (
            .O(N__19137),
            .I(N__19068));
    Span4Mux_v I__4302 (
            .O(N__19134),
            .I(N__19061));
    LocalMux I__4301 (
            .O(N__19131),
            .I(N__19061));
    ClkMux I__4300 (
            .O(N__19130),
            .I(N__19058));
    Span4Mux_v I__4299 (
            .O(N__19127),
            .I(N__19049));
    LocalMux I__4298 (
            .O(N__19124),
            .I(N__19049));
    Span4Mux_h I__4297 (
            .O(N__19119),
            .I(N__19049));
    LocalMux I__4296 (
            .O(N__19116),
            .I(N__19049));
    ClkMux I__4295 (
            .O(N__19115),
            .I(N__19046));
    ClkMux I__4294 (
            .O(N__19114),
            .I(N__19043));
    Span4Mux_v I__4293 (
            .O(N__19111),
            .I(N__19037));
    LocalMux I__4292 (
            .O(N__19108),
            .I(N__19037));
    Span4Mux_v I__4291 (
            .O(N__19105),
            .I(N__19032));
    LocalMux I__4290 (
            .O(N__19102),
            .I(N__19032));
    Span4Mux_v I__4289 (
            .O(N__19097),
            .I(N__19027));
    LocalMux I__4288 (
            .O(N__19094),
            .I(N__19027));
    ClkMux I__4287 (
            .O(N__19093),
            .I(N__19024));
    Span4Mux_h I__4286 (
            .O(N__19090),
            .I(N__19017));
    LocalMux I__4285 (
            .O(N__19087),
            .I(N__19017));
    ClkMux I__4284 (
            .O(N__19086),
            .I(N__19014));
    ClkMux I__4283 (
            .O(N__19085),
            .I(N__19009));
    LocalMux I__4282 (
            .O(N__19082),
            .I(N__19005));
    ClkMux I__4281 (
            .O(N__19081),
            .I(N__19002));
    Span4Mux_v I__4280 (
            .O(N__19074),
            .I(N__18996));
    LocalMux I__4279 (
            .O(N__19071),
            .I(N__18996));
    LocalMux I__4278 (
            .O(N__19068),
            .I(N__18993));
    ClkMux I__4277 (
            .O(N__19067),
            .I(N__18990));
    ClkMux I__4276 (
            .O(N__19066),
            .I(N__18987));
    Span4Mux_v I__4275 (
            .O(N__19061),
            .I(N__18982));
    LocalMux I__4274 (
            .O(N__19058),
            .I(N__18982));
    Span4Mux_v I__4273 (
            .O(N__19049),
            .I(N__18975));
    LocalMux I__4272 (
            .O(N__19046),
            .I(N__18975));
    LocalMux I__4271 (
            .O(N__19043),
            .I(N__18975));
    ClkMux I__4270 (
            .O(N__19042),
            .I(N__18972));
    Span4Mux_v I__4269 (
            .O(N__19037),
            .I(N__18969));
    Span4Mux_s1_h I__4268 (
            .O(N__19032),
            .I(N__18962));
    Span4Mux_v I__4267 (
            .O(N__19027),
            .I(N__18962));
    LocalMux I__4266 (
            .O(N__19024),
            .I(N__18962));
    ClkMux I__4265 (
            .O(N__19023),
            .I(N__18959));
    ClkMux I__4264 (
            .O(N__19022),
            .I(N__18955));
    Span4Mux_v I__4263 (
            .O(N__19017),
            .I(N__18950));
    LocalMux I__4262 (
            .O(N__19014),
            .I(N__18950));
    ClkMux I__4261 (
            .O(N__19013),
            .I(N__18947));
    ClkMux I__4260 (
            .O(N__19012),
            .I(N__18944));
    LocalMux I__4259 (
            .O(N__19009),
            .I(N__18941));
    ClkMux I__4258 (
            .O(N__19008),
            .I(N__18938));
    Span4Mux_v I__4257 (
            .O(N__19005),
            .I(N__18932));
    LocalMux I__4256 (
            .O(N__19002),
            .I(N__18932));
    ClkMux I__4255 (
            .O(N__19001),
            .I(N__18929));
    Span4Mux_v I__4254 (
            .O(N__18996),
            .I(N__18920));
    Span4Mux_v I__4253 (
            .O(N__18993),
            .I(N__18920));
    LocalMux I__4252 (
            .O(N__18990),
            .I(N__18920));
    LocalMux I__4251 (
            .O(N__18987),
            .I(N__18920));
    Span4Mux_v I__4250 (
            .O(N__18982),
            .I(N__18913));
    Span4Mux_v I__4249 (
            .O(N__18975),
            .I(N__18913));
    LocalMux I__4248 (
            .O(N__18972),
            .I(N__18913));
    Span4Mux_h I__4247 (
            .O(N__18969),
            .I(N__18906));
    Span4Mux_h I__4246 (
            .O(N__18962),
            .I(N__18906));
    LocalMux I__4245 (
            .O(N__18959),
            .I(N__18906));
    ClkMux I__4244 (
            .O(N__18958),
            .I(N__18903));
    LocalMux I__4243 (
            .O(N__18955),
            .I(N__18900));
    Span4Mux_v I__4242 (
            .O(N__18950),
            .I(N__18895));
    LocalMux I__4241 (
            .O(N__18947),
            .I(N__18895));
    LocalMux I__4240 (
            .O(N__18944),
            .I(N__18891));
    Sp12to4 I__4239 (
            .O(N__18941),
            .I(N__18886));
    LocalMux I__4238 (
            .O(N__18938),
            .I(N__18886));
    ClkMux I__4237 (
            .O(N__18937),
            .I(N__18883));
    Span4Mux_h I__4236 (
            .O(N__18932),
            .I(N__18878));
    LocalMux I__4235 (
            .O(N__18929),
            .I(N__18878));
    IoSpan4Mux I__4234 (
            .O(N__18920),
            .I(N__18873));
    IoSpan4Mux I__4233 (
            .O(N__18913),
            .I(N__18873));
    Span4Mux_v I__4232 (
            .O(N__18906),
            .I(N__18868));
    LocalMux I__4231 (
            .O(N__18903),
            .I(N__18868));
    Span4Mux_v I__4230 (
            .O(N__18900),
            .I(N__18863));
    Span4Mux_h I__4229 (
            .O(N__18895),
            .I(N__18863));
    ClkMux I__4228 (
            .O(N__18894),
            .I(N__18860));
    Span12Mux_s5_h I__4227 (
            .O(N__18891),
            .I(N__18851));
    Span12Mux_s7_v I__4226 (
            .O(N__18886),
            .I(N__18851));
    LocalMux I__4225 (
            .O(N__18883),
            .I(N__18851));
    Sp12to4 I__4224 (
            .O(N__18878),
            .I(N__18851));
    Odrv4 I__4223 (
            .O(N__18873),
            .I(fpga_osc));
    Odrv4 I__4222 (
            .O(N__18868),
            .I(fpga_osc));
    Odrv4 I__4221 (
            .O(N__18863),
            .I(fpga_osc));
    LocalMux I__4220 (
            .O(N__18860),
            .I(fpga_osc));
    Odrv12 I__4219 (
            .O(N__18851),
            .I(fpga_osc));
    InMux I__4218 (
            .O(N__18840),
            .I(N__18728));
    InMux I__4217 (
            .O(N__18839),
            .I(N__18728));
    InMux I__4216 (
            .O(N__18838),
            .I(N__18728));
    InMux I__4215 (
            .O(N__18837),
            .I(N__18728));
    InMux I__4214 (
            .O(N__18836),
            .I(N__18719));
    InMux I__4213 (
            .O(N__18835),
            .I(N__18719));
    InMux I__4212 (
            .O(N__18834),
            .I(N__18719));
    InMux I__4211 (
            .O(N__18833),
            .I(N__18719));
    InMux I__4210 (
            .O(N__18832),
            .I(N__18710));
    InMux I__4209 (
            .O(N__18831),
            .I(N__18710));
    InMux I__4208 (
            .O(N__18830),
            .I(N__18710));
    InMux I__4207 (
            .O(N__18829),
            .I(N__18710));
    InMux I__4206 (
            .O(N__18828),
            .I(N__18701));
    InMux I__4205 (
            .O(N__18827),
            .I(N__18701));
    InMux I__4204 (
            .O(N__18826),
            .I(N__18701));
    InMux I__4203 (
            .O(N__18825),
            .I(N__18701));
    InMux I__4202 (
            .O(N__18824),
            .I(N__18692));
    InMux I__4201 (
            .O(N__18823),
            .I(N__18692));
    InMux I__4200 (
            .O(N__18822),
            .I(N__18692));
    InMux I__4199 (
            .O(N__18821),
            .I(N__18692));
    InMux I__4198 (
            .O(N__18820),
            .I(N__18683));
    InMux I__4197 (
            .O(N__18819),
            .I(N__18683));
    InMux I__4196 (
            .O(N__18818),
            .I(N__18683));
    InMux I__4195 (
            .O(N__18817),
            .I(N__18683));
    InMux I__4194 (
            .O(N__18816),
            .I(N__18674));
    InMux I__4193 (
            .O(N__18815),
            .I(N__18674));
    InMux I__4192 (
            .O(N__18814),
            .I(N__18674));
    InMux I__4191 (
            .O(N__18813),
            .I(N__18674));
    InMux I__4190 (
            .O(N__18812),
            .I(N__18667));
    InMux I__4189 (
            .O(N__18811),
            .I(N__18667));
    InMux I__4188 (
            .O(N__18810),
            .I(N__18667));
    InMux I__4187 (
            .O(N__18809),
            .I(N__18658));
    InMux I__4186 (
            .O(N__18808),
            .I(N__18658));
    InMux I__4185 (
            .O(N__18807),
            .I(N__18658));
    InMux I__4184 (
            .O(N__18806),
            .I(N__18658));
    InMux I__4183 (
            .O(N__18805),
            .I(N__18651));
    InMux I__4182 (
            .O(N__18804),
            .I(N__18651));
    InMux I__4181 (
            .O(N__18803),
            .I(N__18651));
    InMux I__4180 (
            .O(N__18802),
            .I(N__18642));
    InMux I__4179 (
            .O(N__18801),
            .I(N__18642));
    InMux I__4178 (
            .O(N__18800),
            .I(N__18642));
    InMux I__4177 (
            .O(N__18799),
            .I(N__18642));
    InMux I__4176 (
            .O(N__18798),
            .I(N__18635));
    InMux I__4175 (
            .O(N__18797),
            .I(N__18635));
    InMux I__4174 (
            .O(N__18796),
            .I(N__18635));
    InMux I__4173 (
            .O(N__18795),
            .I(N__18626));
    InMux I__4172 (
            .O(N__18794),
            .I(N__18626));
    InMux I__4171 (
            .O(N__18793),
            .I(N__18626));
    InMux I__4170 (
            .O(N__18792),
            .I(N__18626));
    InMux I__4169 (
            .O(N__18791),
            .I(N__18619));
    InMux I__4168 (
            .O(N__18790),
            .I(N__18619));
    InMux I__4167 (
            .O(N__18789),
            .I(N__18619));
    InMux I__4166 (
            .O(N__18788),
            .I(N__18610));
    InMux I__4165 (
            .O(N__18787),
            .I(N__18610));
    InMux I__4164 (
            .O(N__18786),
            .I(N__18610));
    InMux I__4163 (
            .O(N__18785),
            .I(N__18610));
    InMux I__4162 (
            .O(N__18784),
            .I(N__18601));
    InMux I__4161 (
            .O(N__18783),
            .I(N__18601));
    InMux I__4160 (
            .O(N__18782),
            .I(N__18601));
    InMux I__4159 (
            .O(N__18781),
            .I(N__18601));
    InMux I__4158 (
            .O(N__18780),
            .I(N__18598));
    InMux I__4157 (
            .O(N__18779),
            .I(N__18595));
    InMux I__4156 (
            .O(N__18778),
            .I(N__18592));
    InMux I__4155 (
            .O(N__18777),
            .I(N__18585));
    InMux I__4154 (
            .O(N__18776),
            .I(N__18585));
    InMux I__4153 (
            .O(N__18775),
            .I(N__18585));
    InMux I__4152 (
            .O(N__18774),
            .I(N__18578));
    InMux I__4151 (
            .O(N__18773),
            .I(N__18578));
    InMux I__4150 (
            .O(N__18772),
            .I(N__18578));
    InMux I__4149 (
            .O(N__18771),
            .I(N__18569));
    InMux I__4148 (
            .O(N__18770),
            .I(N__18569));
    InMux I__4147 (
            .O(N__18769),
            .I(N__18569));
    InMux I__4146 (
            .O(N__18768),
            .I(N__18569));
    InMux I__4145 (
            .O(N__18767),
            .I(N__18562));
    InMux I__4144 (
            .O(N__18766),
            .I(N__18562));
    InMux I__4143 (
            .O(N__18765),
            .I(N__18562));
    InMux I__4142 (
            .O(N__18764),
            .I(N__18559));
    InMux I__4141 (
            .O(N__18763),
            .I(N__18550));
    InMux I__4140 (
            .O(N__18762),
            .I(N__18550));
    InMux I__4139 (
            .O(N__18761),
            .I(N__18550));
    InMux I__4138 (
            .O(N__18760),
            .I(N__18550));
    InMux I__4137 (
            .O(N__18759),
            .I(N__18543));
    InMux I__4136 (
            .O(N__18758),
            .I(N__18543));
    InMux I__4135 (
            .O(N__18757),
            .I(N__18543));
    InMux I__4134 (
            .O(N__18756),
            .I(N__18538));
    InMux I__4133 (
            .O(N__18755),
            .I(N__18538));
    InMux I__4132 (
            .O(N__18754),
            .I(N__18529));
    InMux I__4131 (
            .O(N__18753),
            .I(N__18529));
    InMux I__4130 (
            .O(N__18752),
            .I(N__18529));
    InMux I__4129 (
            .O(N__18751),
            .I(N__18529));
    InMux I__4128 (
            .O(N__18750),
            .I(N__18520));
    InMux I__4127 (
            .O(N__18749),
            .I(N__18520));
    InMux I__4126 (
            .O(N__18748),
            .I(N__18520));
    InMux I__4125 (
            .O(N__18747),
            .I(N__18520));
    InMux I__4124 (
            .O(N__18746),
            .I(N__18517));
    InMux I__4123 (
            .O(N__18745),
            .I(N__18510));
    InMux I__4122 (
            .O(N__18744),
            .I(N__18510));
    InMux I__4121 (
            .O(N__18743),
            .I(N__18510));
    InMux I__4120 (
            .O(N__18742),
            .I(N__18507));
    InMux I__4119 (
            .O(N__18741),
            .I(N__18504));
    InMux I__4118 (
            .O(N__18740),
            .I(N__18501));
    InMux I__4117 (
            .O(N__18739),
            .I(N__18498));
    InMux I__4116 (
            .O(N__18738),
            .I(N__18495));
    InMux I__4115 (
            .O(N__18737),
            .I(N__18492));
    LocalMux I__4114 (
            .O(N__18728),
            .I(N__18482));
    LocalMux I__4113 (
            .O(N__18719),
            .I(N__18478));
    LocalMux I__4112 (
            .O(N__18710),
            .I(N__18469));
    LocalMux I__4111 (
            .O(N__18701),
            .I(N__18465));
    LocalMux I__4110 (
            .O(N__18692),
            .I(N__18462));
    LocalMux I__4109 (
            .O(N__18683),
            .I(N__18459));
    LocalMux I__4108 (
            .O(N__18674),
            .I(N__18456));
    LocalMux I__4107 (
            .O(N__18667),
            .I(N__18453));
    LocalMux I__4106 (
            .O(N__18658),
            .I(N__18450));
    LocalMux I__4105 (
            .O(N__18651),
            .I(N__18447));
    LocalMux I__4104 (
            .O(N__18642),
            .I(N__18444));
    LocalMux I__4103 (
            .O(N__18635),
            .I(N__18440));
    LocalMux I__4102 (
            .O(N__18626),
            .I(N__18437));
    LocalMux I__4101 (
            .O(N__18619),
            .I(N__18434));
    LocalMux I__4100 (
            .O(N__18610),
            .I(N__18430));
    LocalMux I__4099 (
            .O(N__18601),
            .I(N__18427));
    LocalMux I__4098 (
            .O(N__18598),
            .I(N__18424));
    LocalMux I__4097 (
            .O(N__18595),
            .I(N__18421));
    LocalMux I__4096 (
            .O(N__18592),
            .I(N__18418));
    LocalMux I__4095 (
            .O(N__18585),
            .I(N__18415));
    LocalMux I__4094 (
            .O(N__18578),
            .I(N__18412));
    LocalMux I__4093 (
            .O(N__18569),
            .I(N__18409));
    LocalMux I__4092 (
            .O(N__18562),
            .I(N__18406));
    LocalMux I__4091 (
            .O(N__18559),
            .I(N__18403));
    LocalMux I__4090 (
            .O(N__18550),
            .I(N__18400));
    LocalMux I__4089 (
            .O(N__18543),
            .I(N__18397));
    LocalMux I__4088 (
            .O(N__18538),
            .I(N__18394));
    LocalMux I__4087 (
            .O(N__18529),
            .I(N__18391));
    LocalMux I__4086 (
            .O(N__18520),
            .I(N__18388));
    LocalMux I__4085 (
            .O(N__18517),
            .I(N__18385));
    LocalMux I__4084 (
            .O(N__18510),
            .I(N__18382));
    LocalMux I__4083 (
            .O(N__18507),
            .I(N__18379));
    LocalMux I__4082 (
            .O(N__18504),
            .I(N__18376));
    LocalMux I__4081 (
            .O(N__18501),
            .I(N__18373));
    LocalMux I__4080 (
            .O(N__18498),
            .I(N__18370));
    LocalMux I__4079 (
            .O(N__18495),
            .I(N__18367));
    LocalMux I__4078 (
            .O(N__18492),
            .I(N__18364));
    CEMux I__4077 (
            .O(N__18491),
            .I(N__18255));
    CEMux I__4076 (
            .O(N__18490),
            .I(N__18255));
    CEMux I__4075 (
            .O(N__18489),
            .I(N__18255));
    CEMux I__4074 (
            .O(N__18488),
            .I(N__18255));
    CEMux I__4073 (
            .O(N__18487),
            .I(N__18255));
    CEMux I__4072 (
            .O(N__18486),
            .I(N__18255));
    CEMux I__4071 (
            .O(N__18485),
            .I(N__18255));
    Glb2LocalMux I__4070 (
            .O(N__18482),
            .I(N__18255));
    CEMux I__4069 (
            .O(N__18481),
            .I(N__18255));
    Glb2LocalMux I__4068 (
            .O(N__18478),
            .I(N__18255));
    CEMux I__4067 (
            .O(N__18477),
            .I(N__18255));
    CEMux I__4066 (
            .O(N__18476),
            .I(N__18255));
    CEMux I__4065 (
            .O(N__18475),
            .I(N__18255));
    CEMux I__4064 (
            .O(N__18474),
            .I(N__18255));
    CEMux I__4063 (
            .O(N__18473),
            .I(N__18255));
    CEMux I__4062 (
            .O(N__18472),
            .I(N__18255));
    Glb2LocalMux I__4061 (
            .O(N__18469),
            .I(N__18255));
    CEMux I__4060 (
            .O(N__18468),
            .I(N__18255));
    Glb2LocalMux I__4059 (
            .O(N__18465),
            .I(N__18255));
    Glb2LocalMux I__4058 (
            .O(N__18462),
            .I(N__18255));
    Glb2LocalMux I__4057 (
            .O(N__18459),
            .I(N__18255));
    Glb2LocalMux I__4056 (
            .O(N__18456),
            .I(N__18255));
    Glb2LocalMux I__4055 (
            .O(N__18453),
            .I(N__18255));
    Glb2LocalMux I__4054 (
            .O(N__18450),
            .I(N__18255));
    Glb2LocalMux I__4053 (
            .O(N__18447),
            .I(N__18255));
    Glb2LocalMux I__4052 (
            .O(N__18444),
            .I(N__18255));
    CEMux I__4051 (
            .O(N__18443),
            .I(N__18255));
    Glb2LocalMux I__4050 (
            .O(N__18440),
            .I(N__18255));
    Glb2LocalMux I__4049 (
            .O(N__18437),
            .I(N__18255));
    Glb2LocalMux I__4048 (
            .O(N__18434),
            .I(N__18255));
    CEMux I__4047 (
            .O(N__18433),
            .I(N__18255));
    Glb2LocalMux I__4046 (
            .O(N__18430),
            .I(N__18255));
    Glb2LocalMux I__4045 (
            .O(N__18427),
            .I(N__18255));
    Glb2LocalMux I__4044 (
            .O(N__18424),
            .I(N__18255));
    Glb2LocalMux I__4043 (
            .O(N__18421),
            .I(N__18255));
    Glb2LocalMux I__4042 (
            .O(N__18418),
            .I(N__18255));
    Glb2LocalMux I__4041 (
            .O(N__18415),
            .I(N__18255));
    Glb2LocalMux I__4040 (
            .O(N__18412),
            .I(N__18255));
    Glb2LocalMux I__4039 (
            .O(N__18409),
            .I(N__18255));
    Glb2LocalMux I__4038 (
            .O(N__18406),
            .I(N__18255));
    Glb2LocalMux I__4037 (
            .O(N__18403),
            .I(N__18255));
    Glb2LocalMux I__4036 (
            .O(N__18400),
            .I(N__18255));
    Glb2LocalMux I__4035 (
            .O(N__18397),
            .I(N__18255));
    Glb2LocalMux I__4034 (
            .O(N__18394),
            .I(N__18255));
    Glb2LocalMux I__4033 (
            .O(N__18391),
            .I(N__18255));
    Glb2LocalMux I__4032 (
            .O(N__18388),
            .I(N__18255));
    Glb2LocalMux I__4031 (
            .O(N__18385),
            .I(N__18255));
    Glb2LocalMux I__4030 (
            .O(N__18382),
            .I(N__18255));
    Glb2LocalMux I__4029 (
            .O(N__18379),
            .I(N__18255));
    Glb2LocalMux I__4028 (
            .O(N__18376),
            .I(N__18255));
    Glb2LocalMux I__4027 (
            .O(N__18373),
            .I(N__18255));
    Glb2LocalMux I__4026 (
            .O(N__18370),
            .I(N__18255));
    Glb2LocalMux I__4025 (
            .O(N__18367),
            .I(N__18255));
    Glb2LocalMux I__4024 (
            .O(N__18364),
            .I(N__18255));
    GlobalMux I__4023 (
            .O(N__18255),
            .I(N__18252));
    gio2CtrlBuf I__4022 (
            .O(N__18252),
            .I(N_49_g));
    CascadeMux I__4021 (
            .O(N__18249),
            .I(\ALL_SYS_PWRGD.un4_count_9_cascade_ ));
    InMux I__4020 (
            .O(N__18246),
            .I(N__18243));
    LocalMux I__4019 (
            .O(N__18243),
            .I(N__18239));
    InMux I__4018 (
            .O(N__18242),
            .I(N__18236));
    Odrv4 I__4017 (
            .O(N__18239),
            .I(\ALL_SYS_PWRGD.N_1_i ));
    LocalMux I__4016 (
            .O(N__18236),
            .I(\ALL_SYS_PWRGD.N_1_i ));
    InMux I__4015 (
            .O(N__18231),
            .I(N__18227));
    InMux I__4014 (
            .O(N__18230),
            .I(N__18224));
    LocalMux I__4013 (
            .O(N__18227),
            .I(\ALL_SYS_PWRGD.countZ0Z_7 ));
    LocalMux I__4012 (
            .O(N__18224),
            .I(\ALL_SYS_PWRGD.countZ0Z_7 ));
    InMux I__4011 (
            .O(N__18219),
            .I(N__18215));
    InMux I__4010 (
            .O(N__18218),
            .I(N__18212));
    LocalMux I__4009 (
            .O(N__18215),
            .I(\ALL_SYS_PWRGD.countZ0Z_6 ));
    LocalMux I__4008 (
            .O(N__18212),
            .I(\ALL_SYS_PWRGD.countZ0Z_6 ));
    CascadeMux I__4007 (
            .O(N__18207),
            .I(N__18203));
    InMux I__4006 (
            .O(N__18206),
            .I(N__18200));
    InMux I__4005 (
            .O(N__18203),
            .I(N__18197));
    LocalMux I__4004 (
            .O(N__18200),
            .I(\ALL_SYS_PWRGD.countZ0Z_8 ));
    LocalMux I__4003 (
            .O(N__18197),
            .I(\ALL_SYS_PWRGD.countZ0Z_8 ));
    InMux I__4002 (
            .O(N__18192),
            .I(N__18188));
    InMux I__4001 (
            .O(N__18191),
            .I(N__18185));
    LocalMux I__4000 (
            .O(N__18188),
            .I(\ALL_SYS_PWRGD.countZ0Z_4 ));
    LocalMux I__3999 (
            .O(N__18185),
            .I(\ALL_SYS_PWRGD.countZ0Z_4 ));
    InMux I__3998 (
            .O(N__18180),
            .I(N__18177));
    LocalMux I__3997 (
            .O(N__18177),
            .I(\ALL_SYS_PWRGD.un4_count_8 ));
    InMux I__3996 (
            .O(N__18174),
            .I(N__18170));
    InMux I__3995 (
            .O(N__18173),
            .I(N__18167));
    LocalMux I__3994 (
            .O(N__18170),
            .I(\ALL_SYS_PWRGD.countZ0Z_3 ));
    LocalMux I__3993 (
            .O(N__18167),
            .I(\ALL_SYS_PWRGD.countZ0Z_3 ));
    InMux I__3992 (
            .O(N__18162),
            .I(N__18158));
    InMux I__3991 (
            .O(N__18161),
            .I(N__18155));
    LocalMux I__3990 (
            .O(N__18158),
            .I(\ALL_SYS_PWRGD.countZ0Z_11 ));
    LocalMux I__3989 (
            .O(N__18155),
            .I(\ALL_SYS_PWRGD.countZ0Z_11 ));
    CascadeMux I__3988 (
            .O(N__18150),
            .I(N__18146));
    InMux I__3987 (
            .O(N__18149),
            .I(N__18143));
    InMux I__3986 (
            .O(N__18146),
            .I(N__18140));
    LocalMux I__3985 (
            .O(N__18143),
            .I(\ALL_SYS_PWRGD.countZ0Z_5 ));
    LocalMux I__3984 (
            .O(N__18140),
            .I(\ALL_SYS_PWRGD.countZ0Z_5 ));
    InMux I__3983 (
            .O(N__18135),
            .I(N__18131));
    InMux I__3982 (
            .O(N__18134),
            .I(N__18128));
    LocalMux I__3981 (
            .O(N__18131),
            .I(\ALL_SYS_PWRGD.countZ0Z_2 ));
    LocalMux I__3980 (
            .O(N__18128),
            .I(\ALL_SYS_PWRGD.countZ0Z_2 ));
    InMux I__3979 (
            .O(N__18123),
            .I(N__18120));
    LocalMux I__3978 (
            .O(N__18120),
            .I(\ALL_SYS_PWRGD.un4_count_10 ));
    InMux I__3977 (
            .O(N__18117),
            .I(N__18114));
    LocalMux I__3976 (
            .O(N__18114),
            .I(N__18111));
    Span4Mux_v I__3975 (
            .O(N__18111),
            .I(N__18107));
    InMux I__3974 (
            .O(N__18110),
            .I(N__18104));
    Span4Mux_v I__3973 (
            .O(N__18107),
            .I(N__18101));
    LocalMux I__3972 (
            .O(N__18104),
            .I(N__18098));
    Odrv4 I__3971 (
            .O(N__18101),
            .I(vddq_ok));
    Odrv4 I__3970 (
            .O(N__18098),
            .I(vddq_ok));
    InMux I__3969 (
            .O(N__18093),
            .I(N__18090));
    LocalMux I__3968 (
            .O(N__18090),
            .I(v5s_ok));
    InMux I__3967 (
            .O(N__18087),
            .I(N__18084));
    LocalMux I__3966 (
            .O(N__18084),
            .I(N__18081));
    Span4Mux_v I__3965 (
            .O(N__18081),
            .I(N__18078));
    Odrv4 I__3964 (
            .O(N__18078),
            .I(vccst_cpu_ok));
    InMux I__3963 (
            .O(N__18075),
            .I(N__18072));
    LocalMux I__3962 (
            .O(N__18072),
            .I(N__18066));
    InMux I__3961 (
            .O(N__18071),
            .I(N__18061));
    InMux I__3960 (
            .O(N__18070),
            .I(N__18061));
    InMux I__3959 (
            .O(N__18069),
            .I(N__18058));
    Span12Mux_s4_h I__3958 (
            .O(N__18066),
            .I(N__18055));
    LocalMux I__3957 (
            .O(N__18061),
            .I(N__18052));
    LocalMux I__3956 (
            .O(N__18058),
            .I(N__18049));
    Odrv12 I__3955 (
            .O(N__18055),
            .I(rsmrst_pwrgd_signal));
    Odrv4 I__3954 (
            .O(N__18052),
            .I(rsmrst_pwrgd_signal));
    Odrv4 I__3953 (
            .O(N__18049),
            .I(rsmrst_pwrgd_signal));
    CascadeMux I__3952 (
            .O(N__18042),
            .I(\ALL_SYS_PWRGD.m4_0_0_a2_1_cascade_ ));
    InMux I__3951 (
            .O(N__18039),
            .I(N__18036));
    LocalMux I__3950 (
            .O(N__18036),
            .I(N__18033));
    Span12Mux_v I__3949 (
            .O(N__18033),
            .I(N__18030));
    Odrv12 I__3948 (
            .O(N__18030),
            .I(v33s_ok));
    InMux I__3947 (
            .O(N__18027),
            .I(N__18024));
    LocalMux I__3946 (
            .O(N__18024),
            .I(N__18020));
    InMux I__3945 (
            .O(N__18023),
            .I(N__18016));
    Span4Mux_v I__3944 (
            .O(N__18020),
            .I(N__18012));
    InMux I__3943 (
            .O(N__18019),
            .I(N__18009));
    LocalMux I__3942 (
            .O(N__18016),
            .I(N__18006));
    InMux I__3941 (
            .O(N__18015),
            .I(N__18003));
    Odrv4 I__3940 (
            .O(N__18012),
            .I(\ALL_SYS_PWRGD.N_245 ));
    LocalMux I__3939 (
            .O(N__18009),
            .I(\ALL_SYS_PWRGD.N_245 ));
    Odrv4 I__3938 (
            .O(N__18006),
            .I(\ALL_SYS_PWRGD.N_245 ));
    LocalMux I__3937 (
            .O(N__18003),
            .I(\ALL_SYS_PWRGD.N_245 ));
    InMux I__3936 (
            .O(N__17994),
            .I(N__17990));
    InMux I__3935 (
            .O(N__17993),
            .I(N__17987));
    LocalMux I__3934 (
            .O(N__17990),
            .I(\ALL_SYS_PWRGD.countZ0Z_14 ));
    LocalMux I__3933 (
            .O(N__17987),
            .I(\ALL_SYS_PWRGD.countZ0Z_14 ));
    InMux I__3932 (
            .O(N__17982),
            .I(N__17978));
    InMux I__3931 (
            .O(N__17981),
            .I(N__17975));
    LocalMux I__3930 (
            .O(N__17978),
            .I(\ALL_SYS_PWRGD.countZ0Z_13 ));
    LocalMux I__3929 (
            .O(N__17975),
            .I(\ALL_SYS_PWRGD.countZ0Z_13 ));
    CascadeMux I__3928 (
            .O(N__17970),
            .I(N__17966));
    InMux I__3927 (
            .O(N__17969),
            .I(N__17963));
    InMux I__3926 (
            .O(N__17966),
            .I(N__17960));
    LocalMux I__3925 (
            .O(N__17963),
            .I(\ALL_SYS_PWRGD.countZ0Z_15 ));
    LocalMux I__3924 (
            .O(N__17960),
            .I(\ALL_SYS_PWRGD.countZ0Z_15 ));
    InMux I__3923 (
            .O(N__17955),
            .I(N__17951));
    InMux I__3922 (
            .O(N__17954),
            .I(N__17948));
    LocalMux I__3921 (
            .O(N__17951),
            .I(\ALL_SYS_PWRGD.countZ0Z_12 ));
    LocalMux I__3920 (
            .O(N__17948),
            .I(\ALL_SYS_PWRGD.countZ0Z_12 ));
    InMux I__3919 (
            .O(N__17943),
            .I(N__17940));
    LocalMux I__3918 (
            .O(N__17940),
            .I(N__17937));
    Odrv4 I__3917 (
            .O(N__17937),
            .I(\ALL_SYS_PWRGD.un4_count_11 ));
    SRMux I__3916 (
            .O(N__17934),
            .I(N__17930));
    SRMux I__3915 (
            .O(N__17933),
            .I(N__17927));
    LocalMux I__3914 (
            .O(N__17930),
            .I(N__17922));
    LocalMux I__3913 (
            .O(N__17927),
            .I(N__17919));
    SRMux I__3912 (
            .O(N__17926),
            .I(N__17916));
    InMux I__3911 (
            .O(N__17925),
            .I(N__17913));
    Span4Mux_s1_h I__3910 (
            .O(N__17922),
            .I(N__17910));
    Sp12to4 I__3909 (
            .O(N__17919),
            .I(N__17905));
    LocalMux I__3908 (
            .O(N__17916),
            .I(N__17905));
    LocalMux I__3907 (
            .O(N__17913),
            .I(N__17902));
    Odrv4 I__3906 (
            .O(N__17910),
            .I(\ALL_SYS_PWRGD.curr_state_RNIDP9H7Z0Z_1 ));
    Odrv12 I__3905 (
            .O(N__17905),
            .I(\ALL_SYS_PWRGD.curr_state_RNIDP9H7Z0Z_1 ));
    Odrv4 I__3904 (
            .O(N__17902),
            .I(\ALL_SYS_PWRGD.curr_state_RNIDP9H7Z0Z_1 ));
    CEMux I__3903 (
            .O(N__17895),
            .I(N__17892));
    LocalMux I__3902 (
            .O(N__17892),
            .I(N__17889));
    Span4Mux_v I__3901 (
            .O(N__17889),
            .I(N__17886));
    Span4Mux_s0_h I__3900 (
            .O(N__17886),
            .I(N__17883));
    Odrv4 I__3899 (
            .O(N__17883),
            .I(\ALL_SYS_PWRGD.N_49_4 ));
    InMux I__3898 (
            .O(N__17880),
            .I(N__17876));
    InMux I__3897 (
            .O(N__17879),
            .I(N__17873));
    LocalMux I__3896 (
            .O(N__17876),
            .I(N__17868));
    LocalMux I__3895 (
            .O(N__17873),
            .I(N__17868));
    Span4Mux_s2_h I__3894 (
            .O(N__17868),
            .I(N__17865));
    Odrv4 I__3893 (
            .O(N__17865),
            .I(\POWERLED.N_48 ));
    CascadeMux I__3892 (
            .O(N__17862),
            .I(N__17857));
    CascadeMux I__3891 (
            .O(N__17861),
            .I(N__17854));
    InMux I__3890 (
            .O(N__17860),
            .I(N__17851));
    InMux I__3889 (
            .O(N__17857),
            .I(N__17848));
    InMux I__3888 (
            .O(N__17854),
            .I(N__17845));
    LocalMux I__3887 (
            .O(N__17851),
            .I(N__17842));
    LocalMux I__3886 (
            .O(N__17848),
            .I(\POWERLED.count_offZ0Z_0 ));
    LocalMux I__3885 (
            .O(N__17845),
            .I(\POWERLED.count_offZ0Z_0 ));
    Odrv4 I__3884 (
            .O(N__17842),
            .I(\POWERLED.count_offZ0Z_0 ));
    InMux I__3883 (
            .O(N__17835),
            .I(N__17831));
    InMux I__3882 (
            .O(N__17834),
            .I(N__17828));
    LocalMux I__3881 (
            .O(N__17831),
            .I(\POWERLED.count_offZ0Z_9 ));
    LocalMux I__3880 (
            .O(N__17828),
            .I(\POWERLED.count_offZ0Z_9 ));
    CascadeMux I__3879 (
            .O(N__17823),
            .I(N__17819));
    InMux I__3878 (
            .O(N__17822),
            .I(N__17816));
    InMux I__3877 (
            .O(N__17819),
            .I(N__17813));
    LocalMux I__3876 (
            .O(N__17816),
            .I(\POWERLED.count_offZ0Z_8 ));
    LocalMux I__3875 (
            .O(N__17813),
            .I(\POWERLED.count_offZ0Z_8 ));
    InMux I__3874 (
            .O(N__17808),
            .I(N__17805));
    LocalMux I__3873 (
            .O(N__17805),
            .I(\POWERLED.func_state_ns_0_a2_9_0 ));
    InMux I__3872 (
            .O(N__17802),
            .I(N__17798));
    InMux I__3871 (
            .O(N__17801),
            .I(N__17795));
    LocalMux I__3870 (
            .O(N__17798),
            .I(\POWERLED.count_offZ0Z_10 ));
    LocalMux I__3869 (
            .O(N__17795),
            .I(\POWERLED.count_offZ0Z_10 ));
    InMux I__3868 (
            .O(N__17790),
            .I(N__17786));
    InMux I__3867 (
            .O(N__17789),
            .I(N__17783));
    LocalMux I__3866 (
            .O(N__17786),
            .I(N__17780));
    LocalMux I__3865 (
            .O(N__17783),
            .I(\POWERLED.count_offZ0Z_14 ));
    Odrv4 I__3864 (
            .O(N__17780),
            .I(\POWERLED.count_offZ0Z_14 ));
    CascadeMux I__3863 (
            .O(N__17775),
            .I(N__17771));
    InMux I__3862 (
            .O(N__17774),
            .I(N__17768));
    InMux I__3861 (
            .O(N__17771),
            .I(N__17765));
    LocalMux I__3860 (
            .O(N__17768),
            .I(\POWERLED.count_offZ0Z_11 ));
    LocalMux I__3859 (
            .O(N__17765),
            .I(\POWERLED.count_offZ0Z_11 ));
    InMux I__3858 (
            .O(N__17760),
            .I(N__17757));
    LocalMux I__3857 (
            .O(N__17757),
            .I(\POWERLED.func_state_ns_0_a2_10_0 ));
    InMux I__3856 (
            .O(N__17754),
            .I(N__17750));
    InMux I__3855 (
            .O(N__17753),
            .I(N__17747));
    LocalMux I__3854 (
            .O(N__17750),
            .I(\POWERLED.count_offZ0Z_13 ));
    LocalMux I__3853 (
            .O(N__17747),
            .I(\POWERLED.count_offZ0Z_13 ));
    InMux I__3852 (
            .O(N__17742),
            .I(N__17738));
    InMux I__3851 (
            .O(N__17741),
            .I(N__17735));
    LocalMux I__3850 (
            .O(N__17738),
            .I(\POWERLED.count_offZ0Z_12 ));
    LocalMux I__3849 (
            .O(N__17735),
            .I(\POWERLED.count_offZ0Z_12 ));
    CascadeMux I__3848 (
            .O(N__17730),
            .I(N__17726));
    InMux I__3847 (
            .O(N__17729),
            .I(N__17723));
    InMux I__3846 (
            .O(N__17726),
            .I(N__17720));
    LocalMux I__3845 (
            .O(N__17723),
            .I(\POWERLED.count_offZ0Z_15 ));
    LocalMux I__3844 (
            .O(N__17720),
            .I(\POWERLED.count_offZ0Z_15 ));
    InMux I__3843 (
            .O(N__17715),
            .I(N__17711));
    InMux I__3842 (
            .O(N__17714),
            .I(N__17708));
    LocalMux I__3841 (
            .O(N__17711),
            .I(N__17705));
    LocalMux I__3840 (
            .O(N__17708),
            .I(\POWERLED.count_offZ0Z_1 ));
    Odrv4 I__3839 (
            .O(N__17705),
            .I(\POWERLED.count_offZ0Z_1 ));
    InMux I__3838 (
            .O(N__17700),
            .I(N__17697));
    LocalMux I__3837 (
            .O(N__17697),
            .I(\POWERLED.func_state_ns_0_a2_11_0 ));
    InMux I__3836 (
            .O(N__17694),
            .I(N__17691));
    LocalMux I__3835 (
            .O(N__17691),
            .I(N__17688));
    Span12Mux_s6_h I__3834 (
            .O(N__17688),
            .I(N__17684));
    InMux I__3833 (
            .O(N__17687),
            .I(N__17681));
    Odrv12 I__3832 (
            .O(N__17684),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    LocalMux I__3831 (
            .O(N__17681),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    InMux I__3830 (
            .O(N__17676),
            .I(N__17671));
    InMux I__3829 (
            .O(N__17675),
            .I(N__17667));
    InMux I__3828 (
            .O(N__17674),
            .I(N__17663));
    LocalMux I__3827 (
            .O(N__17671),
            .I(N__17660));
    InMux I__3826 (
            .O(N__17670),
            .I(N__17657));
    LocalMux I__3825 (
            .O(N__17667),
            .I(N__17654));
    CascadeMux I__3824 (
            .O(N__17666),
            .I(N__17650));
    LocalMux I__3823 (
            .O(N__17663),
            .I(N__17646));
    Span4Mux_v I__3822 (
            .O(N__17660),
            .I(N__17641));
    LocalMux I__3821 (
            .O(N__17657),
            .I(N__17641));
    Span4Mux_v I__3820 (
            .O(N__17654),
            .I(N__17638));
    InMux I__3819 (
            .O(N__17653),
            .I(N__17635));
    InMux I__3818 (
            .O(N__17650),
            .I(N__17630));
    InMux I__3817 (
            .O(N__17649),
            .I(N__17630));
    Span4Mux_v I__3816 (
            .O(N__17646),
            .I(N__17627));
    Span4Mux_h I__3815 (
            .O(N__17641),
            .I(N__17624));
    Sp12to4 I__3814 (
            .O(N__17638),
            .I(N__17617));
    LocalMux I__3813 (
            .O(N__17635),
            .I(N__17617));
    LocalMux I__3812 (
            .O(N__17630),
            .I(N__17617));
    Odrv4 I__3811 (
            .O(N__17627),
            .I(N_55));
    Odrv4 I__3810 (
            .O(N__17624),
            .I(N_55));
    Odrv12 I__3809 (
            .O(N__17617),
            .I(N_55));
    IoInMux I__3808 (
            .O(N__17610),
            .I(N__17607));
    LocalMux I__3807 (
            .O(N__17607),
            .I(N__17604));
    Odrv4 I__3806 (
            .O(N__17604),
            .I(vpp_en));
    InMux I__3805 (
            .O(N__17601),
            .I(N__17598));
    LocalMux I__3804 (
            .O(N__17598),
            .I(\ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa ));
    InMux I__3803 (
            .O(N__17595),
            .I(N__17585));
    InMux I__3802 (
            .O(N__17594),
            .I(N__17585));
    InMux I__3801 (
            .O(N__17593),
            .I(N__17582));
    InMux I__3800 (
            .O(N__17592),
            .I(N__17579));
    InMux I__3799 (
            .O(N__17591),
            .I(N__17576));
    InMux I__3798 (
            .O(N__17590),
            .I(N__17573));
    LocalMux I__3797 (
            .O(N__17585),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__3796 (
            .O(N__17582),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__3795 (
            .O(N__17579),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__3794 (
            .O(N__17576),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__3793 (
            .O(N__17573),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__3792 (
            .O(N__17562),
            .I(N__17558));
    InMux I__3791 (
            .O(N__17561),
            .I(N__17549));
    InMux I__3790 (
            .O(N__17558),
            .I(N__17549));
    InMux I__3789 (
            .O(N__17557),
            .I(N__17546));
    InMux I__3788 (
            .O(N__17556),
            .I(N__17543));
    InMux I__3787 (
            .O(N__17555),
            .I(N__17538));
    InMux I__3786 (
            .O(N__17554),
            .I(N__17538));
    LocalMux I__3785 (
            .O(N__17549),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__3784 (
            .O(N__17546),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__3783 (
            .O(N__17543),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__3782 (
            .O(N__17538),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_0 ));
    CascadeMux I__3781 (
            .O(N__17529),
            .I(N__17525));
    InMux I__3780 (
            .O(N__17528),
            .I(N__17522));
    InMux I__3779 (
            .O(N__17525),
            .I(N__17519));
    LocalMux I__3778 (
            .O(N__17522),
            .I(\ALL_SYS_PWRGD.un1_curr_state10_0 ));
    LocalMux I__3777 (
            .O(N__17519),
            .I(\ALL_SYS_PWRGD.un1_curr_state10_0 ));
    InMux I__3776 (
            .O(N__17514),
            .I(N__17510));
    InMux I__3775 (
            .O(N__17513),
            .I(N__17507));
    LocalMux I__3774 (
            .O(N__17510),
            .I(\ALL_SYS_PWRGD.countZ0Z_9 ));
    LocalMux I__3773 (
            .O(N__17507),
            .I(\ALL_SYS_PWRGD.countZ0Z_9 ));
    InMux I__3772 (
            .O(N__17502),
            .I(N__17498));
    InMux I__3771 (
            .O(N__17501),
            .I(N__17495));
    LocalMux I__3770 (
            .O(N__17498),
            .I(\ALL_SYS_PWRGD.countZ0Z_1 ));
    LocalMux I__3769 (
            .O(N__17495),
            .I(\ALL_SYS_PWRGD.countZ0Z_1 ));
    CascadeMux I__3768 (
            .O(N__17490),
            .I(N__17486));
    InMux I__3767 (
            .O(N__17489),
            .I(N__17483));
    InMux I__3766 (
            .O(N__17486),
            .I(N__17480));
    LocalMux I__3765 (
            .O(N__17483),
            .I(\ALL_SYS_PWRGD.countZ0Z_10 ));
    LocalMux I__3764 (
            .O(N__17480),
            .I(\ALL_SYS_PWRGD.countZ0Z_10 ));
    InMux I__3763 (
            .O(N__17475),
            .I(N__17471));
    InMux I__3762 (
            .O(N__17474),
            .I(N__17468));
    LocalMux I__3761 (
            .O(N__17471),
            .I(\ALL_SYS_PWRGD.countZ0Z_0 ));
    LocalMux I__3760 (
            .O(N__17468),
            .I(\ALL_SYS_PWRGD.countZ0Z_0 ));
    InMux I__3759 (
            .O(N__17463),
            .I(\POWERLED.un1_count_off_1_cry_8 ));
    InMux I__3758 (
            .O(N__17460),
            .I(\POWERLED.un1_count_off_1_cry_9 ));
    InMux I__3757 (
            .O(N__17457),
            .I(\POWERLED.un1_count_off_1_cry_10 ));
    InMux I__3756 (
            .O(N__17454),
            .I(\POWERLED.un1_count_off_1_cry_11 ));
    InMux I__3755 (
            .O(N__17451),
            .I(\POWERLED.un1_count_off_1_cry_12 ));
    InMux I__3754 (
            .O(N__17448),
            .I(\POWERLED.un1_count_off_1_cry_13 ));
    InMux I__3753 (
            .O(N__17445),
            .I(\POWERLED.un1_count_off_1_cry_14 ));
    InMux I__3752 (
            .O(N__17442),
            .I(N__17438));
    InMux I__3751 (
            .O(N__17441),
            .I(N__17435));
    LocalMux I__3750 (
            .O(N__17438),
            .I(N__17432));
    LocalMux I__3749 (
            .O(N__17435),
            .I(\POWERLED.count_offZ0Z_4 ));
    Odrv4 I__3748 (
            .O(N__17432),
            .I(\POWERLED.count_offZ0Z_4 ));
    CascadeMux I__3747 (
            .O(N__17427),
            .I(N__17424));
    InMux I__3746 (
            .O(N__17424),
            .I(N__17420));
    InMux I__3745 (
            .O(N__17423),
            .I(N__17417));
    LocalMux I__3744 (
            .O(N__17420),
            .I(N__17414));
    LocalMux I__3743 (
            .O(N__17417),
            .I(\POWERLED.count_offZ0Z_7 ));
    Odrv4 I__3742 (
            .O(N__17414),
            .I(\POWERLED.count_offZ0Z_7 ));
    InMux I__3741 (
            .O(N__17409),
            .I(N__17405));
    InMux I__3740 (
            .O(N__17408),
            .I(N__17402));
    LocalMux I__3739 (
            .O(N__17405),
            .I(N__17399));
    LocalMux I__3738 (
            .O(N__17402),
            .I(\POWERLED.count_offZ0Z_3 ));
    Odrv4 I__3737 (
            .O(N__17399),
            .I(\POWERLED.count_offZ0Z_3 ));
    CascadeMux I__3736 (
            .O(N__17394),
            .I(\POWERLED.func_state_ns_0_a2_8_0_cascade_ ));
    InMux I__3735 (
            .O(N__17391),
            .I(N__17384));
    InMux I__3734 (
            .O(N__17390),
            .I(N__17381));
    InMux I__3733 (
            .O(N__17389),
            .I(N__17374));
    InMux I__3732 (
            .O(N__17388),
            .I(N__17374));
    InMux I__3731 (
            .O(N__17387),
            .I(N__17374));
    LocalMux I__3730 (
            .O(N__17384),
            .I(N__17363));
    LocalMux I__3729 (
            .O(N__17381),
            .I(N__17363));
    LocalMux I__3728 (
            .O(N__17374),
            .I(N__17363));
    InMux I__3727 (
            .O(N__17373),
            .I(N__17354));
    InMux I__3726 (
            .O(N__17372),
            .I(N__17354));
    InMux I__3725 (
            .O(N__17371),
            .I(N__17354));
    InMux I__3724 (
            .O(N__17370),
            .I(N__17354));
    Span4Mux_v I__3723 (
            .O(N__17363),
            .I(N__17349));
    LocalMux I__3722 (
            .O(N__17354),
            .I(N__17349));
    Odrv4 I__3721 (
            .O(N__17349),
            .I(\POWERLED.count_off_RNIIKVR3Z0Z_10 ));
    InMux I__3720 (
            .O(N__17346),
            .I(\POWERLED.un1_count_off_1_cry_0 ));
    InMux I__3719 (
            .O(N__17343),
            .I(\POWERLED.un1_count_off_1_cry_1 ));
    InMux I__3718 (
            .O(N__17340),
            .I(\POWERLED.un1_count_off_1_cry_2 ));
    InMux I__3717 (
            .O(N__17337),
            .I(\POWERLED.un1_count_off_1_cry_3 ));
    InMux I__3716 (
            .O(N__17334),
            .I(\POWERLED.un1_count_off_1_cry_4 ));
    InMux I__3715 (
            .O(N__17331),
            .I(\POWERLED.un1_count_off_1_cry_5 ));
    InMux I__3714 (
            .O(N__17328),
            .I(\POWERLED.un1_count_off_1_cry_6 ));
    InMux I__3713 (
            .O(N__17325),
            .I(bfn_11_11_0_));
    InMux I__3712 (
            .O(N__17322),
            .I(bfn_11_8_0_));
    InMux I__3711 (
            .O(N__17319),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_8 ));
    InMux I__3710 (
            .O(N__17316),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_9 ));
    InMux I__3709 (
            .O(N__17313),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_10 ));
    InMux I__3708 (
            .O(N__17310),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_11 ));
    InMux I__3707 (
            .O(N__17307),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_12 ));
    InMux I__3706 (
            .O(N__17304),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_13 ));
    CascadeMux I__3705 (
            .O(N__17301),
            .I(N__17294));
    IoInMux I__3704 (
            .O(N__17300),
            .I(N__17289));
    CascadeMux I__3703 (
            .O(N__17299),
            .I(N__17285));
    InMux I__3702 (
            .O(N__17298),
            .I(N__17282));
    InMux I__3701 (
            .O(N__17297),
            .I(N__17279));
    InMux I__3700 (
            .O(N__17294),
            .I(N__17273));
    InMux I__3699 (
            .O(N__17293),
            .I(N__17273));
    InMux I__3698 (
            .O(N__17292),
            .I(N__17270));
    LocalMux I__3697 (
            .O(N__17289),
            .I(N__17267));
    InMux I__3696 (
            .O(N__17288),
            .I(N__17261));
    InMux I__3695 (
            .O(N__17285),
            .I(N__17261));
    LocalMux I__3694 (
            .O(N__17282),
            .I(N__17257));
    LocalMux I__3693 (
            .O(N__17279),
            .I(N__17254));
    InMux I__3692 (
            .O(N__17278),
            .I(N__17251));
    LocalMux I__3691 (
            .O(N__17273),
            .I(N__17248));
    LocalMux I__3690 (
            .O(N__17270),
            .I(N__17245));
    IoSpan4Mux I__3689 (
            .O(N__17267),
            .I(N__17242));
    InMux I__3688 (
            .O(N__17266),
            .I(N__17239));
    LocalMux I__3687 (
            .O(N__17261),
            .I(N__17236));
    InMux I__3686 (
            .O(N__17260),
            .I(N__17233));
    Span4Mux_h I__3685 (
            .O(N__17257),
            .I(N__17227));
    Span4Mux_v I__3684 (
            .O(N__17254),
            .I(N__17227));
    LocalMux I__3683 (
            .O(N__17251),
            .I(N__17224));
    Span4Mux_h I__3682 (
            .O(N__17248),
            .I(N__17219));
    Span4Mux_s3_v I__3681 (
            .O(N__17245),
            .I(N__17219));
    Span4Mux_s3_h I__3680 (
            .O(N__17242),
            .I(N__17214));
    LocalMux I__3679 (
            .O(N__17239),
            .I(N__17214));
    Span4Mux_v I__3678 (
            .O(N__17236),
            .I(N__17209));
    LocalMux I__3677 (
            .O(N__17233),
            .I(N__17209));
    InMux I__3676 (
            .O(N__17232),
            .I(N__17206));
    Span4Mux_h I__3675 (
            .O(N__17227),
            .I(N__17201));
    Span4Mux_v I__3674 (
            .O(N__17224),
            .I(N__17201));
    Span4Mux_v I__3673 (
            .O(N__17219),
            .I(N__17192));
    Span4Mux_h I__3672 (
            .O(N__17214),
            .I(N__17192));
    Span4Mux_h I__3671 (
            .O(N__17209),
            .I(N__17192));
    LocalMux I__3670 (
            .O(N__17206),
            .I(N__17192));
    Odrv4 I__3669 (
            .O(N__17201),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3668 (
            .O(N__17192),
            .I(CONSTANT_ONE_NET));
    InMux I__3667 (
            .O(N__17187),
            .I(bfn_11_9_0_));
    InMux I__3666 (
            .O(N__17184),
            .I(N__17180));
    InMux I__3665 (
            .O(N__17183),
            .I(N__17177));
    LocalMux I__3664 (
            .O(N__17180),
            .I(\ALL_SYS_PWRGD.N_247 ));
    LocalMux I__3663 (
            .O(N__17177),
            .I(\ALL_SYS_PWRGD.N_247 ));
    CascadeMux I__3662 (
            .O(N__17172),
            .I(\ALL_SYS_PWRGD.N_186_cascade_ ));
    InMux I__3661 (
            .O(N__17169),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_0 ));
    InMux I__3660 (
            .O(N__17166),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_1 ));
    InMux I__3659 (
            .O(N__17163),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_2 ));
    InMux I__3658 (
            .O(N__17160),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_3 ));
    InMux I__3657 (
            .O(N__17157),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_4 ));
    InMux I__3656 (
            .O(N__17154),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_5 ));
    InMux I__3655 (
            .O(N__17151),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_6 ));
    InMux I__3654 (
            .O(N__17148),
            .I(N__17145));
    LocalMux I__3653 (
            .O(N__17145),
            .I(N__17142));
    Odrv12 I__3652 (
            .O(N__17142),
            .I(\POWERLED.count_clk_137_tz_0 ));
    InMux I__3651 (
            .O(N__17139),
            .I(N__17136));
    LocalMux I__3650 (
            .O(N__17136),
            .I(\POWERLED.un2_slp_s3n_2_0 ));
    InMux I__3649 (
            .O(N__17133),
            .I(N__17129));
    InMux I__3648 (
            .O(N__17132),
            .I(N__17126));
    LocalMux I__3647 (
            .O(N__17129),
            .I(\POWERLED.count_clkZ0Z_11 ));
    LocalMux I__3646 (
            .O(N__17126),
            .I(\POWERLED.count_clkZ0Z_11 ));
    InMux I__3645 (
            .O(N__17121),
            .I(N__17117));
    InMux I__3644 (
            .O(N__17120),
            .I(N__17114));
    LocalMux I__3643 (
            .O(N__17117),
            .I(\POWERLED.count_clkZ0Z_10 ));
    LocalMux I__3642 (
            .O(N__17114),
            .I(\POWERLED.count_clkZ0Z_10 ));
    CascadeMux I__3641 (
            .O(N__17109),
            .I(N__17105));
    InMux I__3640 (
            .O(N__17108),
            .I(N__17102));
    InMux I__3639 (
            .O(N__17105),
            .I(N__17099));
    LocalMux I__3638 (
            .O(N__17102),
            .I(\POWERLED.count_clkZ0Z_12 ));
    LocalMux I__3637 (
            .O(N__17099),
            .I(\POWERLED.count_clkZ0Z_12 ));
    InMux I__3636 (
            .O(N__17094),
            .I(N__17090));
    InMux I__3635 (
            .O(N__17093),
            .I(N__17087));
    LocalMux I__3634 (
            .O(N__17090),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__3633 (
            .O(N__17087),
            .I(\POWERLED.count_clkZ0Z_0 ));
    InMux I__3632 (
            .O(N__17082),
            .I(N__17078));
    InMux I__3631 (
            .O(N__17081),
            .I(N__17075));
    LocalMux I__3630 (
            .O(N__17078),
            .I(N__17072));
    LocalMux I__3629 (
            .O(N__17075),
            .I(\POWERLED.count_clkZ0Z_15 ));
    Odrv4 I__3628 (
            .O(N__17072),
            .I(\POWERLED.count_clkZ0Z_15 ));
    InMux I__3627 (
            .O(N__17067),
            .I(N__17063));
    InMux I__3626 (
            .O(N__17066),
            .I(N__17060));
    LocalMux I__3625 (
            .O(N__17063),
            .I(\POWERLED.count_clkZ0Z_14 ));
    LocalMux I__3624 (
            .O(N__17060),
            .I(\POWERLED.count_clkZ0Z_14 ));
    CascadeMux I__3623 (
            .O(N__17055),
            .I(\POWERLED.count_clk_0_sqmuxa_5_0_o2_4_cascade_ ));
    InMux I__3622 (
            .O(N__17052),
            .I(N__17048));
    InMux I__3621 (
            .O(N__17051),
            .I(N__17045));
    LocalMux I__3620 (
            .O(N__17048),
            .I(\POWERLED.count_clkZ0Z_13 ));
    LocalMux I__3619 (
            .O(N__17045),
            .I(\POWERLED.count_clkZ0Z_13 ));
    InMux I__3618 (
            .O(N__17040),
            .I(N__17037));
    LocalMux I__3617 (
            .O(N__17037),
            .I(N__17032));
    InMux I__3616 (
            .O(N__17036),
            .I(N__17027));
    InMux I__3615 (
            .O(N__17035),
            .I(N__17027));
    Odrv4 I__3614 (
            .O(N__17032),
            .I(\POWERLED.N_136 ));
    LocalMux I__3613 (
            .O(N__17027),
            .I(\POWERLED.N_136 ));
    SRMux I__3612 (
            .O(N__17022),
            .I(N__17018));
    SRMux I__3611 (
            .O(N__17021),
            .I(N__17015));
    LocalMux I__3610 (
            .O(N__17018),
            .I(N__17011));
    LocalMux I__3609 (
            .O(N__17015),
            .I(N__17008));
    SRMux I__3608 (
            .O(N__17014),
            .I(N__17005));
    Span4Mux_s2_v I__3607 (
            .O(N__17011),
            .I(N__17001));
    Span4Mux_h I__3606 (
            .O(N__17008),
            .I(N__16996));
    LocalMux I__3605 (
            .O(N__17005),
            .I(N__16996));
    InMux I__3604 (
            .O(N__17004),
            .I(N__16993));
    Odrv4 I__3603 (
            .O(N__17001),
            .I(\POWERLED.count_clk_RNIOH1J11Z0Z_7 ));
    Odrv4 I__3602 (
            .O(N__16996),
            .I(\POWERLED.count_clk_RNIOH1J11Z0Z_7 ));
    LocalMux I__3601 (
            .O(N__16993),
            .I(\POWERLED.count_clk_RNIOH1J11Z0Z_7 ));
    CEMux I__3600 (
            .O(N__16986),
            .I(N__16983));
    LocalMux I__3599 (
            .O(N__16983),
            .I(N__16980));
    Odrv4 I__3598 (
            .O(N__16980),
            .I(\POWERLED.N_49_0 ));
    IoInMux I__3597 (
            .O(N__16977),
            .I(N__16974));
    LocalMux I__3596 (
            .O(N__16974),
            .I(N__16971));
    Span4Mux_s3_v I__3595 (
            .O(N__16971),
            .I(N__16965));
    IoInMux I__3594 (
            .O(N__16970),
            .I(N__16962));
    InMux I__3593 (
            .O(N__16969),
            .I(N__16957));
    InMux I__3592 (
            .O(N__16968),
            .I(N__16957));
    Span4Mux_v I__3591 (
            .O(N__16965),
            .I(N__16954));
    LocalMux I__3590 (
            .O(N__16962),
            .I(N__16951));
    LocalMux I__3589 (
            .O(N__16957),
            .I(N__16948));
    Span4Mux_v I__3588 (
            .O(N__16954),
            .I(N__16945));
    Span12Mux_s4_v I__3587 (
            .O(N__16951),
            .I(N__16942));
    Span4Mux_h I__3586 (
            .O(N__16948),
            .I(N__16939));
    Odrv4 I__3585 (
            .O(N__16945),
            .I(vccst_pwrgd));
    Odrv12 I__3584 (
            .O(N__16942),
            .I(vccst_pwrgd));
    Odrv4 I__3583 (
            .O(N__16939),
            .I(vccst_pwrgd));
    InMux I__3582 (
            .O(N__16932),
            .I(N__16929));
    LocalMux I__3581 (
            .O(N__16929),
            .I(\ALL_SYS_PWRGD.N_186 ));
    InMux I__3580 (
            .O(N__16926),
            .I(N__16923));
    LocalMux I__3579 (
            .O(N__16923),
            .I(\POWERLED.N_207 ));
    InMux I__3578 (
            .O(N__16920),
            .I(N__16917));
    LocalMux I__3577 (
            .O(N__16917),
            .I(\POWERLED.count_off_1_sqmuxa_i_a6_0_3 ));
    IoInMux I__3576 (
            .O(N__16914),
            .I(N__16911));
    LocalMux I__3575 (
            .O(N__16911),
            .I(N__16902));
    InMux I__3574 (
            .O(N__16910),
            .I(N__16899));
    CascadeMux I__3573 (
            .O(N__16909),
            .I(N__16896));
    CascadeMux I__3572 (
            .O(N__16908),
            .I(N__16891));
    InMux I__3571 (
            .O(N__16907),
            .I(N__16884));
    InMux I__3570 (
            .O(N__16906),
            .I(N__16884));
    InMux I__3569 (
            .O(N__16905),
            .I(N__16884));
    IoSpan4Mux I__3568 (
            .O(N__16902),
            .I(N__16881));
    LocalMux I__3567 (
            .O(N__16899),
            .I(N__16878));
    InMux I__3566 (
            .O(N__16896),
            .I(N__16873));
    InMux I__3565 (
            .O(N__16895),
            .I(N__16873));
    InMux I__3564 (
            .O(N__16894),
            .I(N__16868));
    InMux I__3563 (
            .O(N__16891),
            .I(N__16868));
    LocalMux I__3562 (
            .O(N__16884),
            .I(N__16865));
    Span4Mux_s1_h I__3561 (
            .O(N__16881),
            .I(N__16861));
    Span4Mux_v I__3560 (
            .O(N__16878),
            .I(N__16856));
    LocalMux I__3559 (
            .O(N__16873),
            .I(N__16856));
    LocalMux I__3558 (
            .O(N__16868),
            .I(N__16853));
    Span4Mux_h I__3557 (
            .O(N__16865),
            .I(N__16850));
    InMux I__3556 (
            .O(N__16864),
            .I(N__16847));
    Span4Mux_h I__3555 (
            .O(N__16861),
            .I(N__16844));
    Span4Mux_v I__3554 (
            .O(N__16856),
            .I(N__16841));
    Span4Mux_v I__3553 (
            .O(N__16853),
            .I(N__16838));
    Sp12to4 I__3552 (
            .O(N__16850),
            .I(N__16833));
    LocalMux I__3551 (
            .O(N__16847),
            .I(N__16833));
    Span4Mux_h I__3550 (
            .O(N__16844),
            .I(N__16826));
    Span4Mux_v I__3549 (
            .O(N__16841),
            .I(N__16826));
    Span4Mux_v I__3548 (
            .O(N__16838),
            .I(N__16826));
    Span12Mux_v I__3547 (
            .O(N__16833),
            .I(N__16823));
    Odrv4 I__3546 (
            .O(N__16826),
            .I(gpio_fpga_soc_4));
    Odrv12 I__3545 (
            .O(N__16823),
            .I(gpio_fpga_soc_4));
    InMux I__3544 (
            .O(N__16818),
            .I(N__16815));
    LocalMux I__3543 (
            .O(N__16815),
            .I(N__16812));
    Odrv4 I__3542 (
            .O(N__16812),
            .I(\POWERLED.count_off_1_sqmuxa_i_a6_0_1 ));
    InMux I__3541 (
            .O(N__16809),
            .I(N__16804));
    InMux I__3540 (
            .O(N__16808),
            .I(N__16801));
    InMux I__3539 (
            .O(N__16807),
            .I(N__16798));
    LocalMux I__3538 (
            .O(N__16804),
            .I(N__16795));
    LocalMux I__3537 (
            .O(N__16801),
            .I(\POWERLED.N_243 ));
    LocalMux I__3536 (
            .O(N__16798),
            .I(\POWERLED.N_243 ));
    Odrv4 I__3535 (
            .O(N__16795),
            .I(\POWERLED.N_243 ));
    InMux I__3534 (
            .O(N__16788),
            .I(N__16784));
    CascadeMux I__3533 (
            .O(N__16787),
            .I(N__16778));
    LocalMux I__3532 (
            .O(N__16784),
            .I(N__16775));
    IoInMux I__3531 (
            .O(N__16783),
            .I(N__16772));
    InMux I__3530 (
            .O(N__16782),
            .I(N__16769));
    InMux I__3529 (
            .O(N__16781),
            .I(N__16764));
    InMux I__3528 (
            .O(N__16778),
            .I(N__16764));
    Span4Mux_v I__3527 (
            .O(N__16775),
            .I(N__16761));
    LocalMux I__3526 (
            .O(N__16772),
            .I(N__16758));
    LocalMux I__3525 (
            .O(N__16769),
            .I(N__16755));
    LocalMux I__3524 (
            .O(N__16764),
            .I(N__16752));
    Span4Mux_h I__3523 (
            .O(N__16761),
            .I(N__16749));
    Span4Mux_s2_h I__3522 (
            .O(N__16758),
            .I(N__16742));
    Span4Mux_v I__3521 (
            .O(N__16755),
            .I(N__16742));
    Span4Mux_h I__3520 (
            .O(N__16752),
            .I(N__16742));
    Odrv4 I__3519 (
            .O(N__16749),
            .I(vccst_en));
    Odrv4 I__3518 (
            .O(N__16742),
            .I(vccst_en));
    CascadeMux I__3517 (
            .O(N__16737),
            .I(\POWERLED.un2_slp_s3n_2_0_a6_3_0_cascade_ ));
    InMux I__3516 (
            .O(N__16734),
            .I(N__16731));
    LocalMux I__3515 (
            .O(N__16731),
            .I(\POWERLED.un2_slp_s3n_2_0_1_0 ));
    CascadeMux I__3514 (
            .O(N__16728),
            .I(\POWERLED.un2_slp_s3n_2_0_1_cascade_ ));
    InMux I__3513 (
            .O(N__16725),
            .I(N__16722));
    LocalMux I__3512 (
            .O(N__16722),
            .I(N__16718));
    InMux I__3511 (
            .O(N__16721),
            .I(N__16715));
    Span4Mux_h I__3510 (
            .O(N__16718),
            .I(N__16712));
    LocalMux I__3509 (
            .O(N__16715),
            .I(\POWERLED.N_251 ));
    Odrv4 I__3508 (
            .O(N__16712),
            .I(\POWERLED.N_251 ));
    InMux I__3507 (
            .O(N__16707),
            .I(N__16697));
    InMux I__3506 (
            .O(N__16706),
            .I(N__16694));
    CascadeMux I__3505 (
            .O(N__16705),
            .I(N__16690));
    CascadeMux I__3504 (
            .O(N__16704),
            .I(N__16687));
    InMux I__3503 (
            .O(N__16703),
            .I(N__16684));
    InMux I__3502 (
            .O(N__16702),
            .I(N__16681));
    InMux I__3501 (
            .O(N__16701),
            .I(N__16676));
    InMux I__3500 (
            .O(N__16700),
            .I(N__16676));
    LocalMux I__3499 (
            .O(N__16697),
            .I(N__16671));
    LocalMux I__3498 (
            .O(N__16694),
            .I(N__16671));
    InMux I__3497 (
            .O(N__16693),
            .I(N__16664));
    InMux I__3496 (
            .O(N__16690),
            .I(N__16664));
    InMux I__3495 (
            .O(N__16687),
            .I(N__16664));
    LocalMux I__3494 (
            .O(N__16684),
            .I(\POWERLED.count_clkZ0Z_7 ));
    LocalMux I__3493 (
            .O(N__16681),
            .I(\POWERLED.count_clkZ0Z_7 ));
    LocalMux I__3492 (
            .O(N__16676),
            .I(\POWERLED.count_clkZ0Z_7 ));
    Odrv4 I__3491 (
            .O(N__16671),
            .I(\POWERLED.count_clkZ0Z_7 ));
    LocalMux I__3490 (
            .O(N__16664),
            .I(\POWERLED.count_clkZ0Z_7 ));
    InMux I__3489 (
            .O(N__16653),
            .I(N__16650));
    LocalMux I__3488 (
            .O(N__16650),
            .I(\POWERLED.count_clk_0_sqmuxa_5_0_a6_1 ));
    InMux I__3487 (
            .O(N__16647),
            .I(N__16641));
    InMux I__3486 (
            .O(N__16646),
            .I(N__16634));
    InMux I__3485 (
            .O(N__16645),
            .I(N__16634));
    InMux I__3484 (
            .O(N__16644),
            .I(N__16634));
    LocalMux I__3483 (
            .O(N__16641),
            .I(\POWERLED.count_clkZ0Z_5 ));
    LocalMux I__3482 (
            .O(N__16634),
            .I(\POWERLED.count_clkZ0Z_5 ));
    CascadeMux I__3481 (
            .O(N__16629),
            .I(N__16624));
    InMux I__3480 (
            .O(N__16628),
            .I(N__16620));
    InMux I__3479 (
            .O(N__16627),
            .I(N__16613));
    InMux I__3478 (
            .O(N__16624),
            .I(N__16613));
    InMux I__3477 (
            .O(N__16623),
            .I(N__16613));
    LocalMux I__3476 (
            .O(N__16620),
            .I(\POWERLED.count_clkZ0Z_9 ));
    LocalMux I__3475 (
            .O(N__16613),
            .I(\POWERLED.count_clkZ0Z_9 ));
    CascadeMux I__3474 (
            .O(N__16608),
            .I(N__16602));
    InMux I__3473 (
            .O(N__16607),
            .I(N__16599));
    InMux I__3472 (
            .O(N__16606),
            .I(N__16596));
    InMux I__3471 (
            .O(N__16605),
            .I(N__16591));
    InMux I__3470 (
            .O(N__16602),
            .I(N__16591));
    LocalMux I__3469 (
            .O(N__16599),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__3468 (
            .O(N__16596),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__3467 (
            .O(N__16591),
            .I(\POWERLED.count_clkZ0Z_1 ));
    InMux I__3466 (
            .O(N__16584),
            .I(N__16578));
    InMux I__3465 (
            .O(N__16583),
            .I(N__16575));
    InMux I__3464 (
            .O(N__16582),
            .I(N__16570));
    InMux I__3463 (
            .O(N__16581),
            .I(N__16570));
    LocalMux I__3462 (
            .O(N__16578),
            .I(\POWERLED.N_146 ));
    LocalMux I__3461 (
            .O(N__16575),
            .I(\POWERLED.N_146 ));
    LocalMux I__3460 (
            .O(N__16570),
            .I(\POWERLED.N_146 ));
    CascadeMux I__3459 (
            .O(N__16563),
            .I(N__16559));
    InMux I__3458 (
            .O(N__16562),
            .I(N__16551));
    InMux I__3457 (
            .O(N__16559),
            .I(N__16551));
    InMux I__3456 (
            .O(N__16558),
            .I(N__16544));
    InMux I__3455 (
            .O(N__16557),
            .I(N__16544));
    InMux I__3454 (
            .O(N__16556),
            .I(N__16544));
    LocalMux I__3453 (
            .O(N__16551),
            .I(N__16539));
    LocalMux I__3452 (
            .O(N__16544),
            .I(N__16539));
    Odrv12 I__3451 (
            .O(N__16539),
            .I(\VPP_VDDQ.N_238 ));
    InMux I__3450 (
            .O(N__16536),
            .I(N__16532));
    InMux I__3449 (
            .O(N__16535),
            .I(N__16529));
    LocalMux I__3448 (
            .O(N__16532),
            .I(N__16521));
    LocalMux I__3447 (
            .O(N__16529),
            .I(N__16518));
    InMux I__3446 (
            .O(N__16528),
            .I(N__16515));
    InMux I__3445 (
            .O(N__16527),
            .I(N__16512));
    InMux I__3444 (
            .O(N__16526),
            .I(N__16505));
    InMux I__3443 (
            .O(N__16525),
            .I(N__16505));
    InMux I__3442 (
            .O(N__16524),
            .I(N__16505));
    Span4Mux_h I__3441 (
            .O(N__16521),
            .I(N__16502));
    Span4Mux_h I__3440 (
            .O(N__16518),
            .I(N__16497));
    LocalMux I__3439 (
            .O(N__16515),
            .I(N__16497));
    LocalMux I__3438 (
            .O(N__16512),
            .I(N__16494));
    LocalMux I__3437 (
            .O(N__16505),
            .I(N__16491));
    Span4Mux_v I__3436 (
            .O(N__16502),
            .I(N__16488));
    Span4Mux_h I__3435 (
            .O(N__16497),
            .I(N__16485));
    Span4Mux_h I__3434 (
            .O(N__16494),
            .I(N__16480));
    Span4Mux_v I__3433 (
            .O(N__16491),
            .I(N__16480));
    Span4Mux_h I__3432 (
            .O(N__16488),
            .I(N__16477));
    Span4Mux_v I__3431 (
            .O(N__16485),
            .I(N__16474));
    IoSpan4Mux I__3430 (
            .O(N__16480),
            .I(N__16471));
    Odrv4 I__3429 (
            .O(N__16477),
            .I(slp_s3n));
    Odrv4 I__3428 (
            .O(N__16474),
            .I(slp_s3n));
    Odrv4 I__3427 (
            .O(N__16471),
            .I(slp_s3n));
    InMux I__3426 (
            .O(N__16464),
            .I(N__16461));
    LocalMux I__3425 (
            .O(N__16461),
            .I(N__16453));
    InMux I__3424 (
            .O(N__16460),
            .I(N__16448));
    InMux I__3423 (
            .O(N__16459),
            .I(N__16448));
    InMux I__3422 (
            .O(N__16458),
            .I(N__16441));
    InMux I__3421 (
            .O(N__16457),
            .I(N__16441));
    InMux I__3420 (
            .O(N__16456),
            .I(N__16441));
    Span4Mux_v I__3419 (
            .O(N__16453),
            .I(N__16436));
    LocalMux I__3418 (
            .O(N__16448),
            .I(N__16436));
    LocalMux I__3417 (
            .O(N__16441),
            .I(N__16432));
    Span4Mux_h I__3416 (
            .O(N__16436),
            .I(N__16429));
    InMux I__3415 (
            .O(N__16435),
            .I(N__16426));
    Span12Mux_s8_h I__3414 (
            .O(N__16432),
            .I(N__16423));
    Span4Mux_v I__3413 (
            .O(N__16429),
            .I(N__16420));
    LocalMux I__3412 (
            .O(N__16426),
            .I(N__16417));
    Odrv12 I__3411 (
            .O(N__16423),
            .I(slp_s4n));
    Odrv4 I__3410 (
            .O(N__16420),
            .I(slp_s4n));
    Odrv12 I__3409 (
            .O(N__16417),
            .I(slp_s4n));
    InMux I__3408 (
            .O(N__16410),
            .I(N__16407));
    LocalMux I__3407 (
            .O(N__16407),
            .I(N__16404));
    Span4Mux_h I__3406 (
            .O(N__16404),
            .I(N__16401));
    Odrv4 I__3405 (
            .O(N__16401),
            .I(\POWERLED.dutycycle_lm_0_1_2 ));
    InMux I__3404 (
            .O(N__16398),
            .I(N__16392));
    InMux I__3403 (
            .O(N__16397),
            .I(N__16389));
    InMux I__3402 (
            .O(N__16396),
            .I(N__16386));
    InMux I__3401 (
            .O(N__16395),
            .I(N__16383));
    LocalMux I__3400 (
            .O(N__16392),
            .I(N__16378));
    LocalMux I__3399 (
            .O(N__16389),
            .I(N__16378));
    LocalMux I__3398 (
            .O(N__16386),
            .I(\POWERLED.N_88 ));
    LocalMux I__3397 (
            .O(N__16383),
            .I(\POWERLED.N_88 ));
    Odrv4 I__3396 (
            .O(N__16378),
            .I(\POWERLED.N_88 ));
    CascadeMux I__3395 (
            .O(N__16371),
            .I(\POWERLED.N_205_cascade_ ));
    InMux I__3394 (
            .O(N__16368),
            .I(N__16362));
    InMux I__3393 (
            .O(N__16367),
            .I(N__16362));
    LocalMux I__3392 (
            .O(N__16362),
            .I(\POWERLED.N_203_4 ));
    CascadeMux I__3391 (
            .O(N__16359),
            .I(\POWERLED.count_clk_0_sqmuxa_5_0_a6_3_cascade_ ));
    InMux I__3390 (
            .O(N__16356),
            .I(N__16351));
    InMux I__3389 (
            .O(N__16355),
            .I(N__16346));
    InMux I__3388 (
            .O(N__16354),
            .I(N__16346));
    LocalMux I__3387 (
            .O(N__16351),
            .I(N__16338));
    LocalMux I__3386 (
            .O(N__16346),
            .I(N__16338));
    InMux I__3385 (
            .O(N__16345),
            .I(N__16333));
    InMux I__3384 (
            .O(N__16344),
            .I(N__16333));
    InMux I__3383 (
            .O(N__16343),
            .I(N__16330));
    Odrv4 I__3382 (
            .O(N__16338),
            .I(\POWERLED.N_226 ));
    LocalMux I__3381 (
            .O(N__16333),
            .I(\POWERLED.N_226 ));
    LocalMux I__3380 (
            .O(N__16330),
            .I(\POWERLED.N_226 ));
    InMux I__3379 (
            .O(N__16323),
            .I(N__16319));
    InMux I__3378 (
            .O(N__16322),
            .I(N__16316));
    LocalMux I__3377 (
            .O(N__16319),
            .I(N__16311));
    LocalMux I__3376 (
            .O(N__16316),
            .I(N__16311));
    Span4Mux_v I__3375 (
            .O(N__16311),
            .I(N__16308));
    Odrv4 I__3374 (
            .O(N__16308),
            .I(\POWERLED.N_200_2 ));
    InMux I__3373 (
            .O(N__16305),
            .I(N__16302));
    LocalMux I__3372 (
            .O(N__16302),
            .I(\POWERLED.N_217 ));
    CascadeMux I__3371 (
            .O(N__16299),
            .I(N__16294));
    InMux I__3370 (
            .O(N__16298),
            .I(N__16289));
    InMux I__3369 (
            .O(N__16297),
            .I(N__16289));
    InMux I__3368 (
            .O(N__16294),
            .I(N__16280));
    LocalMux I__3367 (
            .O(N__16289),
            .I(N__16277));
    InMux I__3366 (
            .O(N__16288),
            .I(N__16270));
    InMux I__3365 (
            .O(N__16287),
            .I(N__16270));
    InMux I__3364 (
            .O(N__16286),
            .I(N__16270));
    InMux I__3363 (
            .O(N__16285),
            .I(N__16267));
    InMux I__3362 (
            .O(N__16284),
            .I(N__16264));
    InMux I__3361 (
            .O(N__16283),
            .I(N__16261));
    LocalMux I__3360 (
            .O(N__16280),
            .I(N__16254));
    Span4Mux_v I__3359 (
            .O(N__16277),
            .I(N__16254));
    LocalMux I__3358 (
            .O(N__16270),
            .I(N__16254));
    LocalMux I__3357 (
            .O(N__16267),
            .I(\POWERLED.func_stateZ0Z_1 ));
    LocalMux I__3356 (
            .O(N__16264),
            .I(\POWERLED.func_stateZ0Z_1 ));
    LocalMux I__3355 (
            .O(N__16261),
            .I(\POWERLED.func_stateZ0Z_1 ));
    Odrv4 I__3354 (
            .O(N__16254),
            .I(\POWERLED.func_stateZ0Z_1 ));
    InMux I__3353 (
            .O(N__16245),
            .I(N__16242));
    LocalMux I__3352 (
            .O(N__16242),
            .I(\POWERLED.N_141 ));
    InMux I__3351 (
            .O(N__16239),
            .I(N__16236));
    LocalMux I__3350 (
            .O(N__16236),
            .I(\POWERLED.N_149 ));
    InMux I__3349 (
            .O(N__16233),
            .I(N__16224));
    InMux I__3348 (
            .O(N__16232),
            .I(N__16219));
    InMux I__3347 (
            .O(N__16231),
            .I(N__16219));
    InMux I__3346 (
            .O(N__16230),
            .I(N__16210));
    InMux I__3345 (
            .O(N__16229),
            .I(N__16210));
    InMux I__3344 (
            .O(N__16228),
            .I(N__16210));
    InMux I__3343 (
            .O(N__16227),
            .I(N__16210));
    LocalMux I__3342 (
            .O(N__16224),
            .I(N__16207));
    LocalMux I__3341 (
            .O(N__16219),
            .I(N__16202));
    LocalMux I__3340 (
            .O(N__16210),
            .I(N__16202));
    Span4Mux_s3_h I__3339 (
            .O(N__16207),
            .I(N__16197));
    Span4Mux_v I__3338 (
            .O(N__16202),
            .I(N__16197));
    Odrv4 I__3337 (
            .O(N__16197),
            .I(\POWERLED.N_222 ));
    CascadeMux I__3336 (
            .O(N__16194),
            .I(\POWERLED.N_149_cascade_ ));
    InMux I__3335 (
            .O(N__16191),
            .I(N__16184));
    InMux I__3334 (
            .O(N__16190),
            .I(N__16184));
    CascadeMux I__3333 (
            .O(N__16189),
            .I(N__16181));
    LocalMux I__3332 (
            .O(N__16184),
            .I(N__16178));
    InMux I__3331 (
            .O(N__16181),
            .I(N__16175));
    Span12Mux_s10_v I__3330 (
            .O(N__16178),
            .I(N__16170));
    LocalMux I__3329 (
            .O(N__16175),
            .I(N__16170));
    Odrv12 I__3328 (
            .O(N__16170),
            .I(\POWERLED.N_228 ));
    CascadeMux I__3327 (
            .O(N__16167),
            .I(N__16164));
    InMux I__3326 (
            .O(N__16164),
            .I(N__16161));
    LocalMux I__3325 (
            .O(N__16161),
            .I(\POWERLED.func_state_ns_i_0_0_1 ));
    InMux I__3324 (
            .O(N__16158),
            .I(N__16155));
    LocalMux I__3323 (
            .O(N__16155),
            .I(N__16150));
    InMux I__3322 (
            .O(N__16154),
            .I(N__16147));
    InMux I__3321 (
            .O(N__16153),
            .I(N__16144));
    Span4Mux_v I__3320 (
            .O(N__16150),
            .I(N__16141));
    LocalMux I__3319 (
            .O(N__16147),
            .I(N__16138));
    LocalMux I__3318 (
            .O(N__16144),
            .I(\POWERLED.N_248 ));
    Odrv4 I__3317 (
            .O(N__16141),
            .I(\POWERLED.N_248 ));
    Odrv4 I__3316 (
            .O(N__16138),
            .I(\POWERLED.N_248 ));
    InMux I__3315 (
            .O(N__16131),
            .I(N__16128));
    LocalMux I__3314 (
            .O(N__16128),
            .I(N__16125));
    Span4Mux_s3_h I__3313 (
            .O(N__16125),
            .I(N__16119));
    InMux I__3312 (
            .O(N__16124),
            .I(N__16116));
    InMux I__3311 (
            .O(N__16123),
            .I(N__16113));
    InMux I__3310 (
            .O(N__16122),
            .I(N__16110));
    Odrv4 I__3309 (
            .O(N__16119),
            .I(\POWERLED.N_127 ));
    LocalMux I__3308 (
            .O(N__16116),
            .I(\POWERLED.N_127 ));
    LocalMux I__3307 (
            .O(N__16113),
            .I(\POWERLED.N_127 ));
    LocalMux I__3306 (
            .O(N__16110),
            .I(\POWERLED.N_127 ));
    InMux I__3305 (
            .O(N__16101),
            .I(N__16098));
    LocalMux I__3304 (
            .O(N__16098),
            .I(N__16095));
    Odrv4 I__3303 (
            .O(N__16095),
            .I(\POWERLED.N_179 ));
    InMux I__3302 (
            .O(N__16092),
            .I(N__16089));
    LocalMux I__3301 (
            .O(N__16089),
            .I(\POWERLED.N_211 ));
    CascadeMux I__3300 (
            .O(N__16086),
            .I(N__16080));
    CascadeMux I__3299 (
            .O(N__16085),
            .I(N__16077));
    InMux I__3298 (
            .O(N__16084),
            .I(N__16074));
    CascadeMux I__3297 (
            .O(N__16083),
            .I(N__16071));
    InMux I__3296 (
            .O(N__16080),
            .I(N__16067));
    InMux I__3295 (
            .O(N__16077),
            .I(N__16064));
    LocalMux I__3294 (
            .O(N__16074),
            .I(N__16058));
    InMux I__3293 (
            .O(N__16071),
            .I(N__16051));
    InMux I__3292 (
            .O(N__16070),
            .I(N__16051));
    LocalMux I__3291 (
            .O(N__16067),
            .I(N__16048));
    LocalMux I__3290 (
            .O(N__16064),
            .I(N__16045));
    InMux I__3289 (
            .O(N__16063),
            .I(N__16038));
    InMux I__3288 (
            .O(N__16062),
            .I(N__16038));
    InMux I__3287 (
            .O(N__16061),
            .I(N__16038));
    Span4Mux_v I__3286 (
            .O(N__16058),
            .I(N__16035));
    InMux I__3285 (
            .O(N__16057),
            .I(N__16030));
    InMux I__3284 (
            .O(N__16056),
            .I(N__16030));
    LocalMux I__3283 (
            .O(N__16051),
            .I(N__16025));
    Span4Mux_h I__3282 (
            .O(N__16048),
            .I(N__16025));
    Odrv12 I__3281 (
            .O(N__16045),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__3280 (
            .O(N__16038),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv4 I__3279 (
            .O(N__16035),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__3278 (
            .O(N__16030),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv4 I__3277 (
            .O(N__16025),
            .I(\POWERLED.func_stateZ0Z_0 ));
    CascadeMux I__3276 (
            .O(N__16014),
            .I(\POWERLED.N_88_cascade_ ));
    CascadeMux I__3275 (
            .O(N__16011),
            .I(\POWERLED.dutycycle_3_sqmuxa_1_i_0_1_1_cascade_ ));
    InMux I__3274 (
            .O(N__16008),
            .I(N__16004));
    InMux I__3273 (
            .O(N__16007),
            .I(N__16001));
    LocalMux I__3272 (
            .O(N__16004),
            .I(N__15996));
    LocalMux I__3271 (
            .O(N__16001),
            .I(N__15996));
    Span4Mux_h I__3270 (
            .O(N__15996),
            .I(N__15993));
    Odrv4 I__3269 (
            .O(N__15993),
            .I(\POWERLED.N_366_1 ));
    InMux I__3268 (
            .O(N__15990),
            .I(N__15987));
    LocalMux I__3267 (
            .O(N__15987),
            .I(\POWERLED.count_clk_1_sqmuxa_5_0_2 ));
    InMux I__3266 (
            .O(N__15984),
            .I(N__15980));
    InMux I__3265 (
            .O(N__15983),
            .I(N__15977));
    LocalMux I__3264 (
            .O(N__15980),
            .I(\COUNTER.counterZ0Z_26 ));
    LocalMux I__3263 (
            .O(N__15977),
            .I(\COUNTER.counterZ0Z_26 ));
    InMux I__3262 (
            .O(N__15972),
            .I(N__15968));
    InMux I__3261 (
            .O(N__15971),
            .I(N__15965));
    LocalMux I__3260 (
            .O(N__15968),
            .I(\COUNTER.counterZ0Z_25 ));
    LocalMux I__3259 (
            .O(N__15965),
            .I(\COUNTER.counterZ0Z_25 ));
    CascadeMux I__3258 (
            .O(N__15960),
            .I(N__15956));
    InMux I__3257 (
            .O(N__15959),
            .I(N__15953));
    InMux I__3256 (
            .O(N__15956),
            .I(N__15950));
    LocalMux I__3255 (
            .O(N__15953),
            .I(\COUNTER.counterZ0Z_27 ));
    LocalMux I__3254 (
            .O(N__15950),
            .I(\COUNTER.counterZ0Z_27 ));
    InMux I__3253 (
            .O(N__15945),
            .I(N__15941));
    InMux I__3252 (
            .O(N__15944),
            .I(N__15938));
    LocalMux I__3251 (
            .O(N__15941),
            .I(\COUNTER.counterZ0Z_24 ));
    LocalMux I__3250 (
            .O(N__15938),
            .I(\COUNTER.counterZ0Z_24 ));
    InMux I__3249 (
            .O(N__15933),
            .I(N__15930));
    LocalMux I__3248 (
            .O(N__15930),
            .I(N__15927));
    Odrv4 I__3247 (
            .O(N__15927),
            .I(\COUNTER.un4_counter_6_and ));
    InMux I__3246 (
            .O(N__15924),
            .I(N__15920));
    InMux I__3245 (
            .O(N__15923),
            .I(N__15917));
    LocalMux I__3244 (
            .O(N__15920),
            .I(\COUNTER.counterZ0Z_22 ));
    LocalMux I__3243 (
            .O(N__15917),
            .I(\COUNTER.counterZ0Z_22 ));
    InMux I__3242 (
            .O(N__15912),
            .I(N__15908));
    InMux I__3241 (
            .O(N__15911),
            .I(N__15905));
    LocalMux I__3240 (
            .O(N__15908),
            .I(\COUNTER.counterZ0Z_21 ));
    LocalMux I__3239 (
            .O(N__15905),
            .I(\COUNTER.counterZ0Z_21 ));
    CascadeMux I__3238 (
            .O(N__15900),
            .I(N__15896));
    InMux I__3237 (
            .O(N__15899),
            .I(N__15893));
    InMux I__3236 (
            .O(N__15896),
            .I(N__15890));
    LocalMux I__3235 (
            .O(N__15893),
            .I(\COUNTER.counterZ0Z_23 ));
    LocalMux I__3234 (
            .O(N__15890),
            .I(\COUNTER.counterZ0Z_23 ));
    InMux I__3233 (
            .O(N__15885),
            .I(N__15881));
    InMux I__3232 (
            .O(N__15884),
            .I(N__15878));
    LocalMux I__3231 (
            .O(N__15881),
            .I(\COUNTER.counterZ0Z_20 ));
    LocalMux I__3230 (
            .O(N__15878),
            .I(\COUNTER.counterZ0Z_20 ));
    InMux I__3229 (
            .O(N__15873),
            .I(N__15870));
    LocalMux I__3228 (
            .O(N__15870),
            .I(N__15867));
    Odrv12 I__3227 (
            .O(N__15867),
            .I(\COUNTER.un4_counter_5_and ));
    CascadeMux I__3226 (
            .O(N__15864),
            .I(N__15857));
    InMux I__3225 (
            .O(N__15863),
            .I(N__15853));
    InMux I__3224 (
            .O(N__15862),
            .I(N__15850));
    InMux I__3223 (
            .O(N__15861),
            .I(N__15845));
    InMux I__3222 (
            .O(N__15860),
            .I(N__15845));
    InMux I__3221 (
            .O(N__15857),
            .I(N__15842));
    InMux I__3220 (
            .O(N__15856),
            .I(N__15839));
    LocalMux I__3219 (
            .O(N__15853),
            .I(N__15836));
    LocalMux I__3218 (
            .O(N__15850),
            .I(\POWERLED.N_214 ));
    LocalMux I__3217 (
            .O(N__15845),
            .I(\POWERLED.N_214 ));
    LocalMux I__3216 (
            .O(N__15842),
            .I(\POWERLED.N_214 ));
    LocalMux I__3215 (
            .O(N__15839),
            .I(\POWERLED.N_214 ));
    Odrv4 I__3214 (
            .O(N__15836),
            .I(\POWERLED.N_214 ));
    InMux I__3213 (
            .O(N__15825),
            .I(N__15821));
    InMux I__3212 (
            .O(N__15824),
            .I(N__15818));
    LocalMux I__3211 (
            .O(N__15821),
            .I(N__15815));
    LocalMux I__3210 (
            .O(N__15818),
            .I(\POWERLED.N_250 ));
    Odrv4 I__3209 (
            .O(N__15815),
            .I(\POWERLED.N_250 ));
    InMux I__3208 (
            .O(N__15810),
            .I(N__15807));
    LocalMux I__3207 (
            .O(N__15807),
            .I(\POWERLED.N_178 ));
    CascadeMux I__3206 (
            .O(N__15804),
            .I(\POWERLED.N_148_cascade_ ));
    CascadeMux I__3205 (
            .O(N__15801),
            .I(\POWERLED.N_208_cascade_ ));
    InMux I__3204 (
            .O(N__15798),
            .I(N__15795));
    LocalMux I__3203 (
            .O(N__15795),
            .I(\POWERLED.func_state_ns_i_0_1_1 ));
    InMux I__3202 (
            .O(N__15792),
            .I(N__15789));
    LocalMux I__3201 (
            .O(N__15789),
            .I(\COUNTER.counter_1_cry_5_THRU_CO ));
    InMux I__3200 (
            .O(N__15786),
            .I(N__15783));
    LocalMux I__3199 (
            .O(N__15783),
            .I(\COUNTER.counter_1_cry_4_THRU_CO ));
    InMux I__3198 (
            .O(N__15780),
            .I(N__15768));
    InMux I__3197 (
            .O(N__15779),
            .I(N__15768));
    InMux I__3196 (
            .O(N__15778),
            .I(N__15761));
    InMux I__3195 (
            .O(N__15777),
            .I(N__15761));
    InMux I__3194 (
            .O(N__15776),
            .I(N__15761));
    InMux I__3193 (
            .O(N__15775),
            .I(N__15754));
    InMux I__3192 (
            .O(N__15774),
            .I(N__15754));
    InMux I__3191 (
            .O(N__15773),
            .I(N__15754));
    LocalMux I__3190 (
            .O(N__15768),
            .I(N__15751));
    LocalMux I__3189 (
            .O(N__15761),
            .I(\COUNTER.un4_counter_7_THRU_CO ));
    LocalMux I__3188 (
            .O(N__15754),
            .I(\COUNTER.un4_counter_7_THRU_CO ));
    Odrv12 I__3187 (
            .O(N__15751),
            .I(\COUNTER.un4_counter_7_THRU_CO ));
    CascadeMux I__3186 (
            .O(N__15744),
            .I(N__15739));
    InMux I__3185 (
            .O(N__15743),
            .I(N__15733));
    InMux I__3184 (
            .O(N__15742),
            .I(N__15733));
    InMux I__3183 (
            .O(N__15739),
            .I(N__15730));
    InMux I__3182 (
            .O(N__15738),
            .I(N__15727));
    LocalMux I__3181 (
            .O(N__15733),
            .I(\COUNTER.counterZ0Z_0 ));
    LocalMux I__3180 (
            .O(N__15730),
            .I(\COUNTER.counterZ0Z_0 ));
    LocalMux I__3179 (
            .O(N__15727),
            .I(\COUNTER.counterZ0Z_0 ));
    InMux I__3178 (
            .O(N__15720),
            .I(N__15715));
    InMux I__3177 (
            .O(N__15719),
            .I(N__15710));
    InMux I__3176 (
            .O(N__15718),
            .I(N__15710));
    LocalMux I__3175 (
            .O(N__15715),
            .I(\COUNTER.counterZ0Z_6 ));
    LocalMux I__3174 (
            .O(N__15710),
            .I(\COUNTER.counterZ0Z_6 ));
    InMux I__3173 (
            .O(N__15705),
            .I(N__15700));
    InMux I__3172 (
            .O(N__15704),
            .I(N__15695));
    InMux I__3171 (
            .O(N__15703),
            .I(N__15695));
    LocalMux I__3170 (
            .O(N__15700),
            .I(\COUNTER.counterZ0Z_5 ));
    LocalMux I__3169 (
            .O(N__15695),
            .I(\COUNTER.counterZ0Z_5 ));
    CascadeMux I__3168 (
            .O(N__15690),
            .I(N__15686));
    InMux I__3167 (
            .O(N__15689),
            .I(N__15683));
    InMux I__3166 (
            .O(N__15686),
            .I(N__15680));
    LocalMux I__3165 (
            .O(N__15683),
            .I(\COUNTER.counterZ0Z_7 ));
    LocalMux I__3164 (
            .O(N__15680),
            .I(\COUNTER.counterZ0Z_7 ));
    InMux I__3163 (
            .O(N__15675),
            .I(N__15670));
    InMux I__3162 (
            .O(N__15674),
            .I(N__15665));
    InMux I__3161 (
            .O(N__15673),
            .I(N__15665));
    LocalMux I__3160 (
            .O(N__15670),
            .I(\COUNTER.counterZ0Z_1 ));
    LocalMux I__3159 (
            .O(N__15665),
            .I(\COUNTER.counterZ0Z_1 ));
    InMux I__3158 (
            .O(N__15660),
            .I(N__15657));
    LocalMux I__3157 (
            .O(N__15657),
            .I(\COUNTER.un4_counter_1_and ));
    InMux I__3156 (
            .O(N__15654),
            .I(N__15650));
    InMux I__3155 (
            .O(N__15653),
            .I(N__15647));
    LocalMux I__3154 (
            .O(N__15650),
            .I(\COUNTER.counterZ0Z_18 ));
    LocalMux I__3153 (
            .O(N__15647),
            .I(\COUNTER.counterZ0Z_18 ));
    InMux I__3152 (
            .O(N__15642),
            .I(N__15638));
    InMux I__3151 (
            .O(N__15641),
            .I(N__15635));
    LocalMux I__3150 (
            .O(N__15638),
            .I(\COUNTER.counterZ0Z_17 ));
    LocalMux I__3149 (
            .O(N__15635),
            .I(\COUNTER.counterZ0Z_17 ));
    CascadeMux I__3148 (
            .O(N__15630),
            .I(N__15626));
    InMux I__3147 (
            .O(N__15629),
            .I(N__15623));
    InMux I__3146 (
            .O(N__15626),
            .I(N__15620));
    LocalMux I__3145 (
            .O(N__15623),
            .I(\COUNTER.counterZ0Z_19 ));
    LocalMux I__3144 (
            .O(N__15620),
            .I(\COUNTER.counterZ0Z_19 ));
    InMux I__3143 (
            .O(N__15615),
            .I(N__15611));
    InMux I__3142 (
            .O(N__15614),
            .I(N__15608));
    LocalMux I__3141 (
            .O(N__15611),
            .I(\COUNTER.counterZ0Z_16 ));
    LocalMux I__3140 (
            .O(N__15608),
            .I(\COUNTER.counterZ0Z_16 ));
    InMux I__3139 (
            .O(N__15603),
            .I(N__15600));
    LocalMux I__3138 (
            .O(N__15600),
            .I(N__15597));
    Odrv4 I__3137 (
            .O(N__15597),
            .I(\COUNTER.un4_counter_4_and ));
    InMux I__3136 (
            .O(N__15594),
            .I(N__15590));
    InMux I__3135 (
            .O(N__15593),
            .I(N__15587));
    LocalMux I__3134 (
            .O(N__15590),
            .I(\COUNTER.counterZ0Z_10 ));
    LocalMux I__3133 (
            .O(N__15587),
            .I(\COUNTER.counterZ0Z_10 ));
    InMux I__3132 (
            .O(N__15582),
            .I(N__15578));
    InMux I__3131 (
            .O(N__15581),
            .I(N__15575));
    LocalMux I__3130 (
            .O(N__15578),
            .I(\COUNTER.counterZ0Z_9 ));
    LocalMux I__3129 (
            .O(N__15575),
            .I(\COUNTER.counterZ0Z_9 ));
    CascadeMux I__3128 (
            .O(N__15570),
            .I(N__15566));
    InMux I__3127 (
            .O(N__15569),
            .I(N__15563));
    InMux I__3126 (
            .O(N__15566),
            .I(N__15560));
    LocalMux I__3125 (
            .O(N__15563),
            .I(\COUNTER.counterZ0Z_11 ));
    LocalMux I__3124 (
            .O(N__15560),
            .I(\COUNTER.counterZ0Z_11 ));
    InMux I__3123 (
            .O(N__15555),
            .I(N__15551));
    InMux I__3122 (
            .O(N__15554),
            .I(N__15548));
    LocalMux I__3121 (
            .O(N__15551),
            .I(\COUNTER.counterZ0Z_8 ));
    LocalMux I__3120 (
            .O(N__15548),
            .I(\COUNTER.counterZ0Z_8 ));
    InMux I__3119 (
            .O(N__15543),
            .I(N__15540));
    LocalMux I__3118 (
            .O(N__15540),
            .I(N__15537));
    Odrv4 I__3117 (
            .O(N__15537),
            .I(\COUNTER.un4_counter_2_and ));
    InMux I__3116 (
            .O(N__15534),
            .I(N__15530));
    InMux I__3115 (
            .O(N__15533),
            .I(N__15527));
    LocalMux I__3114 (
            .O(N__15530),
            .I(\COUNTER.counterZ0Z_14 ));
    LocalMux I__3113 (
            .O(N__15527),
            .I(\COUNTER.counterZ0Z_14 ));
    InMux I__3112 (
            .O(N__15522),
            .I(N__15518));
    InMux I__3111 (
            .O(N__15521),
            .I(N__15515));
    LocalMux I__3110 (
            .O(N__15518),
            .I(\COUNTER.counterZ0Z_13 ));
    LocalMux I__3109 (
            .O(N__15515),
            .I(\COUNTER.counterZ0Z_13 ));
    CascadeMux I__3108 (
            .O(N__15510),
            .I(N__15506));
    InMux I__3107 (
            .O(N__15509),
            .I(N__15503));
    InMux I__3106 (
            .O(N__15506),
            .I(N__15500));
    LocalMux I__3105 (
            .O(N__15503),
            .I(\COUNTER.counterZ0Z_15 ));
    LocalMux I__3104 (
            .O(N__15500),
            .I(\COUNTER.counterZ0Z_15 ));
    InMux I__3103 (
            .O(N__15495),
            .I(N__15491));
    InMux I__3102 (
            .O(N__15494),
            .I(N__15488));
    LocalMux I__3101 (
            .O(N__15491),
            .I(\COUNTER.counterZ0Z_12 ));
    LocalMux I__3100 (
            .O(N__15488),
            .I(\COUNTER.counterZ0Z_12 ));
    InMux I__3099 (
            .O(N__15483),
            .I(N__15480));
    LocalMux I__3098 (
            .O(N__15480),
            .I(N__15477));
    Odrv4 I__3097 (
            .O(N__15477),
            .I(\COUNTER.un4_counter_3_and ));
    InMux I__3096 (
            .O(N__15474),
            .I(N__15471));
    LocalMux I__3095 (
            .O(N__15471),
            .I(N__15468));
    Span4Mux_v I__3094 (
            .O(N__15468),
            .I(N__15465));
    Odrv4 I__3093 (
            .O(N__15465),
            .I(\COUNTER.un4_counter_7_and ));
    InMux I__3092 (
            .O(N__15462),
            .I(bfn_9_5_0_));
    CascadeMux I__3091 (
            .O(N__15459),
            .I(\COUNTER.un4_counter_7_THRU_CO_cascade_ ));
    InMux I__3090 (
            .O(N__15456),
            .I(bfn_8_15_0_));
    InMux I__3089 (
            .O(N__15453),
            .I(N__15449));
    InMux I__3088 (
            .O(N__15452),
            .I(N__15446));
    LocalMux I__3087 (
            .O(N__15449),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    LocalMux I__3086 (
            .O(N__15446),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    InMux I__3085 (
            .O(N__15441),
            .I(N__15437));
    InMux I__3084 (
            .O(N__15440),
            .I(N__15434));
    LocalMux I__3083 (
            .O(N__15437),
            .I(\PCH_PWRGD.countZ0Z_1 ));
    LocalMux I__3082 (
            .O(N__15434),
            .I(\PCH_PWRGD.countZ0Z_1 ));
    CascadeMux I__3081 (
            .O(N__15429),
            .I(N__15425));
    InMux I__3080 (
            .O(N__15428),
            .I(N__15422));
    InMux I__3079 (
            .O(N__15425),
            .I(N__15419));
    LocalMux I__3078 (
            .O(N__15422),
            .I(\PCH_PWRGD.countZ0Z_10 ));
    LocalMux I__3077 (
            .O(N__15419),
            .I(\PCH_PWRGD.countZ0Z_10 ));
    InMux I__3076 (
            .O(N__15414),
            .I(N__15410));
    InMux I__3075 (
            .O(N__15413),
            .I(N__15407));
    LocalMux I__3074 (
            .O(N__15410),
            .I(\PCH_PWRGD.countZ0Z_2 ));
    LocalMux I__3073 (
            .O(N__15407),
            .I(\PCH_PWRGD.countZ0Z_2 ));
    CascadeMux I__3072 (
            .O(N__15402),
            .I(\PCH_PWRGD.un4_count_9_cascade_ ));
    CascadeMux I__3071 (
            .O(N__15399),
            .I(N__15395));
    CascadeMux I__3070 (
            .O(N__15398),
            .I(N__15392));
    InMux I__3069 (
            .O(N__15395),
            .I(N__15389));
    InMux I__3068 (
            .O(N__15392),
            .I(N__15386));
    LocalMux I__3067 (
            .O(N__15389),
            .I(N__15380));
    LocalMux I__3066 (
            .O(N__15386),
            .I(N__15380));
    InMux I__3065 (
            .O(N__15385),
            .I(N__15377));
    Span4Mux_v I__3064 (
            .O(N__15380),
            .I(N__15372));
    LocalMux I__3063 (
            .O(N__15377),
            .I(N__15372));
    Odrv4 I__3062 (
            .O(N__15372),
            .I(\PCH_PWRGD.N_1_i ));
    InMux I__3061 (
            .O(N__15369),
            .I(N__15365));
    InMux I__3060 (
            .O(N__15368),
            .I(N__15362));
    LocalMux I__3059 (
            .O(N__15365),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    LocalMux I__3058 (
            .O(N__15362),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    InMux I__3057 (
            .O(N__15357),
            .I(N__15353));
    InMux I__3056 (
            .O(N__15356),
            .I(N__15350));
    LocalMux I__3055 (
            .O(N__15353),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    LocalMux I__3054 (
            .O(N__15350),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    CascadeMux I__3053 (
            .O(N__15345),
            .I(N__15341));
    InMux I__3052 (
            .O(N__15344),
            .I(N__15338));
    InMux I__3051 (
            .O(N__15341),
            .I(N__15335));
    LocalMux I__3050 (
            .O(N__15338),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    LocalMux I__3049 (
            .O(N__15335),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    InMux I__3048 (
            .O(N__15330),
            .I(N__15326));
    InMux I__3047 (
            .O(N__15329),
            .I(N__15323));
    LocalMux I__3046 (
            .O(N__15326),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    LocalMux I__3045 (
            .O(N__15323),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    InMux I__3044 (
            .O(N__15318),
            .I(N__15315));
    LocalMux I__3043 (
            .O(N__15315),
            .I(\PCH_PWRGD.un4_count_11 ));
    InMux I__3042 (
            .O(N__15312),
            .I(N__15308));
    InMux I__3041 (
            .O(N__15311),
            .I(N__15305));
    LocalMux I__3040 (
            .O(N__15308),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    LocalMux I__3039 (
            .O(N__15305),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    InMux I__3038 (
            .O(N__15300),
            .I(N__15296));
    InMux I__3037 (
            .O(N__15299),
            .I(N__15293));
    LocalMux I__3036 (
            .O(N__15296),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    LocalMux I__3035 (
            .O(N__15293),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    CascadeMux I__3034 (
            .O(N__15288),
            .I(N__15284));
    InMux I__3033 (
            .O(N__15287),
            .I(N__15281));
    InMux I__3032 (
            .O(N__15284),
            .I(N__15278));
    LocalMux I__3031 (
            .O(N__15281),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    LocalMux I__3030 (
            .O(N__15278),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    InMux I__3029 (
            .O(N__15273),
            .I(N__15269));
    InMux I__3028 (
            .O(N__15272),
            .I(N__15266));
    LocalMux I__3027 (
            .O(N__15269),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    LocalMux I__3026 (
            .O(N__15266),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    InMux I__3025 (
            .O(N__15261),
            .I(N__15258));
    LocalMux I__3024 (
            .O(N__15258),
            .I(\PCH_PWRGD.un4_count_10 ));
    InMux I__3023 (
            .O(N__15255),
            .I(N__15251));
    InMux I__3022 (
            .O(N__15254),
            .I(N__15248));
    LocalMux I__3021 (
            .O(N__15251),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    LocalMux I__3020 (
            .O(N__15248),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    InMux I__3019 (
            .O(N__15243),
            .I(N__15239));
    InMux I__3018 (
            .O(N__15242),
            .I(N__15236));
    LocalMux I__3017 (
            .O(N__15239),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    LocalMux I__3016 (
            .O(N__15236),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    CascadeMux I__3015 (
            .O(N__15231),
            .I(N__15227));
    InMux I__3014 (
            .O(N__15230),
            .I(N__15224));
    InMux I__3013 (
            .O(N__15227),
            .I(N__15221));
    LocalMux I__3012 (
            .O(N__15224),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    LocalMux I__3011 (
            .O(N__15221),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    InMux I__3010 (
            .O(N__15216),
            .I(N__15212));
    InMux I__3009 (
            .O(N__15215),
            .I(N__15209));
    LocalMux I__3008 (
            .O(N__15212),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    LocalMux I__3007 (
            .O(N__15209),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    InMux I__3006 (
            .O(N__15204),
            .I(N__15201));
    LocalMux I__3005 (
            .O(N__15201),
            .I(\PCH_PWRGD.un4_count_8 ));
    InMux I__3004 (
            .O(N__15198),
            .I(N__15195));
    LocalMux I__3003 (
            .O(N__15195),
            .I(\COUNTER.un4_counter_0_and ));
    InMux I__3002 (
            .O(N__15192),
            .I(N__15186));
    InMux I__3001 (
            .O(N__15191),
            .I(N__15179));
    InMux I__3000 (
            .O(N__15190),
            .I(N__15179));
    InMux I__2999 (
            .O(N__15189),
            .I(N__15179));
    LocalMux I__2998 (
            .O(N__15186),
            .I(\POWERLED.count_clkZ0Z_6 ));
    LocalMux I__2997 (
            .O(N__15179),
            .I(\POWERLED.count_clkZ0Z_6 ));
    InMux I__2996 (
            .O(N__15174),
            .I(\POWERLED.un1_count_clk_1_cry_5 ));
    InMux I__2995 (
            .O(N__15171),
            .I(\POWERLED.un1_count_clk_1_cry_6 ));
    CascadeMux I__2994 (
            .O(N__15168),
            .I(N__15165));
    InMux I__2993 (
            .O(N__15165),
            .I(N__15158));
    InMux I__2992 (
            .O(N__15164),
            .I(N__15158));
    InMux I__2991 (
            .O(N__15163),
            .I(N__15155));
    LocalMux I__2990 (
            .O(N__15158),
            .I(N__15152));
    LocalMux I__2989 (
            .O(N__15155),
            .I(\POWERLED.count_clkZ0Z_8 ));
    Odrv4 I__2988 (
            .O(N__15152),
            .I(\POWERLED.count_clkZ0Z_8 ));
    InMux I__2987 (
            .O(N__15147),
            .I(bfn_8_14_0_));
    InMux I__2986 (
            .O(N__15144),
            .I(\POWERLED.un1_count_clk_1_cry_8 ));
    InMux I__2985 (
            .O(N__15141),
            .I(\POWERLED.un1_count_clk_1_cry_9 ));
    InMux I__2984 (
            .O(N__15138),
            .I(\POWERLED.un1_count_clk_1_cry_10 ));
    InMux I__2983 (
            .O(N__15135),
            .I(\POWERLED.un1_count_clk_1_cry_11 ));
    InMux I__2982 (
            .O(N__15132),
            .I(\POWERLED.un1_count_clk_1_cry_12 ));
    InMux I__2981 (
            .O(N__15129),
            .I(\POWERLED.un1_count_clk_1_cry_13 ));
    CascadeMux I__2980 (
            .O(N__15126),
            .I(\POWERLED.count_clk_0_sqmuxa_5_0_o2_0_0_cascade_ ));
    CascadeMux I__2979 (
            .O(N__15123),
            .I(\POWERLED.N_141_cascade_ ));
    CascadeMux I__2978 (
            .O(N__15120),
            .I(N__15116));
    InMux I__2977 (
            .O(N__15119),
            .I(N__15113));
    InMux I__2976 (
            .O(N__15116),
            .I(N__15110));
    LocalMux I__2975 (
            .O(N__15113),
            .I(N__15105));
    LocalMux I__2974 (
            .O(N__15110),
            .I(N__15105));
    Odrv4 I__2973 (
            .O(N__15105),
            .I(\POWERLED.count_clk_1_sqmuxa_5_i ));
    InMux I__2972 (
            .O(N__15102),
            .I(\POWERLED.un1_count_clk_1_cry_0 ));
    InMux I__2971 (
            .O(N__15099),
            .I(N__15094));
    InMux I__2970 (
            .O(N__15098),
            .I(N__15089));
    InMux I__2969 (
            .O(N__15097),
            .I(N__15089));
    LocalMux I__2968 (
            .O(N__15094),
            .I(\POWERLED.count_clkZ0Z_2 ));
    LocalMux I__2967 (
            .O(N__15089),
            .I(\POWERLED.count_clkZ0Z_2 ));
    InMux I__2966 (
            .O(N__15084),
            .I(\POWERLED.un1_count_clk_1_cry_1 ));
    InMux I__2965 (
            .O(N__15081),
            .I(N__15076));
    InMux I__2964 (
            .O(N__15080),
            .I(N__15073));
    InMux I__2963 (
            .O(N__15079),
            .I(N__15070));
    LocalMux I__2962 (
            .O(N__15076),
            .I(\POWERLED.count_clkZ0Z_3 ));
    LocalMux I__2961 (
            .O(N__15073),
            .I(\POWERLED.count_clkZ0Z_3 ));
    LocalMux I__2960 (
            .O(N__15070),
            .I(\POWERLED.count_clkZ0Z_3 ));
    InMux I__2959 (
            .O(N__15063),
            .I(\POWERLED.un1_count_clk_1_cry_2 ));
    InMux I__2958 (
            .O(N__15060),
            .I(N__15055));
    InMux I__2957 (
            .O(N__15059),
            .I(N__15050));
    InMux I__2956 (
            .O(N__15058),
            .I(N__15050));
    LocalMux I__2955 (
            .O(N__15055),
            .I(\POWERLED.count_clkZ0Z_4 ));
    LocalMux I__2954 (
            .O(N__15050),
            .I(\POWERLED.count_clkZ0Z_4 ));
    InMux I__2953 (
            .O(N__15045),
            .I(\POWERLED.un1_count_clk_1_cry_3 ));
    InMux I__2952 (
            .O(N__15042),
            .I(\POWERLED.un1_count_clk_1_cry_4 ));
    CascadeMux I__2951 (
            .O(N__15039),
            .I(N__15030));
    CascadeMux I__2950 (
            .O(N__15038),
            .I(N__15025));
    InMux I__2949 (
            .O(N__15037),
            .I(N__15022));
    InMux I__2948 (
            .O(N__15036),
            .I(N__15019));
    InMux I__2947 (
            .O(N__15035),
            .I(N__15014));
    InMux I__2946 (
            .O(N__15034),
            .I(N__15014));
    InMux I__2945 (
            .O(N__15033),
            .I(N__15011));
    InMux I__2944 (
            .O(N__15030),
            .I(N__15002));
    InMux I__2943 (
            .O(N__15029),
            .I(N__15002));
    InMux I__2942 (
            .O(N__15028),
            .I(N__15002));
    InMux I__2941 (
            .O(N__15025),
            .I(N__15002));
    LocalMux I__2940 (
            .O(N__15022),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__2939 (
            .O(N__15019),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__2938 (
            .O(N__15014),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__2937 (
            .O(N__15011),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__2936 (
            .O(N__15002),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    CascadeMux I__2935 (
            .O(N__14991),
            .I(N__14987));
    CascadeMux I__2934 (
            .O(N__14990),
            .I(N__14977));
    InMux I__2933 (
            .O(N__14987),
            .I(N__14974));
    InMux I__2932 (
            .O(N__14986),
            .I(N__14971));
    InMux I__2931 (
            .O(N__14985),
            .I(N__14962));
    InMux I__2930 (
            .O(N__14984),
            .I(N__14962));
    InMux I__2929 (
            .O(N__14983),
            .I(N__14962));
    InMux I__2928 (
            .O(N__14982),
            .I(N__14962));
    InMux I__2927 (
            .O(N__14981),
            .I(N__14955));
    InMux I__2926 (
            .O(N__14980),
            .I(N__14955));
    InMux I__2925 (
            .O(N__14977),
            .I(N__14955));
    LocalMux I__2924 (
            .O(N__14974),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__2923 (
            .O(N__14971),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__2922 (
            .O(N__14962),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__2921 (
            .O(N__14955),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    CascadeMux I__2920 (
            .O(N__14946),
            .I(N__14939));
    CascadeMux I__2919 (
            .O(N__14945),
            .I(N__14936));
    CascadeMux I__2918 (
            .O(N__14944),
            .I(N__14931));
    InMux I__2917 (
            .O(N__14943),
            .I(N__14925));
    InMux I__2916 (
            .O(N__14942),
            .I(N__14925));
    InMux I__2915 (
            .O(N__14939),
            .I(N__14922));
    InMux I__2914 (
            .O(N__14936),
            .I(N__14917));
    InMux I__2913 (
            .O(N__14935),
            .I(N__14917));
    InMux I__2912 (
            .O(N__14934),
            .I(N__14910));
    InMux I__2911 (
            .O(N__14931),
            .I(N__14910));
    InMux I__2910 (
            .O(N__14930),
            .I(N__14910));
    LocalMux I__2909 (
            .O(N__14925),
            .I(N__14907));
    LocalMux I__2908 (
            .O(N__14922),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__2907 (
            .O(N__14917),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__2906 (
            .O(N__14910),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__2905 (
            .O(N__14907),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    InMux I__2904 (
            .O(N__14898),
            .I(N__14887));
    InMux I__2903 (
            .O(N__14897),
            .I(N__14887));
    InMux I__2902 (
            .O(N__14896),
            .I(N__14882));
    InMux I__2901 (
            .O(N__14895),
            .I(N__14877));
    InMux I__2900 (
            .O(N__14894),
            .I(N__14877));
    InMux I__2899 (
            .O(N__14893),
            .I(N__14872));
    InMux I__2898 (
            .O(N__14892),
            .I(N__14872));
    LocalMux I__2897 (
            .O(N__14887),
            .I(N__14869));
    InMux I__2896 (
            .O(N__14886),
            .I(N__14864));
    InMux I__2895 (
            .O(N__14885),
            .I(N__14864));
    LocalMux I__2894 (
            .O(N__14882),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__2893 (
            .O(N__14877),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__2892 (
            .O(N__14872),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__2891 (
            .O(N__14869),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__2890 (
            .O(N__14864),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    InMux I__2889 (
            .O(N__14853),
            .I(N__14850));
    LocalMux I__2888 (
            .O(N__14850),
            .I(\POWERLED.un2_slp_s3n_2_0_o2_3_7 ));
    CascadeMux I__2887 (
            .O(N__14847),
            .I(\POWERLED.un2_slp_s3n_2_0_o2_3_8_cascade_ ));
    InMux I__2886 (
            .O(N__14844),
            .I(N__14841));
    LocalMux I__2885 (
            .O(N__14841),
            .I(\POWERLED.un2_slp_s3n_2_0_o2_3_6 ));
    CascadeMux I__2884 (
            .O(N__14838),
            .I(N__14835));
    InMux I__2883 (
            .O(N__14835),
            .I(N__14830));
    InMux I__2882 (
            .O(N__14834),
            .I(N__14825));
    InMux I__2881 (
            .O(N__14833),
            .I(N__14825));
    LocalMux I__2880 (
            .O(N__14830),
            .I(N__14820));
    LocalMux I__2879 (
            .O(N__14825),
            .I(N__14820));
    Span4Mux_v I__2878 (
            .O(N__14820),
            .I(N__14817));
    Odrv4 I__2877 (
            .O(N__14817),
            .I(\POWERLED.N_112 ));
    CascadeMux I__2876 (
            .O(N__14814),
            .I(\POWERLED.N_177_5_cascade_ ));
    InMux I__2875 (
            .O(N__14811),
            .I(N__14808));
    LocalMux I__2874 (
            .O(N__14808),
            .I(\POWERLED.N_177_5 ));
    CascadeMux I__2873 (
            .O(N__14805),
            .I(\POWERLED.N_368_0_i_i_a6_0_cascade_ ));
    CascadeMux I__2872 (
            .O(N__14802),
            .I(N__14792));
    CascadeMux I__2871 (
            .O(N__14801),
            .I(N__14788));
    CascadeMux I__2870 (
            .O(N__14800),
            .I(N__14784));
    CascadeMux I__2869 (
            .O(N__14799),
            .I(N__14780));
    CascadeMux I__2868 (
            .O(N__14798),
            .I(N__14775));
    CascadeMux I__2867 (
            .O(N__14797),
            .I(N__14771));
    CascadeMux I__2866 (
            .O(N__14796),
            .I(N__14766));
    InMux I__2865 (
            .O(N__14795),
            .I(N__14763));
    InMux I__2864 (
            .O(N__14792),
            .I(N__14746));
    InMux I__2863 (
            .O(N__14791),
            .I(N__14746));
    InMux I__2862 (
            .O(N__14788),
            .I(N__14746));
    InMux I__2861 (
            .O(N__14787),
            .I(N__14746));
    InMux I__2860 (
            .O(N__14784),
            .I(N__14746));
    InMux I__2859 (
            .O(N__14783),
            .I(N__14746));
    InMux I__2858 (
            .O(N__14780),
            .I(N__14746));
    InMux I__2857 (
            .O(N__14779),
            .I(N__14746));
    InMux I__2856 (
            .O(N__14778),
            .I(N__14735));
    InMux I__2855 (
            .O(N__14775),
            .I(N__14735));
    InMux I__2854 (
            .O(N__14774),
            .I(N__14735));
    InMux I__2853 (
            .O(N__14771),
            .I(N__14735));
    InMux I__2852 (
            .O(N__14770),
            .I(N__14735));
    InMux I__2851 (
            .O(N__14769),
            .I(N__14730));
    InMux I__2850 (
            .O(N__14766),
            .I(N__14730));
    LocalMux I__2849 (
            .O(N__14763),
            .I(\POWERLED.N_177 ));
    LocalMux I__2848 (
            .O(N__14746),
            .I(\POWERLED.N_177 ));
    LocalMux I__2847 (
            .O(N__14735),
            .I(\POWERLED.N_177 ));
    LocalMux I__2846 (
            .O(N__14730),
            .I(\POWERLED.N_177 ));
    IoInMux I__2845 (
            .O(N__14721),
            .I(N__14718));
    LocalMux I__2844 (
            .O(N__14718),
            .I(N__14714));
    InMux I__2843 (
            .O(N__14717),
            .I(N__14711));
    IoSpan4Mux I__2842 (
            .O(N__14714),
            .I(N__14706));
    LocalMux I__2841 (
            .O(N__14711),
            .I(N__14703));
    InMux I__2840 (
            .O(N__14710),
            .I(N__14700));
    InMux I__2839 (
            .O(N__14709),
            .I(N__14697));
    Span4Mux_s3_h I__2838 (
            .O(N__14706),
            .I(N__14687));
    Span4Mux_v I__2837 (
            .O(N__14703),
            .I(N__14687));
    LocalMux I__2836 (
            .O(N__14700),
            .I(N__14687));
    LocalMux I__2835 (
            .O(N__14697),
            .I(N__14687));
    InMux I__2834 (
            .O(N__14696),
            .I(N__14684));
    Span4Mux_h I__2833 (
            .O(N__14687),
            .I(N__14678));
    LocalMux I__2832 (
            .O(N__14684),
            .I(N__14675));
    InMux I__2831 (
            .O(N__14683),
            .I(N__14672));
    InMux I__2830 (
            .O(N__14682),
            .I(N__14667));
    InMux I__2829 (
            .O(N__14681),
            .I(N__14667));
    Odrv4 I__2828 (
            .O(N__14678),
            .I(rsmrstn));
    Odrv12 I__2827 (
            .O(N__14675),
            .I(rsmrstn));
    LocalMux I__2826 (
            .O(N__14672),
            .I(rsmrstn));
    LocalMux I__2825 (
            .O(N__14667),
            .I(rsmrstn));
    InMux I__2824 (
            .O(N__14658),
            .I(N__14655));
    LocalMux I__2823 (
            .O(N__14655),
            .I(\POWERLED.dutycycle_s_1 ));
    InMux I__2822 (
            .O(N__14652),
            .I(N__14648));
    InMux I__2821 (
            .O(N__14651),
            .I(N__14641));
    LocalMux I__2820 (
            .O(N__14648),
            .I(N__14638));
    CascadeMux I__2819 (
            .O(N__14647),
            .I(N__14635));
    CascadeMux I__2818 (
            .O(N__14646),
            .I(N__14630));
    InMux I__2817 (
            .O(N__14645),
            .I(N__14625));
    InMux I__2816 (
            .O(N__14644),
            .I(N__14625));
    LocalMux I__2815 (
            .O(N__14641),
            .I(N__14622));
    Span4Mux_v I__2814 (
            .O(N__14638),
            .I(N__14619));
    InMux I__2813 (
            .O(N__14635),
            .I(N__14616));
    CascadeMux I__2812 (
            .O(N__14634),
            .I(N__14612));
    CascadeMux I__2811 (
            .O(N__14633),
            .I(N__14609));
    InMux I__2810 (
            .O(N__14630),
            .I(N__14606));
    LocalMux I__2809 (
            .O(N__14625),
            .I(N__14603));
    Span12Mux_s7_h I__2808 (
            .O(N__14622),
            .I(N__14600));
    Span4Mux_h I__2807 (
            .O(N__14619),
            .I(N__14595));
    LocalMux I__2806 (
            .O(N__14616),
            .I(N__14595));
    InMux I__2805 (
            .O(N__14615),
            .I(N__14588));
    InMux I__2804 (
            .O(N__14612),
            .I(N__14588));
    InMux I__2803 (
            .O(N__14609),
            .I(N__14588));
    LocalMux I__2802 (
            .O(N__14606),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__2801 (
            .O(N__14603),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv12 I__2800 (
            .O(N__14600),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__2799 (
            .O(N__14595),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__2798 (
            .O(N__14588),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    CascadeMux I__2797 (
            .O(N__14577),
            .I(N__14574));
    InMux I__2796 (
            .O(N__14574),
            .I(N__14571));
    LocalMux I__2795 (
            .O(N__14571),
            .I(N__14568));
    Odrv4 I__2794 (
            .O(N__14568),
            .I(\POWERLED.un1_dutycycle_1_axb_1 ));
    InMux I__2793 (
            .O(N__14565),
            .I(N__14559));
    InMux I__2792 (
            .O(N__14564),
            .I(N__14559));
    LocalMux I__2791 (
            .O(N__14559),
            .I(\POWERLED.N_53 ));
    CascadeMux I__2790 (
            .O(N__14556),
            .I(N__14553));
    InMux I__2789 (
            .O(N__14553),
            .I(N__14550));
    LocalMux I__2788 (
            .O(N__14550),
            .I(\POWERLED.dutycycle_s_0 ));
    InMux I__2787 (
            .O(N__14547),
            .I(N__14544));
    LocalMux I__2786 (
            .O(N__14544),
            .I(N__14540));
    CascadeMux I__2785 (
            .O(N__14543),
            .I(N__14536));
    Span4Mux_s3_h I__2784 (
            .O(N__14540),
            .I(N__14531));
    InMux I__2783 (
            .O(N__14539),
            .I(N__14526));
    InMux I__2782 (
            .O(N__14536),
            .I(N__14526));
    InMux I__2781 (
            .O(N__14535),
            .I(N__14523));
    InMux I__2780 (
            .O(N__14534),
            .I(N__14518));
    Span4Mux_h I__2779 (
            .O(N__14531),
            .I(N__14515));
    LocalMux I__2778 (
            .O(N__14526),
            .I(N__14512));
    LocalMux I__2777 (
            .O(N__14523),
            .I(N__14509));
    InMux I__2776 (
            .O(N__14522),
            .I(N__14504));
    InMux I__2775 (
            .O(N__14521),
            .I(N__14504));
    LocalMux I__2774 (
            .O(N__14518),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__2773 (
            .O(N__14515),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__2772 (
            .O(N__14512),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__2771 (
            .O(N__14509),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__2770 (
            .O(N__14504),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    InMux I__2769 (
            .O(N__14493),
            .I(N__14489));
    InMux I__2768 (
            .O(N__14492),
            .I(N__14486));
    LocalMux I__2767 (
            .O(N__14489),
            .I(N__14483));
    LocalMux I__2766 (
            .O(N__14486),
            .I(\POWERLED.dutycycle_s_5 ));
    Odrv4 I__2765 (
            .O(N__14483),
            .I(\POWERLED.dutycycle_s_5 ));
    CascadeMux I__2764 (
            .O(N__14478),
            .I(N__14470));
    CascadeMux I__2763 (
            .O(N__14477),
            .I(N__14467));
    InMux I__2762 (
            .O(N__14476),
            .I(N__14459));
    InMux I__2761 (
            .O(N__14475),
            .I(N__14459));
    InMux I__2760 (
            .O(N__14474),
            .I(N__14459));
    InMux I__2759 (
            .O(N__14473),
            .I(N__14454));
    InMux I__2758 (
            .O(N__14470),
            .I(N__14447));
    InMux I__2757 (
            .O(N__14467),
            .I(N__14447));
    InMux I__2756 (
            .O(N__14466),
            .I(N__14447));
    LocalMux I__2755 (
            .O(N__14459),
            .I(N__14443));
    InMux I__2754 (
            .O(N__14458),
            .I(N__14440));
    InMux I__2753 (
            .O(N__14457),
            .I(N__14437));
    LocalMux I__2752 (
            .O(N__14454),
            .I(N__14426));
    LocalMux I__2751 (
            .O(N__14447),
            .I(N__14423));
    InMux I__2750 (
            .O(N__14446),
            .I(N__14420));
    Span4Mux_h I__2749 (
            .O(N__14443),
            .I(N__14413));
    LocalMux I__2748 (
            .O(N__14440),
            .I(N__14413));
    LocalMux I__2747 (
            .O(N__14437),
            .I(N__14413));
    InMux I__2746 (
            .O(N__14436),
            .I(N__14404));
    InMux I__2745 (
            .O(N__14435),
            .I(N__14404));
    InMux I__2744 (
            .O(N__14434),
            .I(N__14404));
    InMux I__2743 (
            .O(N__14433),
            .I(N__14404));
    InMux I__2742 (
            .O(N__14432),
            .I(N__14395));
    InMux I__2741 (
            .O(N__14431),
            .I(N__14395));
    InMux I__2740 (
            .O(N__14430),
            .I(N__14395));
    InMux I__2739 (
            .O(N__14429),
            .I(N__14395));
    Odrv12 I__2738 (
            .O(N__14426),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    Odrv4 I__2737 (
            .O(N__14423),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    LocalMux I__2736 (
            .O(N__14420),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    Odrv4 I__2735 (
            .O(N__14413),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    LocalMux I__2734 (
            .O(N__14404),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    LocalMux I__2733 (
            .O(N__14395),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    InMux I__2732 (
            .O(N__14382),
            .I(N__14376));
    InMux I__2731 (
            .O(N__14381),
            .I(N__14376));
    LocalMux I__2730 (
            .O(N__14376),
            .I(N__14371));
    CascadeMux I__2729 (
            .O(N__14375),
            .I(N__14368));
    CascadeMux I__2728 (
            .O(N__14374),
            .I(N__14365));
    Span4Mux_v I__2727 (
            .O(N__14371),
            .I(N__14362));
    InMux I__2726 (
            .O(N__14368),
            .I(N__14359));
    InMux I__2725 (
            .O(N__14365),
            .I(N__14356));
    Odrv4 I__2724 (
            .O(N__14362),
            .I(\POWERLED.N_213 ));
    LocalMux I__2723 (
            .O(N__14359),
            .I(\POWERLED.N_213 ));
    LocalMux I__2722 (
            .O(N__14356),
            .I(\POWERLED.N_213 ));
    CascadeMux I__2721 (
            .O(N__14349),
            .I(N__14345));
    CascadeMux I__2720 (
            .O(N__14348),
            .I(N__14341));
    InMux I__2719 (
            .O(N__14345),
            .I(N__14334));
    InMux I__2718 (
            .O(N__14344),
            .I(N__14334));
    InMux I__2717 (
            .O(N__14341),
            .I(N__14334));
    LocalMux I__2716 (
            .O(N__14334),
            .I(N__14331));
    Odrv4 I__2715 (
            .O(N__14331),
            .I(\POWERLED.dutycycle_fastZ0Z_5 ));
    CascadeMux I__2714 (
            .O(N__14328),
            .I(N__14325));
    InMux I__2713 (
            .O(N__14325),
            .I(N__14315));
    InMux I__2712 (
            .O(N__14324),
            .I(N__14312));
    InMux I__2711 (
            .O(N__14323),
            .I(N__14309));
    InMux I__2710 (
            .O(N__14322),
            .I(N__14302));
    InMux I__2709 (
            .O(N__14321),
            .I(N__14302));
    InMux I__2708 (
            .O(N__14320),
            .I(N__14302));
    InMux I__2707 (
            .O(N__14319),
            .I(N__14297));
    InMux I__2706 (
            .O(N__14318),
            .I(N__14297));
    LocalMux I__2705 (
            .O(N__14315),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__2704 (
            .O(N__14312),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__2703 (
            .O(N__14309),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__2702 (
            .O(N__14302),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__2701 (
            .O(N__14297),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    CascadeMux I__2700 (
            .O(N__14286),
            .I(N__14281));
    CascadeMux I__2699 (
            .O(N__14285),
            .I(N__14278));
    InMux I__2698 (
            .O(N__14284),
            .I(N__14275));
    InMux I__2697 (
            .O(N__14281),
            .I(N__14270));
    InMux I__2696 (
            .O(N__14278),
            .I(N__14267));
    LocalMux I__2695 (
            .O(N__14275),
            .I(N__14264));
    CascadeMux I__2694 (
            .O(N__14274),
            .I(N__14260));
    CascadeMux I__2693 (
            .O(N__14273),
            .I(N__14257));
    LocalMux I__2692 (
            .O(N__14270),
            .I(N__14253));
    LocalMux I__2691 (
            .O(N__14267),
            .I(N__14248));
    Span4Mux_v I__2690 (
            .O(N__14264),
            .I(N__14248));
    InMux I__2689 (
            .O(N__14263),
            .I(N__14245));
    InMux I__2688 (
            .O(N__14260),
            .I(N__14242));
    InMux I__2687 (
            .O(N__14257),
            .I(N__14237));
    InMux I__2686 (
            .O(N__14256),
            .I(N__14237));
    Odrv4 I__2685 (
            .O(N__14253),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    Odrv4 I__2684 (
            .O(N__14248),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    LocalMux I__2683 (
            .O(N__14245),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    LocalMux I__2682 (
            .O(N__14242),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    LocalMux I__2681 (
            .O(N__14237),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    CascadeMux I__2680 (
            .O(N__14226),
            .I(N__14220));
    InMux I__2679 (
            .O(N__14225),
            .I(N__14215));
    CascadeMux I__2678 (
            .O(N__14224),
            .I(N__14212));
    InMux I__2677 (
            .O(N__14223),
            .I(N__14206));
    InMux I__2676 (
            .O(N__14220),
            .I(N__14206));
    CascadeMux I__2675 (
            .O(N__14219),
            .I(N__14203));
    CascadeMux I__2674 (
            .O(N__14218),
            .I(N__14200));
    LocalMux I__2673 (
            .O(N__14215),
            .I(N__14194));
    InMux I__2672 (
            .O(N__14212),
            .I(N__14191));
    InMux I__2671 (
            .O(N__14211),
            .I(N__14188));
    LocalMux I__2670 (
            .O(N__14206),
            .I(N__14185));
    InMux I__2669 (
            .O(N__14203),
            .I(N__14174));
    InMux I__2668 (
            .O(N__14200),
            .I(N__14174));
    InMux I__2667 (
            .O(N__14199),
            .I(N__14174));
    InMux I__2666 (
            .O(N__14198),
            .I(N__14174));
    InMux I__2665 (
            .O(N__14197),
            .I(N__14174));
    Odrv4 I__2664 (
            .O(N__14194),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__2663 (
            .O(N__14191),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__2662 (
            .O(N__14188),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__2661 (
            .O(N__14185),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__2660 (
            .O(N__14174),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    CascadeMux I__2659 (
            .O(N__14163),
            .I(N__14159));
    InMux I__2658 (
            .O(N__14162),
            .I(N__14156));
    InMux I__2657 (
            .O(N__14159),
            .I(N__14153));
    LocalMux I__2656 (
            .O(N__14156),
            .I(N__14146));
    LocalMux I__2655 (
            .O(N__14153),
            .I(N__14143));
    CascadeMux I__2654 (
            .O(N__14152),
            .I(N__14140));
    InMux I__2653 (
            .O(N__14151),
            .I(N__14135));
    InMux I__2652 (
            .O(N__14150),
            .I(N__14132));
    InMux I__2651 (
            .O(N__14149),
            .I(N__14129));
    Span4Mux_h I__2650 (
            .O(N__14146),
            .I(N__14124));
    Span4Mux_h I__2649 (
            .O(N__14143),
            .I(N__14124));
    InMux I__2648 (
            .O(N__14140),
            .I(N__14121));
    InMux I__2647 (
            .O(N__14139),
            .I(N__14116));
    InMux I__2646 (
            .O(N__14138),
            .I(N__14116));
    LocalMux I__2645 (
            .O(N__14135),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__2644 (
            .O(N__14132),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__2643 (
            .O(N__14129),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__2642 (
            .O(N__14124),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__2641 (
            .O(N__14121),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__2640 (
            .O(N__14116),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    InMux I__2639 (
            .O(N__14103),
            .I(N__14099));
    InMux I__2638 (
            .O(N__14102),
            .I(N__14096));
    LocalMux I__2637 (
            .O(N__14099),
            .I(N__14092));
    LocalMux I__2636 (
            .O(N__14096),
            .I(N__14089));
    CascadeMux I__2635 (
            .O(N__14095),
            .I(N__14084));
    Span4Mux_v I__2634 (
            .O(N__14092),
            .I(N__14078));
    Span4Mux_s2_h I__2633 (
            .O(N__14089),
            .I(N__14078));
    CascadeMux I__2632 (
            .O(N__14088),
            .I(N__14074));
    CascadeMux I__2631 (
            .O(N__14087),
            .I(N__14071));
    InMux I__2630 (
            .O(N__14084),
            .I(N__14067));
    InMux I__2629 (
            .O(N__14083),
            .I(N__14064));
    Span4Mux_h I__2628 (
            .O(N__14078),
            .I(N__14061));
    InMux I__2627 (
            .O(N__14077),
            .I(N__14058));
    InMux I__2626 (
            .O(N__14074),
            .I(N__14053));
    InMux I__2625 (
            .O(N__14071),
            .I(N__14053));
    InMux I__2624 (
            .O(N__14070),
            .I(N__14050));
    LocalMux I__2623 (
            .O(N__14067),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__2622 (
            .O(N__14064),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__2621 (
            .O(N__14061),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__2620 (
            .O(N__14058),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__2619 (
            .O(N__14053),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__2618 (
            .O(N__14050),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    CascadeMux I__2617 (
            .O(N__14037),
            .I(N__14030));
    InMux I__2616 (
            .O(N__14036),
            .I(N__14025));
    CascadeMux I__2615 (
            .O(N__14035),
            .I(N__14021));
    CascadeMux I__2614 (
            .O(N__14034),
            .I(N__14018));
    InMux I__2613 (
            .O(N__14033),
            .I(N__14014));
    InMux I__2612 (
            .O(N__14030),
            .I(N__14011));
    InMux I__2611 (
            .O(N__14029),
            .I(N__14008));
    InMux I__2610 (
            .O(N__14028),
            .I(N__14005));
    LocalMux I__2609 (
            .O(N__14025),
            .I(N__14002));
    InMux I__2608 (
            .O(N__14024),
            .I(N__13997));
    InMux I__2607 (
            .O(N__14021),
            .I(N__13997));
    InMux I__2606 (
            .O(N__14018),
            .I(N__13992));
    InMux I__2605 (
            .O(N__14017),
            .I(N__13992));
    LocalMux I__2604 (
            .O(N__14014),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__2603 (
            .O(N__14011),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__2602 (
            .O(N__14008),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__2601 (
            .O(N__14005),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    Odrv4 I__2600 (
            .O(N__14002),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__2599 (
            .O(N__13997),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__2598 (
            .O(N__13992),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    InMux I__2597 (
            .O(N__13977),
            .I(N__13971));
    CascadeMux I__2596 (
            .O(N__13976),
            .I(N__13967));
    CascadeMux I__2595 (
            .O(N__13975),
            .I(N__13961));
    CascadeMux I__2594 (
            .O(N__13974),
            .I(N__13957));
    LocalMux I__2593 (
            .O(N__13971),
            .I(N__13954));
    InMux I__2592 (
            .O(N__13970),
            .I(N__13949));
    InMux I__2591 (
            .O(N__13967),
            .I(N__13946));
    InMux I__2590 (
            .O(N__13966),
            .I(N__13943));
    InMux I__2589 (
            .O(N__13965),
            .I(N__13940));
    InMux I__2588 (
            .O(N__13964),
            .I(N__13935));
    InMux I__2587 (
            .O(N__13961),
            .I(N__13935));
    InMux I__2586 (
            .O(N__13960),
            .I(N__13930));
    InMux I__2585 (
            .O(N__13957),
            .I(N__13930));
    Span4Mux_h I__2584 (
            .O(N__13954),
            .I(N__13927));
    InMux I__2583 (
            .O(N__13953),
            .I(N__13922));
    InMux I__2582 (
            .O(N__13952),
            .I(N__13922));
    LocalMux I__2581 (
            .O(N__13949),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__2580 (
            .O(N__13946),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__2579 (
            .O(N__13943),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__2578 (
            .O(N__13940),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__2577 (
            .O(N__13935),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__2576 (
            .O(N__13930),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    Odrv4 I__2575 (
            .O(N__13927),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__2574 (
            .O(N__13922),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    CascadeMux I__2573 (
            .O(N__13905),
            .I(N__13897));
    CascadeMux I__2572 (
            .O(N__13904),
            .I(N__13890));
    InMux I__2571 (
            .O(N__13903),
            .I(N__13887));
    InMux I__2570 (
            .O(N__13902),
            .I(N__13882));
    InMux I__2569 (
            .O(N__13901),
            .I(N__13882));
    InMux I__2568 (
            .O(N__13900),
            .I(N__13879));
    InMux I__2567 (
            .O(N__13897),
            .I(N__13874));
    InMux I__2566 (
            .O(N__13896),
            .I(N__13874));
    InMux I__2565 (
            .O(N__13895),
            .I(N__13865));
    InMux I__2564 (
            .O(N__13894),
            .I(N__13865));
    InMux I__2563 (
            .O(N__13893),
            .I(N__13865));
    InMux I__2562 (
            .O(N__13890),
            .I(N__13865));
    LocalMux I__2561 (
            .O(N__13887),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__2560 (
            .O(N__13882),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__2559 (
            .O(N__13879),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__2558 (
            .O(N__13874),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__2557 (
            .O(N__13865),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    CascadeMux I__2556 (
            .O(N__13854),
            .I(\POWERLED.un1_dutycycle_1_44_0_cascade_ ));
    CascadeMux I__2555 (
            .O(N__13851),
            .I(N__13848));
    InMux I__2554 (
            .O(N__13848),
            .I(N__13845));
    LocalMux I__2553 (
            .O(N__13845),
            .I(N__13842));
    Odrv4 I__2552 (
            .O(N__13842),
            .I(\POWERLED.dutycycle_RNIF3561Z0Z_9 ));
    InMux I__2551 (
            .O(N__13839),
            .I(\COUNTER.counter_1_cry_30 ));
    CascadeMux I__2550 (
            .O(N__13836),
            .I(N__13833));
    InMux I__2549 (
            .O(N__13833),
            .I(N__13827));
    InMux I__2548 (
            .O(N__13832),
            .I(N__13827));
    LocalMux I__2547 (
            .O(N__13827),
            .I(\COUNTER.counterZ0Z_30 ));
    CascadeMux I__2546 (
            .O(N__13824),
            .I(N__13821));
    InMux I__2545 (
            .O(N__13821),
            .I(N__13815));
    InMux I__2544 (
            .O(N__13820),
            .I(N__13815));
    LocalMux I__2543 (
            .O(N__13815),
            .I(\COUNTER.counterZ0Z_29 ));
    CascadeMux I__2542 (
            .O(N__13812),
            .I(N__13808));
    InMux I__2541 (
            .O(N__13811),
            .I(N__13803));
    InMux I__2540 (
            .O(N__13808),
            .I(N__13803));
    LocalMux I__2539 (
            .O(N__13803),
            .I(\COUNTER.counterZ0Z_31 ));
    InMux I__2538 (
            .O(N__13800),
            .I(N__13794));
    InMux I__2537 (
            .O(N__13799),
            .I(N__13794));
    LocalMux I__2536 (
            .O(N__13794),
            .I(\COUNTER.counterZ0Z_28 ));
    InMux I__2535 (
            .O(N__13791),
            .I(N__13787));
    InMux I__2534 (
            .O(N__13790),
            .I(N__13784));
    LocalMux I__2533 (
            .O(N__13787),
            .I(\POWERLED.N_234 ));
    LocalMux I__2532 (
            .O(N__13784),
            .I(\POWERLED.N_234 ));
    CascadeMux I__2531 (
            .O(N__13779),
            .I(\POWERLED.N_248_cascade_ ));
    InMux I__2530 (
            .O(N__13776),
            .I(N__13770));
    InMux I__2529 (
            .O(N__13775),
            .I(N__13770));
    LocalMux I__2528 (
            .O(N__13770),
            .I(\POWERLED.N_118 ));
    InMux I__2527 (
            .O(N__13767),
            .I(N__13764));
    LocalMux I__2526 (
            .O(N__13764),
            .I(N__13761));
    Odrv12 I__2525 (
            .O(N__13761),
            .I(\POWERLED.dutycycle_RNIFHLJZ0Z_0 ));
    InMux I__2524 (
            .O(N__13758),
            .I(N__13752));
    CascadeMux I__2523 (
            .O(N__13757),
            .I(N__13749));
    CascadeMux I__2522 (
            .O(N__13756),
            .I(N__13745));
    CascadeMux I__2521 (
            .O(N__13755),
            .I(N__13742));
    LocalMux I__2520 (
            .O(N__13752),
            .I(N__13738));
    InMux I__2519 (
            .O(N__13749),
            .I(N__13733));
    InMux I__2518 (
            .O(N__13748),
            .I(N__13733));
    InMux I__2517 (
            .O(N__13745),
            .I(N__13728));
    InMux I__2516 (
            .O(N__13742),
            .I(N__13728));
    InMux I__2515 (
            .O(N__13741),
            .I(N__13725));
    Odrv12 I__2514 (
            .O(N__13738),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__2513 (
            .O(N__13733),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__2512 (
            .O(N__13728),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__2511 (
            .O(N__13725),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    CascadeMux I__2510 (
            .O(N__13716),
            .I(\POWERLED.dutycycle_RNIFHLJZ0Z_0_cascade_ ));
    CascadeMux I__2509 (
            .O(N__13713),
            .I(N__13710));
    InMux I__2508 (
            .O(N__13710),
            .I(N__13707));
    LocalMux I__2507 (
            .O(N__13707),
            .I(N__13704));
    Odrv12 I__2506 (
            .O(N__13704),
            .I(\POWERLED.dutycycle_RNI16B71Z0Z_5 ));
    InMux I__2505 (
            .O(N__13701),
            .I(\COUNTER.counter_1_cry_21 ));
    InMux I__2504 (
            .O(N__13698),
            .I(\COUNTER.counter_1_cry_22 ));
    InMux I__2503 (
            .O(N__13695),
            .I(\COUNTER.counter_1_cry_23 ));
    InMux I__2502 (
            .O(N__13692),
            .I(bfn_8_8_0_));
    InMux I__2501 (
            .O(N__13689),
            .I(\COUNTER.counter_1_cry_25 ));
    InMux I__2500 (
            .O(N__13686),
            .I(\COUNTER.counter_1_cry_26 ));
    InMux I__2499 (
            .O(N__13683),
            .I(\COUNTER.counter_1_cry_27 ));
    InMux I__2498 (
            .O(N__13680),
            .I(\COUNTER.counter_1_cry_28 ));
    InMux I__2497 (
            .O(N__13677),
            .I(\COUNTER.counter_1_cry_29 ));
    InMux I__2496 (
            .O(N__13674),
            .I(\COUNTER.counter_1_cry_12 ));
    InMux I__2495 (
            .O(N__13671),
            .I(\COUNTER.counter_1_cry_13 ));
    InMux I__2494 (
            .O(N__13668),
            .I(\COUNTER.counter_1_cry_14 ));
    InMux I__2493 (
            .O(N__13665),
            .I(\COUNTER.counter_1_cry_15 ));
    InMux I__2492 (
            .O(N__13662),
            .I(bfn_8_7_0_));
    InMux I__2491 (
            .O(N__13659),
            .I(\COUNTER.counter_1_cry_17 ));
    InMux I__2490 (
            .O(N__13656),
            .I(\COUNTER.counter_1_cry_18 ));
    InMux I__2489 (
            .O(N__13653),
            .I(\COUNTER.counter_1_cry_19 ));
    InMux I__2488 (
            .O(N__13650),
            .I(\COUNTER.counter_1_cry_20 ));
    CascadeMux I__2487 (
            .O(N__13647),
            .I(N__13642));
    InMux I__2486 (
            .O(N__13646),
            .I(N__13639));
    InMux I__2485 (
            .O(N__13645),
            .I(N__13634));
    InMux I__2484 (
            .O(N__13642),
            .I(N__13634));
    LocalMux I__2483 (
            .O(N__13639),
            .I(\COUNTER.counterZ0Z_4 ));
    LocalMux I__2482 (
            .O(N__13634),
            .I(\COUNTER.counterZ0Z_4 ));
    InMux I__2481 (
            .O(N__13629),
            .I(N__13626));
    LocalMux I__2480 (
            .O(N__13626),
            .I(\COUNTER.counter_1_cry_3_THRU_CO ));
    InMux I__2479 (
            .O(N__13623),
            .I(\COUNTER.counter_1_cry_3 ));
    InMux I__2478 (
            .O(N__13620),
            .I(\COUNTER.counter_1_cry_4 ));
    InMux I__2477 (
            .O(N__13617),
            .I(\COUNTER.counter_1_cry_5 ));
    InMux I__2476 (
            .O(N__13614),
            .I(\COUNTER.counter_1_cry_6 ));
    InMux I__2475 (
            .O(N__13611),
            .I(\COUNTER.counter_1_cry_7 ));
    InMux I__2474 (
            .O(N__13608),
            .I(bfn_8_6_0_));
    InMux I__2473 (
            .O(N__13605),
            .I(\COUNTER.counter_1_cry_9 ));
    InMux I__2472 (
            .O(N__13602),
            .I(\COUNTER.counter_1_cry_10 ));
    InMux I__2471 (
            .O(N__13599),
            .I(\COUNTER.counter_1_cry_11 ));
    InMux I__2470 (
            .O(N__13596),
            .I(bfn_8_3_0_));
    CEMux I__2469 (
            .O(N__13593),
            .I(N__13590));
    LocalMux I__2468 (
            .O(N__13590),
            .I(N__13587));
    Span4Mux_s2_v I__2467 (
            .O(N__13587),
            .I(N__13584));
    Odrv4 I__2466 (
            .O(N__13584),
            .I(\PCH_PWRGD.N_49_3 ));
    SRMux I__2465 (
            .O(N__13581),
            .I(N__13577));
    SRMux I__2464 (
            .O(N__13580),
            .I(N__13572));
    LocalMux I__2463 (
            .O(N__13577),
            .I(N__13569));
    SRMux I__2462 (
            .O(N__13576),
            .I(N__13566));
    InMux I__2461 (
            .O(N__13575),
            .I(N__13563));
    LocalMux I__2460 (
            .O(N__13572),
            .I(N__13560));
    Span4Mux_h I__2459 (
            .O(N__13569),
            .I(N__13557));
    LocalMux I__2458 (
            .O(N__13566),
            .I(N__13554));
    LocalMux I__2457 (
            .O(N__13563),
            .I(N__13551));
    Odrv4 I__2456 (
            .O(N__13560),
            .I(\PCH_PWRGD.curr_state_RNI7N705Z0Z_0 ));
    Odrv4 I__2455 (
            .O(N__13557),
            .I(\PCH_PWRGD.curr_state_RNI7N705Z0Z_0 ));
    Odrv4 I__2454 (
            .O(N__13554),
            .I(\PCH_PWRGD.curr_state_RNI7N705Z0Z_0 ));
    Odrv4 I__2453 (
            .O(N__13551),
            .I(\PCH_PWRGD.curr_state_RNI7N705Z0Z_0 ));
    InMux I__2452 (
            .O(N__13542),
            .I(N__13537));
    InMux I__2451 (
            .O(N__13541),
            .I(N__13532));
    InMux I__2450 (
            .O(N__13540),
            .I(N__13532));
    LocalMux I__2449 (
            .O(N__13537),
            .I(\COUNTER.counterZ0Z_2 ));
    LocalMux I__2448 (
            .O(N__13532),
            .I(\COUNTER.counterZ0Z_2 ));
    InMux I__2447 (
            .O(N__13527),
            .I(N__13524));
    LocalMux I__2446 (
            .O(N__13524),
            .I(\COUNTER.counter_1_cry_1_THRU_CO ));
    InMux I__2445 (
            .O(N__13521),
            .I(\COUNTER.counter_1_cry_1 ));
    InMux I__2444 (
            .O(N__13518),
            .I(N__13513));
    InMux I__2443 (
            .O(N__13517),
            .I(N__13508));
    InMux I__2442 (
            .O(N__13516),
            .I(N__13508));
    LocalMux I__2441 (
            .O(N__13513),
            .I(\COUNTER.counterZ0Z_3 ));
    LocalMux I__2440 (
            .O(N__13508),
            .I(\COUNTER.counterZ0Z_3 ));
    InMux I__2439 (
            .O(N__13503),
            .I(N__13500));
    LocalMux I__2438 (
            .O(N__13500),
            .I(\COUNTER.counter_1_cry_2_THRU_CO ));
    InMux I__2437 (
            .O(N__13497),
            .I(\COUNTER.counter_1_cry_2 ));
    InMux I__2436 (
            .O(N__13494),
            .I(\PCH_PWRGD.un1_count_1_cry_5 ));
    InMux I__2435 (
            .O(N__13491),
            .I(\PCH_PWRGD.un1_count_1_cry_6 ));
    InMux I__2434 (
            .O(N__13488),
            .I(bfn_8_2_0_));
    InMux I__2433 (
            .O(N__13485),
            .I(\PCH_PWRGD.un1_count_1_cry_8 ));
    InMux I__2432 (
            .O(N__13482),
            .I(\PCH_PWRGD.un1_count_1_cry_9 ));
    InMux I__2431 (
            .O(N__13479),
            .I(\PCH_PWRGD.un1_count_1_cry_10 ));
    InMux I__2430 (
            .O(N__13476),
            .I(\PCH_PWRGD.un1_count_1_cry_11 ));
    InMux I__2429 (
            .O(N__13473),
            .I(\PCH_PWRGD.un1_count_1_cry_12 ));
    InMux I__2428 (
            .O(N__13470),
            .I(\PCH_PWRGD.un1_count_1_cry_13 ));
    InMux I__2427 (
            .O(N__13467),
            .I(N__13463));
    InMux I__2426 (
            .O(N__13466),
            .I(N__13460));
    LocalMux I__2425 (
            .O(N__13463),
            .I(N__13455));
    LocalMux I__2424 (
            .O(N__13460),
            .I(N__13455));
    Odrv4 I__2423 (
            .O(N__13455),
            .I(\VPP_VDDQ.count_esr_RNIRFM64Z0Z_15 ));
    InMux I__2422 (
            .O(N__13452),
            .I(N__13442));
    InMux I__2421 (
            .O(N__13451),
            .I(N__13442));
    InMux I__2420 (
            .O(N__13450),
            .I(N__13433));
    InMux I__2419 (
            .O(N__13449),
            .I(N__13433));
    InMux I__2418 (
            .O(N__13448),
            .I(N__13433));
    InMux I__2417 (
            .O(N__13447),
            .I(N__13433));
    LocalMux I__2416 (
            .O(N__13442),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    LocalMux I__2415 (
            .O(N__13433),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    InMux I__2414 (
            .O(N__13428),
            .I(N__13420));
    InMux I__2413 (
            .O(N__13427),
            .I(N__13413));
    InMux I__2412 (
            .O(N__13426),
            .I(N__13413));
    InMux I__2411 (
            .O(N__13425),
            .I(N__13413));
    InMux I__2410 (
            .O(N__13424),
            .I(N__13408));
    InMux I__2409 (
            .O(N__13423),
            .I(N__13408));
    LocalMux I__2408 (
            .O(N__13420),
            .I(VPP_VDDQ_curr_state_0));
    LocalMux I__2407 (
            .O(N__13413),
            .I(VPP_VDDQ_curr_state_0));
    LocalMux I__2406 (
            .O(N__13408),
            .I(VPP_VDDQ_curr_state_0));
    InMux I__2405 (
            .O(N__13401),
            .I(N__13397));
    CascadeMux I__2404 (
            .O(N__13400),
            .I(N__13394));
    LocalMux I__2403 (
            .O(N__13397),
            .I(N__13391));
    InMux I__2402 (
            .O(N__13394),
            .I(N__13388));
    Odrv4 I__2401 (
            .O(N__13391),
            .I(\PCH_PWRGD.un1_curr_state10_0 ));
    LocalMux I__2400 (
            .O(N__13388),
            .I(\PCH_PWRGD.un1_curr_state10_0 ));
    InMux I__2399 (
            .O(N__13383),
            .I(\PCH_PWRGD.un1_count_1_cry_0 ));
    InMux I__2398 (
            .O(N__13380),
            .I(\PCH_PWRGD.un1_count_1_cry_1 ));
    InMux I__2397 (
            .O(N__13377),
            .I(\PCH_PWRGD.un1_count_1_cry_2 ));
    InMux I__2396 (
            .O(N__13374),
            .I(\PCH_PWRGD.un1_count_1_cry_3 ));
    InMux I__2395 (
            .O(N__13371),
            .I(\PCH_PWRGD.un1_count_1_cry_4 ));
    InMux I__2394 (
            .O(N__13368),
            .I(bfn_7_12_0_));
    InMux I__2393 (
            .O(N__13365),
            .I(\POWERLED.dutycycle_cry_7 ));
    InMux I__2392 (
            .O(N__13362),
            .I(\POWERLED.dutycycle_cry_8 ));
    InMux I__2391 (
            .O(N__13359),
            .I(\POWERLED.dutycycle_cry_9 ));
    InMux I__2390 (
            .O(N__13356),
            .I(\POWERLED.dutycycle_cry_10 ));
    InMux I__2389 (
            .O(N__13353),
            .I(\POWERLED.dutycycle_cry_11 ));
    InMux I__2388 (
            .O(N__13350),
            .I(\POWERLED.dutycycle_cry_12 ));
    InMux I__2387 (
            .O(N__13347),
            .I(\POWERLED.dutycycle_cry_13 ));
    InMux I__2386 (
            .O(N__13344),
            .I(bfn_7_13_0_));
    InMux I__2385 (
            .O(N__13341),
            .I(N__13336));
    InMux I__2384 (
            .O(N__13340),
            .I(N__13331));
    InMux I__2383 (
            .O(N__13339),
            .I(N__13331));
    LocalMux I__2382 (
            .O(N__13336),
            .I(\POWERLED.dutycycle_fastZ0Z_6 ));
    LocalMux I__2381 (
            .O(N__13331),
            .I(\POWERLED.dutycycle_fastZ0Z_6 ));
    CascadeMux I__2380 (
            .O(N__13326),
            .I(N__13323));
    InMux I__2379 (
            .O(N__13323),
            .I(N__13319));
    InMux I__2378 (
            .O(N__13322),
            .I(N__13316));
    LocalMux I__2377 (
            .O(N__13319),
            .I(N__13313));
    LocalMux I__2376 (
            .O(N__13316),
            .I(\POWERLED.dutycycle_fast_RNIBPSKZ0Z_6 ));
    Odrv4 I__2375 (
            .O(N__13313),
            .I(\POWERLED.dutycycle_fast_RNIBPSKZ0Z_6 ));
    CascadeMux I__2374 (
            .O(N__13308),
            .I(N__13305));
    InMux I__2373 (
            .O(N__13305),
            .I(N__13301));
    InMux I__2372 (
            .O(N__13304),
            .I(N__13298));
    LocalMux I__2371 (
            .O(N__13301),
            .I(N__13293));
    LocalMux I__2370 (
            .O(N__13298),
            .I(N__13293));
    Odrv4 I__2369 (
            .O(N__13293),
            .I(\POWERLED.dutycycle ));
    InMux I__2368 (
            .O(N__13290),
            .I(\POWERLED.dutycycle_cry_c_0_THRU_CO ));
    InMux I__2367 (
            .O(N__13287),
            .I(\POWERLED.dutycycle_cry_0 ));
    CascadeMux I__2366 (
            .O(N__13284),
            .I(N__13281));
    InMux I__2365 (
            .O(N__13281),
            .I(N__13278));
    LocalMux I__2364 (
            .O(N__13278),
            .I(\POWERLED.dutycycle_s_2 ));
    InMux I__2363 (
            .O(N__13275),
            .I(\POWERLED.dutycycle_cry_1 ));
    InMux I__2362 (
            .O(N__13272),
            .I(\POWERLED.dutycycle_cry_2 ));
    InMux I__2361 (
            .O(N__13269),
            .I(\POWERLED.dutycycle_cry_3 ));
    InMux I__2360 (
            .O(N__13266),
            .I(\POWERLED.dutycycle_cry_4 ));
    CascadeMux I__2359 (
            .O(N__13263),
            .I(N__13258));
    InMux I__2358 (
            .O(N__13262),
            .I(N__13253));
    InMux I__2357 (
            .O(N__13261),
            .I(N__13253));
    InMux I__2356 (
            .O(N__13258),
            .I(N__13246));
    LocalMux I__2355 (
            .O(N__13253),
            .I(N__13243));
    InMux I__2354 (
            .O(N__13252),
            .I(N__13238));
    InMux I__2353 (
            .O(N__13251),
            .I(N__13238));
    InMux I__2352 (
            .O(N__13250),
            .I(N__13233));
    InMux I__2351 (
            .O(N__13249),
            .I(N__13233));
    LocalMux I__2350 (
            .O(N__13246),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__2349 (
            .O(N__13243),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__2348 (
            .O(N__13238),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__2347 (
            .O(N__13233),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    InMux I__2346 (
            .O(N__13224),
            .I(N__13218));
    InMux I__2345 (
            .O(N__13223),
            .I(N__13218));
    LocalMux I__2344 (
            .O(N__13218),
            .I(\POWERLED.dutycycle_s_6 ));
    InMux I__2343 (
            .O(N__13215),
            .I(\POWERLED.dutycycle_cry_5 ));
    InMux I__2342 (
            .O(N__13212),
            .I(N__13208));
    CascadeMux I__2341 (
            .O(N__13211),
            .I(N__13205));
    LocalMux I__2340 (
            .O(N__13208),
            .I(N__13202));
    InMux I__2339 (
            .O(N__13205),
            .I(N__13199));
    Span4Mux_h I__2338 (
            .O(N__13202),
            .I(N__13196));
    LocalMux I__2337 (
            .O(N__13199),
            .I(N__13193));
    Odrv4 I__2336 (
            .O(N__13196),
            .I(\POWERLED.mult1_un82_sum ));
    Odrv4 I__2335 (
            .O(N__13193),
            .I(\POWERLED.mult1_un82_sum ));
    InMux I__2334 (
            .O(N__13188),
            .I(N__13185));
    LocalMux I__2333 (
            .O(N__13185),
            .I(\POWERLED.mult1_un82_sum_i ));
    CascadeMux I__2332 (
            .O(N__13182),
            .I(N__13178));
    InMux I__2331 (
            .O(N__13181),
            .I(N__13175));
    InMux I__2330 (
            .O(N__13178),
            .I(N__13172));
    LocalMux I__2329 (
            .O(N__13175),
            .I(\POWERLED.dutycycle_fast_RNI8MSKZ0Z_5 ));
    LocalMux I__2328 (
            .O(N__13172),
            .I(\POWERLED.dutycycle_fast_RNI8MSKZ0Z_5 ));
    InMux I__2327 (
            .O(N__13167),
            .I(N__13164));
    LocalMux I__2326 (
            .O(N__13164),
            .I(N__13161));
    Odrv4 I__2325 (
            .O(N__13161),
            .I(\POWERLED.dutycycle_RNI6NI81Z0Z_5 ));
    InMux I__2324 (
            .O(N__13158),
            .I(N__13154));
    CascadeMux I__2323 (
            .O(N__13157),
            .I(N__13151));
    LocalMux I__2322 (
            .O(N__13154),
            .I(N__13148));
    InMux I__2321 (
            .O(N__13151),
            .I(N__13145));
    Odrv4 I__2320 (
            .O(N__13148),
            .I(\POWERLED.dutycycle_fast_RNIVCSKZ0Z_5 ));
    LocalMux I__2319 (
            .O(N__13145),
            .I(\POWERLED.dutycycle_fast_RNIVCSKZ0Z_5 ));
    InMux I__2318 (
            .O(N__13140),
            .I(N__13137));
    LocalMux I__2317 (
            .O(N__13137),
            .I(N__13134));
    Odrv4 I__2316 (
            .O(N__13134),
            .I(\POWERLED.dutycycle_RNIK4I81Z0Z_6 ));
    CascadeMux I__2315 (
            .O(N__13131),
            .I(N__13128));
    InMux I__2314 (
            .O(N__13128),
            .I(N__13124));
    InMux I__2313 (
            .O(N__13127),
            .I(N__13121));
    LocalMux I__2312 (
            .O(N__13124),
            .I(N__13118));
    LocalMux I__2311 (
            .O(N__13121),
            .I(\POWERLED.dutycycle_fast_RNI2GSKZ0Z_6 ));
    Odrv4 I__2310 (
            .O(N__13118),
            .I(\POWERLED.dutycycle_fast_RNI2GSKZ0Z_6 ));
    InMux I__2309 (
            .O(N__13113),
            .I(N__13102));
    InMux I__2308 (
            .O(N__13112),
            .I(N__13102));
    InMux I__2307 (
            .O(N__13111),
            .I(N__13102));
    InMux I__2306 (
            .O(N__13110),
            .I(N__13097));
    InMux I__2305 (
            .O(N__13109),
            .I(N__13097));
    LocalMux I__2304 (
            .O(N__13102),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__2303 (
            .O(N__13097),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    InMux I__2302 (
            .O(N__13092),
            .I(N__13087));
    InMux I__2301 (
            .O(N__13091),
            .I(N__13082));
    InMux I__2300 (
            .O(N__13090),
            .I(N__13082));
    LocalMux I__2299 (
            .O(N__13087),
            .I(\PCH_PWRGD.N_3_i ));
    LocalMux I__2298 (
            .O(N__13082),
            .I(\PCH_PWRGD.N_3_i ));
    CascadeMux I__2297 (
            .O(N__13077),
            .I(N__13070));
    InMux I__2296 (
            .O(N__13076),
            .I(N__13063));
    InMux I__2295 (
            .O(N__13075),
            .I(N__13063));
    InMux I__2294 (
            .O(N__13074),
            .I(N__13063));
    InMux I__2293 (
            .O(N__13073),
            .I(N__13060));
    InMux I__2292 (
            .O(N__13070),
            .I(N__13057));
    LocalMux I__2291 (
            .O(N__13063),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__2290 (
            .O(N__13060),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__2289 (
            .O(N__13057),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    IoInMux I__2288 (
            .O(N__13050),
            .I(N__13047));
    LocalMux I__2287 (
            .O(N__13047),
            .I(N__13044));
    IoSpan4Mux I__2286 (
            .O(N__13044),
            .I(N__13041));
    Span4Mux_s3_h I__2285 (
            .O(N__13041),
            .I(N__13038));
    Sp12to4 I__2284 (
            .O(N__13038),
            .I(N__13034));
    IoInMux I__2283 (
            .O(N__13037),
            .I(N__13031));
    Span12Mux_v I__2282 (
            .O(N__13034),
            .I(N__13026));
    LocalMux I__2281 (
            .O(N__13031),
            .I(N__13026));
    Odrv12 I__2280 (
            .O(N__13026),
            .I(pch_pwrok));
    InMux I__2279 (
            .O(N__13023),
            .I(N__13020));
    LocalMux I__2278 (
            .O(N__13020),
            .I(N__13016));
    CascadeMux I__2277 (
            .O(N__13019),
            .I(N__13013));
    Span4Mux_h I__2276 (
            .O(N__13016),
            .I(N__13010));
    InMux I__2275 (
            .O(N__13013),
            .I(N__13007));
    Sp12to4 I__2274 (
            .O(N__13010),
            .I(N__13002));
    LocalMux I__2273 (
            .O(N__13007),
            .I(N__13002));
    Odrv12 I__2272 (
            .O(N__13002),
            .I(\POWERLED.mult1_un96_sum ));
    InMux I__2271 (
            .O(N__12999),
            .I(N__12996));
    LocalMux I__2270 (
            .O(N__12996),
            .I(N__12993));
    Odrv4 I__2269 (
            .O(N__12993),
            .I(\POWERLED.mult1_un96_sum_i ));
    InMux I__2268 (
            .O(N__12990),
            .I(N__12986));
    InMux I__2267 (
            .O(N__12989),
            .I(N__12983));
    LocalMux I__2266 (
            .O(N__12986),
            .I(N__12978));
    LocalMux I__2265 (
            .O(N__12983),
            .I(N__12978));
    Span4Mux_h I__2264 (
            .O(N__12978),
            .I(N__12975));
    Odrv4 I__2263 (
            .O(N__12975),
            .I(\POWERLED.mult1_un89_sum ));
    InMux I__2262 (
            .O(N__12972),
            .I(N__12969));
    LocalMux I__2261 (
            .O(N__12969),
            .I(N__12966));
    Odrv4 I__2260 (
            .O(N__12966),
            .I(\POWERLED.mult1_un89_sum_i ));
    InMux I__2259 (
            .O(N__12963),
            .I(N__12960));
    LocalMux I__2258 (
            .O(N__12960),
            .I(\POWERLED.N_117 ));
    CascadeMux I__2257 (
            .O(N__12957),
            .I(\POWERLED.N_117_cascade_ ));
    CascadeMux I__2256 (
            .O(N__12954),
            .I(N_154_cascade_));
    InMux I__2255 (
            .O(N__12951),
            .I(N__12948));
    LocalMux I__2254 (
            .O(N__12948),
            .I(N_128));
    CascadeMux I__2253 (
            .O(N__12945),
            .I(N_128_cascade_));
    InMux I__2252 (
            .O(N__12942),
            .I(N__12939));
    LocalMux I__2251 (
            .O(N__12939),
            .I(\VPP_VDDQ.delayed_vddq_pwrgd_0 ));
    SRMux I__2250 (
            .O(N__12936),
            .I(N__12930));
    SRMux I__2249 (
            .O(N__12935),
            .I(N__12927));
    SRMux I__2248 (
            .O(N__12934),
            .I(N__12924));
    InMux I__2247 (
            .O(N__12933),
            .I(N__12921));
    LocalMux I__2246 (
            .O(N__12930),
            .I(G_111));
    LocalMux I__2245 (
            .O(N__12927),
            .I(G_111));
    LocalMux I__2244 (
            .O(N__12924),
            .I(G_111));
    LocalMux I__2243 (
            .O(N__12921),
            .I(G_111));
    CEMux I__2242 (
            .O(N__12912),
            .I(N__12909));
    LocalMux I__2241 (
            .O(N__12909),
            .I(N__12906));
    Odrv4 I__2240 (
            .O(N__12906),
            .I(\VPP_VDDQ.N_49_1 ));
    CascadeMux I__2239 (
            .O(N__12903),
            .I(\PCH_PWRGD.N_3_i_cascade_ ));
    CascadeMux I__2238 (
            .O(N__12900),
            .I(\PCH_PWRGD.un1_curr_state_0_sqmuxa_0_cascade_ ));
    InMux I__2237 (
            .O(N__12897),
            .I(N__12891));
    InMux I__2236 (
            .O(N__12896),
            .I(N__12891));
    LocalMux I__2235 (
            .O(N__12891),
            .I(N__12888));
    Span4Mux_h I__2234 (
            .O(N__12888),
            .I(N__12885));
    Span4Mux_v I__2233 (
            .O(N__12885),
            .I(N__12882));
    Span4Mux_v I__2232 (
            .O(N__12882),
            .I(N__12879));
    Odrv4 I__2231 (
            .O(N__12879),
            .I(vr_ready_vccin));
    CascadeMux I__2230 (
            .O(N__12876),
            .I(N__12872));
    InMux I__2229 (
            .O(N__12875),
            .I(N__12869));
    InMux I__2228 (
            .O(N__12872),
            .I(N__12866));
    LocalMux I__2227 (
            .O(N__12869),
            .I(\POWERLED.dutycycle_RNIO18NZ0Z_9 ));
    LocalMux I__2226 (
            .O(N__12866),
            .I(\POWERLED.dutycycle_RNIO18NZ0Z_9 ));
    CascadeMux I__2225 (
            .O(N__12861),
            .I(N__12858));
    InMux I__2224 (
            .O(N__12858),
            .I(N__12855));
    LocalMux I__2223 (
            .O(N__12855),
            .I(\POWERLED.dutycycle_RNIC8C11Z0Z_15 ));
    InMux I__2222 (
            .O(N__12852),
            .I(N__12849));
    LocalMux I__2221 (
            .O(N__12849),
            .I(N__12846));
    Odrv4 I__2220 (
            .O(N__12846),
            .I(\POWERLED.dutycycle_RNI31MGZ0Z_12 ));
    CascadeMux I__2219 (
            .O(N__12843),
            .I(N__12840));
    InMux I__2218 (
            .O(N__12840),
            .I(N__12837));
    LocalMux I__2217 (
            .O(N__12837),
            .I(N__12834));
    Odrv4 I__2216 (
            .O(N__12834),
            .I(\POWERLED.dutycycle_RNI31MG_0Z0Z_12 ));
    CascadeMux I__2215 (
            .O(N__12831),
            .I(\POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_1_cascade_ ));
    CascadeMux I__2214 (
            .O(N__12828),
            .I(N__12825));
    InMux I__2213 (
            .O(N__12825),
            .I(N__12822));
    LocalMux I__2212 (
            .O(N__12822),
            .I(\POWERLED.dutycycle_RNI75MGZ0Z_15 ));
    InMux I__2211 (
            .O(N__12819),
            .I(N__12815));
    CascadeMux I__2210 (
            .O(N__12818),
            .I(N__12812));
    LocalMux I__2209 (
            .O(N__12815),
            .I(N__12809));
    InMux I__2208 (
            .O(N__12812),
            .I(N__12806));
    Odrv4 I__2207 (
            .O(N__12809),
            .I(\VPP_VDDQ.N_108_i ));
    LocalMux I__2206 (
            .O(N__12806),
            .I(\VPP_VDDQ.N_108_i ));
    CascadeMux I__2205 (
            .O(N__12801),
            .I(\VPP_VDDQ.N_242_cascade_ ));
    CascadeMux I__2204 (
            .O(N__12798),
            .I(N__12794));
    InMux I__2203 (
            .O(N__12797),
            .I(N__12791));
    InMux I__2202 (
            .O(N__12794),
            .I(N__12788));
    LocalMux I__2201 (
            .O(N__12791),
            .I(\POWERLED.dutycycle_fast_RNILMLMZ0Z_6 ));
    LocalMux I__2200 (
            .O(N__12788),
            .I(\POWERLED.dutycycle_fast_RNILMLMZ0Z_6 ));
    CascadeMux I__2199 (
            .O(N__12783),
            .I(N__12780));
    InMux I__2198 (
            .O(N__12780),
            .I(N__12777));
    LocalMux I__2197 (
            .O(N__12777),
            .I(\POWERLED.dutycycle_RNI84C11Z0Z_14 ));
    InMux I__2196 (
            .O(N__12774),
            .I(N__12771));
    LocalMux I__2195 (
            .O(N__12771),
            .I(\POWERLED.dutycycle_RNIQ09G1Z0Z_10 ));
    CascadeMux I__2194 (
            .O(N__12768),
            .I(\POWERLED.un1_dutycycle_1_39_0_cascade_ ));
    CascadeMux I__2193 (
            .O(N__12765),
            .I(N__12762));
    InMux I__2192 (
            .O(N__12762),
            .I(N__12759));
    LocalMux I__2191 (
            .O(N__12759),
            .I(\POWERLED.dutycycle_RNI34C41Z0Z_8 ));
    InMux I__2190 (
            .O(N__12756),
            .I(N__12753));
    LocalMux I__2189 (
            .O(N__12753),
            .I(\POWERLED.dutycycle_RNI73C11Z0Z_15 ));
    InMux I__2188 (
            .O(N__12750),
            .I(N__12747));
    LocalMux I__2187 (
            .O(N__12747),
            .I(\POWERLED.dutycycle_RNIE4FLZ0Z_9 ));
    InMux I__2186 (
            .O(N__12744),
            .I(N__12741));
    LocalMux I__2185 (
            .O(N__12741),
            .I(\POWERLED.dutycycle_RNI2V0PZ0Z_10 ));
    CascadeMux I__2184 (
            .O(N__12738),
            .I(\POWERLED.dutycycle_RNI2V0PZ0Z_10_cascade_ ));
    CascadeMux I__2183 (
            .O(N__12735),
            .I(N__12732));
    InMux I__2182 (
            .O(N__12732),
            .I(N__12729));
    LocalMux I__2181 (
            .O(N__12729),
            .I(\POWERLED.dutycycle_RNI712I1Z0Z_15 ));
    CascadeMux I__2180 (
            .O(N__12726),
            .I(N__12723));
    InMux I__2179 (
            .O(N__12723),
            .I(N__12719));
    InMux I__2178 (
            .O(N__12722),
            .I(N__12716));
    LocalMux I__2177 (
            .O(N__12719),
            .I(N__12713));
    LocalMux I__2176 (
            .O(N__12716),
            .I(\POWERLED.mult1_un68_sum ));
    Odrv4 I__2175 (
            .O(N__12713),
            .I(\POWERLED.mult1_un68_sum ));
    InMux I__2174 (
            .O(N__12708),
            .I(N__12705));
    LocalMux I__2173 (
            .O(N__12705),
            .I(N__12702));
    Odrv4 I__2172 (
            .O(N__12702),
            .I(\POWERLED.mult1_un68_sum_i ));
    InMux I__2171 (
            .O(N__12699),
            .I(N__12696));
    LocalMux I__2170 (
            .O(N__12696),
            .I(\POWERLED.dutycycle_RNI53MGZ0Z_14 ));
    InMux I__2169 (
            .O(N__12693),
            .I(N__12690));
    LocalMux I__2168 (
            .O(N__12690),
            .I(\POWERLED.dutycycle_RNIJNBA1Z0Z_6 ));
    InMux I__2167 (
            .O(N__12687),
            .I(N__12684));
    LocalMux I__2166 (
            .O(N__12684),
            .I(\POWERLED.dutycycle_RNIOQLJZ0Z_4 ));
    CascadeMux I__2165 (
            .O(N__12681),
            .I(\POWERLED.un1_dutycycle_1_34_0_cascade_ ));
    InMux I__2164 (
            .O(N__12678),
            .I(N__12675));
    LocalMux I__2163 (
            .O(N__12675),
            .I(\POWERLED.un1_dutycycle_1_axb_8 ));
    InMux I__2162 (
            .O(N__12672),
            .I(N__12669));
    LocalMux I__2161 (
            .O(N__12669),
            .I(\POWERLED.dutycycle_RNIB1FLZ0Z_8 ));
    InMux I__2160 (
            .O(N__12666),
            .I(N__12663));
    LocalMux I__2159 (
            .O(N__12663),
            .I(N__12659));
    CascadeMux I__2158 (
            .O(N__12662),
            .I(N__12655));
    Span4Mux_h I__2157 (
            .O(N__12659),
            .I(N__12651));
    InMux I__2156 (
            .O(N__12658),
            .I(N__12646));
    InMux I__2155 (
            .O(N__12655),
            .I(N__12646));
    InMux I__2154 (
            .O(N__12654),
            .I(N__12643));
    Odrv4 I__2153 (
            .O(N__12651),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__2152 (
            .O(N__12646),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__2151 (
            .O(N__12643),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    CascadeMux I__2150 (
            .O(N__12636),
            .I(N__12633));
    InMux I__2149 (
            .O(N__12633),
            .I(N__12630));
    LocalMux I__2148 (
            .O(N__12630),
            .I(\POWERLED.mult1_un68_sum_cry_5_s ));
    InMux I__2147 (
            .O(N__12627),
            .I(N__12624));
    LocalMux I__2146 (
            .O(N__12624),
            .I(\POWERLED.mult1_un75_sum_cry_6_s ));
    InMux I__2145 (
            .O(N__12621),
            .I(\POWERLED.mult1_un75_sum_cry_5 ));
    InMux I__2144 (
            .O(N__12618),
            .I(N__12615));
    LocalMux I__2143 (
            .O(N__12615),
            .I(\POWERLED.mult1_un68_sum_cry_6_s ));
    CascadeMux I__2142 (
            .O(N__12612),
            .I(N__12608));
    CascadeMux I__2141 (
            .O(N__12611),
            .I(N__12604));
    InMux I__2140 (
            .O(N__12608),
            .I(N__12597));
    InMux I__2139 (
            .O(N__12607),
            .I(N__12597));
    InMux I__2138 (
            .O(N__12604),
            .I(N__12597));
    LocalMux I__2137 (
            .O(N__12597),
            .I(\POWERLED.mult1_un68_sum_i_0_8 ));
    CascadeMux I__2136 (
            .O(N__12594),
            .I(N__12591));
    InMux I__2135 (
            .O(N__12591),
            .I(N__12588));
    LocalMux I__2134 (
            .O(N__12588),
            .I(\POWERLED.mult1_un82_sum_axb_8 ));
    InMux I__2133 (
            .O(N__12585),
            .I(\POWERLED.mult1_un75_sum_cry_6 ));
    CascadeMux I__2132 (
            .O(N__12582),
            .I(N__12579));
    InMux I__2131 (
            .O(N__12579),
            .I(N__12576));
    LocalMux I__2130 (
            .O(N__12576),
            .I(\POWERLED.mult1_un75_sum_axb_8 ));
    InMux I__2129 (
            .O(N__12573),
            .I(\POWERLED.mult1_un75_sum_cry_7 ));
    InMux I__2128 (
            .O(N__12570),
            .I(N__12567));
    LocalMux I__2127 (
            .O(N__12567),
            .I(N__12563));
    CascadeMux I__2126 (
            .O(N__12566),
            .I(N__12559));
    Span4Mux_h I__2125 (
            .O(N__12563),
            .I(N__12555));
    InMux I__2124 (
            .O(N__12562),
            .I(N__12550));
    InMux I__2123 (
            .O(N__12559),
            .I(N__12550));
    InMux I__2122 (
            .O(N__12558),
            .I(N__12547));
    Odrv4 I__2121 (
            .O(N__12555),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__2120 (
            .O(N__12550),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__2119 (
            .O(N__12547),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    CascadeMux I__2118 (
            .O(N__12540),
            .I(\POWERLED.mult1_un75_sum_s_8_cascade_ ));
    CascadeMux I__2117 (
            .O(N__12537),
            .I(N__12533));
    CascadeMux I__2116 (
            .O(N__12536),
            .I(N__12529));
    InMux I__2115 (
            .O(N__12533),
            .I(N__12522));
    InMux I__2114 (
            .O(N__12532),
            .I(N__12522));
    InMux I__2113 (
            .O(N__12529),
            .I(N__12522));
    LocalMux I__2112 (
            .O(N__12522),
            .I(\POWERLED.mult1_un75_sum_i_0_8 ));
    CascadeMux I__2111 (
            .O(N__12519),
            .I(N__12516));
    InMux I__2110 (
            .O(N__12516),
            .I(N__12513));
    LocalMux I__2109 (
            .O(N__12513),
            .I(\POWERLED.dutycycle_RNIJL1R1Z0Z_6 ));
    CascadeMux I__2108 (
            .O(N__12510),
            .I(\POWERLED.un1_dutycycle_1_19_0_cascade_ ));
    CascadeMux I__2107 (
            .O(N__12507),
            .I(N__12504));
    InMux I__2106 (
            .O(N__12504),
            .I(N__12501));
    LocalMux I__2105 (
            .O(N__12501),
            .I(\POWERLED.dutycycle_RNIEJ021Z0Z_4 ));
    InMux I__2104 (
            .O(N__12498),
            .I(N__12495));
    LocalMux I__2103 (
            .O(N__12495),
            .I(\POWERLED.dutycycle_RNIQAI81Z0Z_4 ));
    CascadeMux I__2102 (
            .O(N__12492),
            .I(N__12489));
    InMux I__2101 (
            .O(N__12489),
            .I(N__12486));
    LocalMux I__2100 (
            .O(N__12486),
            .I(\POWERLED.mult1_un82_sum_cry_5_s ));
    InMux I__2099 (
            .O(N__12483),
            .I(\POWERLED.mult1_un82_sum_cry_4 ));
    InMux I__2098 (
            .O(N__12480),
            .I(N__12477));
    LocalMux I__2097 (
            .O(N__12477),
            .I(\POWERLED.mult1_un82_sum_cry_6_s ));
    InMux I__2096 (
            .O(N__12474),
            .I(\POWERLED.mult1_un82_sum_cry_5 ));
    CascadeMux I__2095 (
            .O(N__12471),
            .I(N__12468));
    InMux I__2094 (
            .O(N__12468),
            .I(N__12465));
    LocalMux I__2093 (
            .O(N__12465),
            .I(\POWERLED.mult1_un89_sum_axb_8 ));
    InMux I__2092 (
            .O(N__12462),
            .I(\POWERLED.mult1_un82_sum_cry_6 ));
    InMux I__2091 (
            .O(N__12459),
            .I(\POWERLED.mult1_un82_sum_cry_7 ));
    InMux I__2090 (
            .O(N__12456),
            .I(N__12453));
    LocalMux I__2089 (
            .O(N__12453),
            .I(N__12449));
    CascadeMux I__2088 (
            .O(N__12452),
            .I(N__12445));
    Span4Mux_h I__2087 (
            .O(N__12449),
            .I(N__12441));
    InMux I__2086 (
            .O(N__12448),
            .I(N__12436));
    InMux I__2085 (
            .O(N__12445),
            .I(N__12436));
    InMux I__2084 (
            .O(N__12444),
            .I(N__12433));
    Odrv4 I__2083 (
            .O(N__12441),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__2082 (
            .O(N__12436),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__2081 (
            .O(N__12433),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    CascadeMux I__2080 (
            .O(N__12426),
            .I(\POWERLED.mult1_un82_sum_s_8_cascade_ ));
    CascadeMux I__2079 (
            .O(N__12423),
            .I(N__12419));
    CascadeMux I__2078 (
            .O(N__12422),
            .I(N__12415));
    InMux I__2077 (
            .O(N__12419),
            .I(N__12408));
    InMux I__2076 (
            .O(N__12418),
            .I(N__12408));
    InMux I__2075 (
            .O(N__12415),
            .I(N__12408));
    LocalMux I__2074 (
            .O(N__12408),
            .I(\POWERLED.mult1_un82_sum_i_0_8 ));
    InMux I__2073 (
            .O(N__12405),
            .I(N__12402));
    LocalMux I__2072 (
            .O(N__12402),
            .I(N__12398));
    InMux I__2071 (
            .O(N__12401),
            .I(N__12395));
    Span4Mux_h I__2070 (
            .O(N__12398),
            .I(N__12392));
    LocalMux I__2069 (
            .O(N__12395),
            .I(N__12389));
    Odrv4 I__2068 (
            .O(N__12392),
            .I(\POWERLED.mult1_un75_sum ));
    Odrv4 I__2067 (
            .O(N__12389),
            .I(\POWERLED.mult1_un75_sum ));
    CascadeMux I__2066 (
            .O(N__12384),
            .I(N__12381));
    InMux I__2065 (
            .O(N__12381),
            .I(N__12378));
    LocalMux I__2064 (
            .O(N__12378),
            .I(\POWERLED.mult1_un75_sum_cry_3_s ));
    InMux I__2063 (
            .O(N__12375),
            .I(\POWERLED.mult1_un75_sum_cry_2 ));
    CascadeMux I__2062 (
            .O(N__12372),
            .I(N__12369));
    InMux I__2061 (
            .O(N__12369),
            .I(N__12366));
    LocalMux I__2060 (
            .O(N__12366),
            .I(\POWERLED.mult1_un68_sum_cry_3_s ));
    InMux I__2059 (
            .O(N__12363),
            .I(N__12360));
    LocalMux I__2058 (
            .O(N__12360),
            .I(\POWERLED.mult1_un75_sum_cry_4_s ));
    InMux I__2057 (
            .O(N__12357),
            .I(\POWERLED.mult1_un75_sum_cry_3 ));
    InMux I__2056 (
            .O(N__12354),
            .I(N__12351));
    LocalMux I__2055 (
            .O(N__12351),
            .I(\POWERLED.mult1_un68_sum_cry_4_s ));
    CascadeMux I__2054 (
            .O(N__12348),
            .I(N__12345));
    InMux I__2053 (
            .O(N__12345),
            .I(N__12342));
    LocalMux I__2052 (
            .O(N__12342),
            .I(\POWERLED.mult1_un75_sum_cry_5_s ));
    InMux I__2051 (
            .O(N__12339),
            .I(\POWERLED.mult1_un75_sum_cry_4 ));
    CascadeMux I__2050 (
            .O(N__12336),
            .I(N__12333));
    InMux I__2049 (
            .O(N__12333),
            .I(N__12330));
    LocalMux I__2048 (
            .O(N__12330),
            .I(\POWERLED.mult1_un89_sum_cry_5_s ));
    InMux I__2047 (
            .O(N__12327),
            .I(\POWERLED.mult1_un89_sum_cry_4 ));
    InMux I__2046 (
            .O(N__12324),
            .I(N__12321));
    LocalMux I__2045 (
            .O(N__12321),
            .I(\POWERLED.mult1_un89_sum_cry_6_s ));
    InMux I__2044 (
            .O(N__12318),
            .I(\POWERLED.mult1_un89_sum_cry_5 ));
    InMux I__2043 (
            .O(N__12315),
            .I(N__12312));
    LocalMux I__2042 (
            .O(N__12312),
            .I(\POWERLED.mult1_un96_sum_axb_8 ));
    InMux I__2041 (
            .O(N__12309),
            .I(\POWERLED.mult1_un89_sum_cry_6 ));
    InMux I__2040 (
            .O(N__12306),
            .I(\POWERLED.mult1_un89_sum_cry_7 ));
    InMux I__2039 (
            .O(N__12303),
            .I(N__12300));
    LocalMux I__2038 (
            .O(N__12300),
            .I(N__12296));
    CascadeMux I__2037 (
            .O(N__12299),
            .I(N__12292));
    Span4Mux_h I__2036 (
            .O(N__12296),
            .I(N__12288));
    InMux I__2035 (
            .O(N__12295),
            .I(N__12283));
    InMux I__2034 (
            .O(N__12292),
            .I(N__12283));
    InMux I__2033 (
            .O(N__12291),
            .I(N__12280));
    Odrv4 I__2032 (
            .O(N__12288),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__2031 (
            .O(N__12283),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__2030 (
            .O(N__12280),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    CascadeMux I__2029 (
            .O(N__12273),
            .I(\POWERLED.mult1_un89_sum_s_8_cascade_ ));
    CascadeMux I__2028 (
            .O(N__12270),
            .I(N__12266));
    CascadeMux I__2027 (
            .O(N__12269),
            .I(N__12262));
    InMux I__2026 (
            .O(N__12266),
            .I(N__12255));
    InMux I__2025 (
            .O(N__12265),
            .I(N__12255));
    InMux I__2024 (
            .O(N__12262),
            .I(N__12255));
    LocalMux I__2023 (
            .O(N__12255),
            .I(\POWERLED.mult1_un89_sum_i_0_8 ));
    InMux I__2022 (
            .O(N__12252),
            .I(N__12249));
    LocalMux I__2021 (
            .O(N__12249),
            .I(N__12246));
    Span4Mux_h I__2020 (
            .O(N__12246),
            .I(N__12243));
    Odrv4 I__2019 (
            .O(N__12243),
            .I(\POWERLED.mult1_un75_sum_i ));
    CascadeMux I__2018 (
            .O(N__12240),
            .I(N__12237));
    InMux I__2017 (
            .O(N__12237),
            .I(N__12234));
    LocalMux I__2016 (
            .O(N__12234),
            .I(\POWERLED.mult1_un82_sum_cry_3_s ));
    InMux I__2015 (
            .O(N__12231),
            .I(\POWERLED.mult1_un82_sum_cry_2 ));
    InMux I__2014 (
            .O(N__12228),
            .I(N__12225));
    LocalMux I__2013 (
            .O(N__12225),
            .I(\POWERLED.mult1_un82_sum_cry_4_s ));
    InMux I__2012 (
            .O(N__12222),
            .I(\POWERLED.mult1_un82_sum_cry_3 ));
    InMux I__2011 (
            .O(N__12219),
            .I(N__12216));
    LocalMux I__2010 (
            .O(N__12216),
            .I(\POWERLED.mult1_un96_sum_cry_4_s ));
    CascadeMux I__2009 (
            .O(N__12213),
            .I(N__12210));
    InMux I__2008 (
            .O(N__12210),
            .I(N__12207));
    LocalMux I__2007 (
            .O(N__12207),
            .I(\POWERLED.mult1_un103_sum_cry_5_s ));
    InMux I__2006 (
            .O(N__12204),
            .I(\POWERLED.mult1_un103_sum_cry_4 ));
    CascadeMux I__2005 (
            .O(N__12201),
            .I(N__12196));
    InMux I__2004 (
            .O(N__12200),
            .I(N__12192));
    InMux I__2003 (
            .O(N__12199),
            .I(N__12187));
    InMux I__2002 (
            .O(N__12196),
            .I(N__12187));
    InMux I__2001 (
            .O(N__12195),
            .I(N__12184));
    LocalMux I__2000 (
            .O(N__12192),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__1999 (
            .O(N__12187),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__1998 (
            .O(N__12184),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    CascadeMux I__1997 (
            .O(N__12177),
            .I(N__12174));
    InMux I__1996 (
            .O(N__12174),
            .I(N__12171));
    LocalMux I__1995 (
            .O(N__12171),
            .I(\POWERLED.mult1_un96_sum_cry_5_s ));
    InMux I__1994 (
            .O(N__12168),
            .I(N__12165));
    LocalMux I__1993 (
            .O(N__12165),
            .I(\POWERLED.mult1_un103_sum_cry_6_s ));
    InMux I__1992 (
            .O(N__12162),
            .I(\POWERLED.mult1_un103_sum_cry_5 ));
    InMux I__1991 (
            .O(N__12159),
            .I(N__12156));
    LocalMux I__1990 (
            .O(N__12156),
            .I(\POWERLED.mult1_un96_sum_cry_6_s ));
    CascadeMux I__1989 (
            .O(N__12153),
            .I(N__12149));
    CascadeMux I__1988 (
            .O(N__12152),
            .I(N__12145));
    InMux I__1987 (
            .O(N__12149),
            .I(N__12138));
    InMux I__1986 (
            .O(N__12148),
            .I(N__12138));
    InMux I__1985 (
            .O(N__12145),
            .I(N__12138));
    LocalMux I__1984 (
            .O(N__12138),
            .I(\POWERLED.mult1_un96_sum_i_0_8 ));
    InMux I__1983 (
            .O(N__12135),
            .I(N__12132));
    LocalMux I__1982 (
            .O(N__12132),
            .I(\POWERLED.mult1_un110_sum_axb_8 ));
    InMux I__1981 (
            .O(N__12129),
            .I(\POWERLED.mult1_un103_sum_cry_6 ));
    CascadeMux I__1980 (
            .O(N__12126),
            .I(N__12123));
    InMux I__1979 (
            .O(N__12123),
            .I(N__12120));
    LocalMux I__1978 (
            .O(N__12120),
            .I(\POWERLED.mult1_un103_sum_axb_8 ));
    InMux I__1977 (
            .O(N__12117),
            .I(\POWERLED.mult1_un103_sum_cry_7 ));
    InMux I__1976 (
            .O(N__12114),
            .I(N__12110));
    CascadeMux I__1975 (
            .O(N__12113),
            .I(N__12106));
    LocalMux I__1974 (
            .O(N__12110),
            .I(N__12102));
    InMux I__1973 (
            .O(N__12109),
            .I(N__12097));
    InMux I__1972 (
            .O(N__12106),
            .I(N__12097));
    InMux I__1971 (
            .O(N__12105),
            .I(N__12094));
    Odrv4 I__1970 (
            .O(N__12102),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__1969 (
            .O(N__12097),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__1968 (
            .O(N__12094),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    CascadeMux I__1967 (
            .O(N__12087),
            .I(\POWERLED.mult1_un103_sum_s_8_cascade_ ));
    CascadeMux I__1966 (
            .O(N__12084),
            .I(N__12080));
    CascadeMux I__1965 (
            .O(N__12083),
            .I(N__12076));
    InMux I__1964 (
            .O(N__12080),
            .I(N__12069));
    InMux I__1963 (
            .O(N__12079),
            .I(N__12069));
    InMux I__1962 (
            .O(N__12076),
            .I(N__12069));
    LocalMux I__1961 (
            .O(N__12069),
            .I(\POWERLED.mult1_un103_sum_i_0_8 ));
    CascadeMux I__1960 (
            .O(N__12066),
            .I(N__12063));
    InMux I__1959 (
            .O(N__12063),
            .I(N__12060));
    LocalMux I__1958 (
            .O(N__12060),
            .I(\POWERLED.mult1_un89_sum_cry_3_s ));
    InMux I__1957 (
            .O(N__12057),
            .I(\POWERLED.mult1_un89_sum_cry_2 ));
    InMux I__1956 (
            .O(N__12054),
            .I(N__12051));
    LocalMux I__1955 (
            .O(N__12051),
            .I(\POWERLED.mult1_un89_sum_cry_4_s ));
    InMux I__1954 (
            .O(N__12048),
            .I(\POWERLED.mult1_un89_sum_cry_3 ));
    InMux I__1953 (
            .O(N__12045),
            .I(N__12041));
    InMux I__1952 (
            .O(N__12044),
            .I(N__12036));
    LocalMux I__1951 (
            .O(N__12041),
            .I(N__12033));
    InMux I__1950 (
            .O(N__12040),
            .I(N__12030));
    InMux I__1949 (
            .O(N__12039),
            .I(N__12027));
    LocalMux I__1948 (
            .O(N__12036),
            .I(N__12022));
    Span4Mux_v I__1947 (
            .O(N__12033),
            .I(N__12022));
    LocalMux I__1946 (
            .O(N__12030),
            .I(\POWERLED.countZ0Z_12 ));
    LocalMux I__1945 (
            .O(N__12027),
            .I(\POWERLED.countZ0Z_12 ));
    Odrv4 I__1944 (
            .O(N__12022),
            .I(\POWERLED.countZ0Z_12 ));
    InMux I__1943 (
            .O(N__12015),
            .I(\POWERLED.un1_count_1_cry_11 ));
    InMux I__1942 (
            .O(N__12012),
            .I(N__12008));
    InMux I__1941 (
            .O(N__12011),
            .I(N__12004));
    LocalMux I__1940 (
            .O(N__12008),
            .I(N__12000));
    InMux I__1939 (
            .O(N__12007),
            .I(N__11997));
    LocalMux I__1938 (
            .O(N__12004),
            .I(N__11994));
    InMux I__1937 (
            .O(N__12003),
            .I(N__11991));
    Span4Mux_h I__1936 (
            .O(N__12000),
            .I(N__11988));
    LocalMux I__1935 (
            .O(N__11997),
            .I(\POWERLED.countZ0Z_13 ));
    Odrv4 I__1934 (
            .O(N__11994),
            .I(\POWERLED.countZ0Z_13 ));
    LocalMux I__1933 (
            .O(N__11991),
            .I(\POWERLED.countZ0Z_13 ));
    Odrv4 I__1932 (
            .O(N__11988),
            .I(\POWERLED.countZ0Z_13 ));
    InMux I__1931 (
            .O(N__11979),
            .I(\POWERLED.un1_count_1_cry_12 ));
    InMux I__1930 (
            .O(N__11976),
            .I(N__11973));
    LocalMux I__1929 (
            .O(N__11973),
            .I(N__11969));
    InMux I__1928 (
            .O(N__11972),
            .I(N__11965));
    Span4Mux_s2_h I__1927 (
            .O(N__11969),
            .I(N__11961));
    InMux I__1926 (
            .O(N__11968),
            .I(N__11958));
    LocalMux I__1925 (
            .O(N__11965),
            .I(N__11955));
    InMux I__1924 (
            .O(N__11964),
            .I(N__11952));
    Span4Mux_h I__1923 (
            .O(N__11961),
            .I(N__11949));
    LocalMux I__1922 (
            .O(N__11958),
            .I(\POWERLED.countZ0Z_14 ));
    Odrv4 I__1921 (
            .O(N__11955),
            .I(\POWERLED.countZ0Z_14 ));
    LocalMux I__1920 (
            .O(N__11952),
            .I(\POWERLED.countZ0Z_14 ));
    Odrv4 I__1919 (
            .O(N__11949),
            .I(\POWERLED.countZ0Z_14 ));
    InMux I__1918 (
            .O(N__11940),
            .I(\POWERLED.un1_count_1_cry_13 ));
    InMux I__1917 (
            .O(N__11937),
            .I(bfn_6_5_0_));
    CascadeMux I__1916 (
            .O(N__11934),
            .I(N__11929));
    InMux I__1915 (
            .O(N__11933),
            .I(N__11926));
    InMux I__1914 (
            .O(N__11932),
            .I(N__11922));
    InMux I__1913 (
            .O(N__11929),
            .I(N__11919));
    LocalMux I__1912 (
            .O(N__11926),
            .I(N__11916));
    InMux I__1911 (
            .O(N__11925),
            .I(N__11913));
    LocalMux I__1910 (
            .O(N__11922),
            .I(N__11908));
    LocalMux I__1909 (
            .O(N__11919),
            .I(N__11908));
    Span12Mux_s11_v I__1908 (
            .O(N__11916),
            .I(N__11905));
    LocalMux I__1907 (
            .O(N__11913),
            .I(N__11900));
    Span4Mux_v I__1906 (
            .O(N__11908),
            .I(N__11900));
    Odrv12 I__1905 (
            .O(N__11905),
            .I(\POWERLED.countZ0Z_15 ));
    Odrv4 I__1904 (
            .O(N__11900),
            .I(\POWERLED.countZ0Z_15 ));
    CEMux I__1903 (
            .O(N__11895),
            .I(N__11892));
    LocalMux I__1902 (
            .O(N__11892),
            .I(N__11889));
    Odrv4 I__1901 (
            .O(N__11889),
            .I(\POWERLED.N_49_5 ));
    SRMux I__1900 (
            .O(N__11886),
            .I(N__11882));
    SRMux I__1899 (
            .O(N__11885),
            .I(N__11879));
    LocalMux I__1898 (
            .O(N__11882),
            .I(N__11875));
    LocalMux I__1897 (
            .O(N__11879),
            .I(N__11872));
    SRMux I__1896 (
            .O(N__11878),
            .I(N__11868));
    Span4Mux_v I__1895 (
            .O(N__11875),
            .I(N__11863));
    Span4Mux_h I__1894 (
            .O(N__11872),
            .I(N__11860));
    SRMux I__1893 (
            .O(N__11871),
            .I(N__11857));
    LocalMux I__1892 (
            .O(N__11868),
            .I(N__11854));
    SRMux I__1891 (
            .O(N__11867),
            .I(N__11851));
    InMux I__1890 (
            .O(N__11866),
            .I(N__11848));
    Odrv4 I__1889 (
            .O(N__11863),
            .I(\POWERLED.curr_state_RNI75RB5Z0Z_0 ));
    Odrv4 I__1888 (
            .O(N__11860),
            .I(\POWERLED.curr_state_RNI75RB5Z0Z_0 ));
    LocalMux I__1887 (
            .O(N__11857),
            .I(\POWERLED.curr_state_RNI75RB5Z0Z_0 ));
    Odrv12 I__1886 (
            .O(N__11854),
            .I(\POWERLED.curr_state_RNI75RB5Z0Z_0 ));
    LocalMux I__1885 (
            .O(N__11851),
            .I(\POWERLED.curr_state_RNI75RB5Z0Z_0 ));
    LocalMux I__1884 (
            .O(N__11848),
            .I(\POWERLED.curr_state_RNI75RB5Z0Z_0 ));
    InMux I__1883 (
            .O(N__11835),
            .I(N__11831));
    InMux I__1882 (
            .O(N__11834),
            .I(N__11828));
    LocalMux I__1881 (
            .O(N__11831),
            .I(N__11825));
    LocalMux I__1880 (
            .O(N__11828),
            .I(N__11822));
    Span4Mux_v I__1879 (
            .O(N__11825),
            .I(N__11817));
    Span4Mux_v I__1878 (
            .O(N__11822),
            .I(N__11817));
    Odrv4 I__1877 (
            .O(N__11817),
            .I(\POWERLED.mult1_un103_sum ));
    CascadeMux I__1876 (
            .O(N__11814),
            .I(N__11811));
    InMux I__1875 (
            .O(N__11811),
            .I(N__11808));
    LocalMux I__1874 (
            .O(N__11808),
            .I(\POWERLED.mult1_un103_sum_cry_3_s ));
    InMux I__1873 (
            .O(N__11805),
            .I(\POWERLED.mult1_un103_sum_cry_2 ));
    CascadeMux I__1872 (
            .O(N__11802),
            .I(N__11799));
    InMux I__1871 (
            .O(N__11799),
            .I(N__11796));
    LocalMux I__1870 (
            .O(N__11796),
            .I(\POWERLED.mult1_un96_sum_cry_3_s ));
    InMux I__1869 (
            .O(N__11793),
            .I(N__11790));
    LocalMux I__1868 (
            .O(N__11790),
            .I(\POWERLED.mult1_un103_sum_cry_4_s ));
    InMux I__1867 (
            .O(N__11787),
            .I(\POWERLED.mult1_un103_sum_cry_3 ));
    InMux I__1866 (
            .O(N__11784),
            .I(N__11780));
    InMux I__1865 (
            .O(N__11783),
            .I(N__11777));
    LocalMux I__1864 (
            .O(N__11780),
            .I(N__11773));
    LocalMux I__1863 (
            .O(N__11777),
            .I(N__11770));
    InMux I__1862 (
            .O(N__11776),
            .I(N__11766));
    Span4Mux_h I__1861 (
            .O(N__11773),
            .I(N__11763));
    Span4Mux_v I__1860 (
            .O(N__11770),
            .I(N__11760));
    InMux I__1859 (
            .O(N__11769),
            .I(N__11757));
    LocalMux I__1858 (
            .O(N__11766),
            .I(\POWERLED.countZ0Z_4 ));
    Odrv4 I__1857 (
            .O(N__11763),
            .I(\POWERLED.countZ0Z_4 ));
    Odrv4 I__1856 (
            .O(N__11760),
            .I(\POWERLED.countZ0Z_4 ));
    LocalMux I__1855 (
            .O(N__11757),
            .I(\POWERLED.countZ0Z_4 ));
    InMux I__1854 (
            .O(N__11748),
            .I(\POWERLED.un1_count_1_cry_3 ));
    InMux I__1853 (
            .O(N__11745),
            .I(N__11741));
    InMux I__1852 (
            .O(N__11744),
            .I(N__11738));
    LocalMux I__1851 (
            .O(N__11741),
            .I(N__11734));
    LocalMux I__1850 (
            .O(N__11738),
            .I(N__11730));
    InMux I__1849 (
            .O(N__11737),
            .I(N__11727));
    Span4Mux_v I__1848 (
            .O(N__11734),
            .I(N__11724));
    InMux I__1847 (
            .O(N__11733),
            .I(N__11721));
    Span4Mux_h I__1846 (
            .O(N__11730),
            .I(N__11718));
    LocalMux I__1845 (
            .O(N__11727),
            .I(\POWERLED.countZ0Z_5 ));
    Odrv4 I__1844 (
            .O(N__11724),
            .I(\POWERLED.countZ0Z_5 ));
    LocalMux I__1843 (
            .O(N__11721),
            .I(\POWERLED.countZ0Z_5 ));
    Odrv4 I__1842 (
            .O(N__11718),
            .I(\POWERLED.countZ0Z_5 ));
    InMux I__1841 (
            .O(N__11709),
            .I(\POWERLED.un1_count_1_cry_4 ));
    InMux I__1840 (
            .O(N__11706),
            .I(N__11702));
    InMux I__1839 (
            .O(N__11705),
            .I(N__11699));
    LocalMux I__1838 (
            .O(N__11702),
            .I(N__11696));
    LocalMux I__1837 (
            .O(N__11699),
            .I(N__11691));
    Span4Mux_s2_h I__1836 (
            .O(N__11696),
            .I(N__11688));
    InMux I__1835 (
            .O(N__11695),
            .I(N__11685));
    InMux I__1834 (
            .O(N__11694),
            .I(N__11682));
    Span4Mux_v I__1833 (
            .O(N__11691),
            .I(N__11679));
    Span4Mux_h I__1832 (
            .O(N__11688),
            .I(N__11676));
    LocalMux I__1831 (
            .O(N__11685),
            .I(\POWERLED.countZ0Z_6 ));
    LocalMux I__1830 (
            .O(N__11682),
            .I(\POWERLED.countZ0Z_6 ));
    Odrv4 I__1829 (
            .O(N__11679),
            .I(\POWERLED.countZ0Z_6 ));
    Odrv4 I__1828 (
            .O(N__11676),
            .I(\POWERLED.countZ0Z_6 ));
    InMux I__1827 (
            .O(N__11667),
            .I(\POWERLED.un1_count_1_cry_5 ));
    InMux I__1826 (
            .O(N__11664),
            .I(N__11660));
    InMux I__1825 (
            .O(N__11663),
            .I(N__11657));
    LocalMux I__1824 (
            .O(N__11660),
            .I(N__11653));
    LocalMux I__1823 (
            .O(N__11657),
            .I(N__11650));
    InMux I__1822 (
            .O(N__11656),
            .I(N__11646));
    Span4Mux_h I__1821 (
            .O(N__11653),
            .I(N__11643));
    Span4Mux_h I__1820 (
            .O(N__11650),
            .I(N__11640));
    InMux I__1819 (
            .O(N__11649),
            .I(N__11637));
    LocalMux I__1818 (
            .O(N__11646),
            .I(\POWERLED.countZ0Z_7 ));
    Odrv4 I__1817 (
            .O(N__11643),
            .I(\POWERLED.countZ0Z_7 ));
    Odrv4 I__1816 (
            .O(N__11640),
            .I(\POWERLED.countZ0Z_7 ));
    LocalMux I__1815 (
            .O(N__11637),
            .I(\POWERLED.countZ0Z_7 ));
    InMux I__1814 (
            .O(N__11628),
            .I(\POWERLED.un1_count_1_cry_6 ));
    InMux I__1813 (
            .O(N__11625),
            .I(N__11621));
    InMux I__1812 (
            .O(N__11624),
            .I(N__11618));
    LocalMux I__1811 (
            .O(N__11621),
            .I(N__11614));
    LocalMux I__1810 (
            .O(N__11618),
            .I(N__11611));
    InMux I__1809 (
            .O(N__11617),
            .I(N__11607));
    Span4Mux_h I__1808 (
            .O(N__11614),
            .I(N__11604));
    Span4Mux_h I__1807 (
            .O(N__11611),
            .I(N__11601));
    InMux I__1806 (
            .O(N__11610),
            .I(N__11598));
    LocalMux I__1805 (
            .O(N__11607),
            .I(\POWERLED.countZ0Z_8 ));
    Odrv4 I__1804 (
            .O(N__11604),
            .I(\POWERLED.countZ0Z_8 ));
    Odrv4 I__1803 (
            .O(N__11601),
            .I(\POWERLED.countZ0Z_8 ));
    LocalMux I__1802 (
            .O(N__11598),
            .I(\POWERLED.countZ0Z_8 ));
    InMux I__1801 (
            .O(N__11589),
            .I(\POWERLED.un1_count_1_cry_7 ));
    InMux I__1800 (
            .O(N__11586),
            .I(N__11582));
    InMux I__1799 (
            .O(N__11585),
            .I(N__11578));
    LocalMux I__1798 (
            .O(N__11582),
            .I(N__11575));
    InMux I__1797 (
            .O(N__11581),
            .I(N__11571));
    LocalMux I__1796 (
            .O(N__11578),
            .I(N__11568));
    Span4Mux_h I__1795 (
            .O(N__11575),
            .I(N__11565));
    InMux I__1794 (
            .O(N__11574),
            .I(N__11562));
    LocalMux I__1793 (
            .O(N__11571),
            .I(\POWERLED.countZ0Z_9 ));
    Odrv4 I__1792 (
            .O(N__11568),
            .I(\POWERLED.countZ0Z_9 ));
    Odrv4 I__1791 (
            .O(N__11565),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__1790 (
            .O(N__11562),
            .I(\POWERLED.countZ0Z_9 ));
    InMux I__1789 (
            .O(N__11553),
            .I(bfn_6_4_0_));
    InMux I__1788 (
            .O(N__11550),
            .I(N__11547));
    LocalMux I__1787 (
            .O(N__11547),
            .I(N__11543));
    InMux I__1786 (
            .O(N__11546),
            .I(N__11538));
    Span4Mux_s2_h I__1785 (
            .O(N__11543),
            .I(N__11535));
    CascadeMux I__1784 (
            .O(N__11542),
            .I(N__11532));
    InMux I__1783 (
            .O(N__11541),
            .I(N__11529));
    LocalMux I__1782 (
            .O(N__11538),
            .I(N__11526));
    Span4Mux_h I__1781 (
            .O(N__11535),
            .I(N__11523));
    InMux I__1780 (
            .O(N__11532),
            .I(N__11520));
    LocalMux I__1779 (
            .O(N__11529),
            .I(\POWERLED.countZ0Z_10 ));
    Odrv4 I__1778 (
            .O(N__11526),
            .I(\POWERLED.countZ0Z_10 ));
    Odrv4 I__1777 (
            .O(N__11523),
            .I(\POWERLED.countZ0Z_10 ));
    LocalMux I__1776 (
            .O(N__11520),
            .I(\POWERLED.countZ0Z_10 ));
    InMux I__1775 (
            .O(N__11511),
            .I(\POWERLED.un1_count_1_cry_9 ));
    InMux I__1774 (
            .O(N__11508),
            .I(N__11504));
    InMux I__1773 (
            .O(N__11507),
            .I(N__11499));
    LocalMux I__1772 (
            .O(N__11504),
            .I(N__11496));
    InMux I__1771 (
            .O(N__11503),
            .I(N__11493));
    InMux I__1770 (
            .O(N__11502),
            .I(N__11490));
    LocalMux I__1769 (
            .O(N__11499),
            .I(N__11485));
    Span4Mux_v I__1768 (
            .O(N__11496),
            .I(N__11485));
    LocalMux I__1767 (
            .O(N__11493),
            .I(\POWERLED.countZ0Z_11 ));
    LocalMux I__1766 (
            .O(N__11490),
            .I(\POWERLED.countZ0Z_11 ));
    Odrv4 I__1765 (
            .O(N__11485),
            .I(\POWERLED.countZ0Z_11 ));
    InMux I__1764 (
            .O(N__11478),
            .I(\POWERLED.un1_count_1_cry_10 ));
    InMux I__1763 (
            .O(N__11475),
            .I(N__11471));
    InMux I__1762 (
            .O(N__11474),
            .I(N__11468));
    LocalMux I__1761 (
            .O(N__11471),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    LocalMux I__1760 (
            .O(N__11468),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    InMux I__1759 (
            .O(N__11463),
            .I(\VPP_VDDQ.un1_count_1_cry_11 ));
    InMux I__1758 (
            .O(N__11460),
            .I(N__11456));
    InMux I__1757 (
            .O(N__11459),
            .I(N__11453));
    LocalMux I__1756 (
            .O(N__11456),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    LocalMux I__1755 (
            .O(N__11453),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    InMux I__1754 (
            .O(N__11448),
            .I(\VPP_VDDQ.un1_count_1_cry_12 ));
    InMux I__1753 (
            .O(N__11445),
            .I(N__11441));
    InMux I__1752 (
            .O(N__11444),
            .I(N__11438));
    LocalMux I__1751 (
            .O(N__11441),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    LocalMux I__1750 (
            .O(N__11438),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    InMux I__1749 (
            .O(N__11433),
            .I(\VPP_VDDQ.un1_count_1_cry_13 ));
    InMux I__1748 (
            .O(N__11430),
            .I(bfn_5_15_0_));
    CascadeMux I__1747 (
            .O(N__11427),
            .I(N__11423));
    InMux I__1746 (
            .O(N__11426),
            .I(N__11420));
    InMux I__1745 (
            .O(N__11423),
            .I(N__11417));
    LocalMux I__1744 (
            .O(N__11420),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    LocalMux I__1743 (
            .O(N__11417),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    InMux I__1742 (
            .O(N__11412),
            .I(N__11409));
    LocalMux I__1741 (
            .O(N__11409),
            .I(N__11406));
    Span4Mux_v I__1740 (
            .O(N__11406),
            .I(N__11401));
    InMux I__1739 (
            .O(N__11405),
            .I(N__11398));
    InMux I__1738 (
            .O(N__11404),
            .I(N__11395));
    Span4Mux_h I__1737 (
            .O(N__11401),
            .I(N__11392));
    LocalMux I__1736 (
            .O(N__11398),
            .I(\POWERLED.countZ0Z_1 ));
    LocalMux I__1735 (
            .O(N__11395),
            .I(\POWERLED.countZ0Z_1 ));
    Odrv4 I__1734 (
            .O(N__11392),
            .I(\POWERLED.countZ0Z_1 ));
    CascadeMux I__1733 (
            .O(N__11385),
            .I(N__11379));
    InMux I__1732 (
            .O(N__11384),
            .I(N__11376));
    InMux I__1731 (
            .O(N__11383),
            .I(N__11373));
    InMux I__1730 (
            .O(N__11382),
            .I(N__11370));
    InMux I__1729 (
            .O(N__11379),
            .I(N__11367));
    LocalMux I__1728 (
            .O(N__11376),
            .I(N__11364));
    LocalMux I__1727 (
            .O(N__11373),
            .I(N__11357));
    LocalMux I__1726 (
            .O(N__11370),
            .I(N__11357));
    LocalMux I__1725 (
            .O(N__11367),
            .I(N__11357));
    Span4Mux_s3_h I__1724 (
            .O(N__11364),
            .I(N__11354));
    Odrv4 I__1723 (
            .O(N__11357),
            .I(\POWERLED.countZ0Z_0 ));
    Odrv4 I__1722 (
            .O(N__11354),
            .I(\POWERLED.countZ0Z_0 ));
    InMux I__1721 (
            .O(N__11349),
            .I(N__11345));
    InMux I__1720 (
            .O(N__11348),
            .I(N__11342));
    LocalMux I__1719 (
            .O(N__11345),
            .I(N__11338));
    LocalMux I__1718 (
            .O(N__11342),
            .I(N__11335));
    InMux I__1717 (
            .O(N__11341),
            .I(N__11331));
    Span4Mux_h I__1716 (
            .O(N__11338),
            .I(N__11328));
    Span4Mux_h I__1715 (
            .O(N__11335),
            .I(N__11325));
    InMux I__1714 (
            .O(N__11334),
            .I(N__11322));
    LocalMux I__1713 (
            .O(N__11331),
            .I(\POWERLED.countZ0Z_2 ));
    Odrv4 I__1712 (
            .O(N__11328),
            .I(\POWERLED.countZ0Z_2 ));
    Odrv4 I__1711 (
            .O(N__11325),
            .I(\POWERLED.countZ0Z_2 ));
    LocalMux I__1710 (
            .O(N__11322),
            .I(\POWERLED.countZ0Z_2 ));
    InMux I__1709 (
            .O(N__11313),
            .I(\POWERLED.un1_count_1_cry_1 ));
    InMux I__1708 (
            .O(N__11310),
            .I(N__11306));
    InMux I__1707 (
            .O(N__11309),
            .I(N__11303));
    LocalMux I__1706 (
            .O(N__11306),
            .I(N__11299));
    LocalMux I__1705 (
            .O(N__11303),
            .I(N__11296));
    InMux I__1704 (
            .O(N__11302),
            .I(N__11292));
    Span4Mux_h I__1703 (
            .O(N__11299),
            .I(N__11289));
    Span4Mux_v I__1702 (
            .O(N__11296),
            .I(N__11286));
    InMux I__1701 (
            .O(N__11295),
            .I(N__11283));
    LocalMux I__1700 (
            .O(N__11292),
            .I(\POWERLED.countZ0Z_3 ));
    Odrv4 I__1699 (
            .O(N__11289),
            .I(\POWERLED.countZ0Z_3 ));
    Odrv4 I__1698 (
            .O(N__11286),
            .I(\POWERLED.countZ0Z_3 ));
    LocalMux I__1697 (
            .O(N__11283),
            .I(\POWERLED.countZ0Z_3 ));
    InMux I__1696 (
            .O(N__11274),
            .I(\POWERLED.un1_count_1_cry_2 ));
    InMux I__1695 (
            .O(N__11271),
            .I(N__11267));
    InMux I__1694 (
            .O(N__11270),
            .I(N__11264));
    LocalMux I__1693 (
            .O(N__11267),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    LocalMux I__1692 (
            .O(N__11264),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    InMux I__1691 (
            .O(N__11259),
            .I(\VPP_VDDQ.un1_count_1_cry_2 ));
    InMux I__1690 (
            .O(N__11256),
            .I(N__11252));
    InMux I__1689 (
            .O(N__11255),
            .I(N__11249));
    LocalMux I__1688 (
            .O(N__11252),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    LocalMux I__1687 (
            .O(N__11249),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    InMux I__1686 (
            .O(N__11244),
            .I(\VPP_VDDQ.un1_count_1_cry_3 ));
    InMux I__1685 (
            .O(N__11241),
            .I(N__11237));
    InMux I__1684 (
            .O(N__11240),
            .I(N__11234));
    LocalMux I__1683 (
            .O(N__11237),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    LocalMux I__1682 (
            .O(N__11234),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    InMux I__1681 (
            .O(N__11229),
            .I(\VPP_VDDQ.un1_count_1_cry_4 ));
    InMux I__1680 (
            .O(N__11226),
            .I(N__11222));
    InMux I__1679 (
            .O(N__11225),
            .I(N__11219));
    LocalMux I__1678 (
            .O(N__11222),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    LocalMux I__1677 (
            .O(N__11219),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    InMux I__1676 (
            .O(N__11214),
            .I(\VPP_VDDQ.un1_count_1_cry_5 ));
    CascadeMux I__1675 (
            .O(N__11211),
            .I(N__11207));
    InMux I__1674 (
            .O(N__11210),
            .I(N__11204));
    InMux I__1673 (
            .O(N__11207),
            .I(N__11201));
    LocalMux I__1672 (
            .O(N__11204),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    LocalMux I__1671 (
            .O(N__11201),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    InMux I__1670 (
            .O(N__11196),
            .I(\VPP_VDDQ.un1_count_1_cry_6 ));
    InMux I__1669 (
            .O(N__11193),
            .I(N__11189));
    InMux I__1668 (
            .O(N__11192),
            .I(N__11186));
    LocalMux I__1667 (
            .O(N__11189),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    LocalMux I__1666 (
            .O(N__11186),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    InMux I__1665 (
            .O(N__11181),
            .I(bfn_5_14_0_));
    InMux I__1664 (
            .O(N__11178),
            .I(N__11174));
    InMux I__1663 (
            .O(N__11177),
            .I(N__11171));
    LocalMux I__1662 (
            .O(N__11174),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    LocalMux I__1661 (
            .O(N__11171),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    InMux I__1660 (
            .O(N__11166),
            .I(\VPP_VDDQ.un1_count_1_cry_8 ));
    CascadeMux I__1659 (
            .O(N__11163),
            .I(N__11159));
    InMux I__1658 (
            .O(N__11162),
            .I(N__11156));
    InMux I__1657 (
            .O(N__11159),
            .I(N__11153));
    LocalMux I__1656 (
            .O(N__11156),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    LocalMux I__1655 (
            .O(N__11153),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    InMux I__1654 (
            .O(N__11148),
            .I(\VPP_VDDQ.un1_count_1_cry_9 ));
    CascadeMux I__1653 (
            .O(N__11145),
            .I(N__11141));
    InMux I__1652 (
            .O(N__11144),
            .I(N__11138));
    InMux I__1651 (
            .O(N__11141),
            .I(N__11135));
    LocalMux I__1650 (
            .O(N__11138),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    LocalMux I__1649 (
            .O(N__11135),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    InMux I__1648 (
            .O(N__11130),
            .I(\VPP_VDDQ.un1_count_1_cry_10 ));
    InMux I__1647 (
            .O(N__11127),
            .I(bfn_5_12_0_));
    InMux I__1646 (
            .O(N__11124),
            .I(\POWERLED.CO2 ));
    InMux I__1645 (
            .O(N__11121),
            .I(N__11118));
    LocalMux I__1644 (
            .O(N__11118),
            .I(\POWERLED.CO2_THRU_CO ));
    CascadeMux I__1643 (
            .O(N__11115),
            .I(N__11112));
    InMux I__1642 (
            .O(N__11112),
            .I(N__11106));
    InMux I__1641 (
            .O(N__11111),
            .I(N__11103));
    InMux I__1640 (
            .O(N__11110),
            .I(N__11098));
    InMux I__1639 (
            .O(N__11109),
            .I(N__11098));
    LocalMux I__1638 (
            .O(N__11106),
            .I(\POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1 ));
    LocalMux I__1637 (
            .O(N__11103),
            .I(\POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1 ));
    LocalMux I__1636 (
            .O(N__11098),
            .I(\POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1 ));
    CascadeMux I__1635 (
            .O(N__11091),
            .I(\POWERLED.CO2_THRU_CO_cascade_ ));
    CascadeMux I__1634 (
            .O(N__11088),
            .I(N__11085));
    InMux I__1633 (
            .O(N__11085),
            .I(N__11080));
    InMux I__1632 (
            .O(N__11084),
            .I(N__11077));
    InMux I__1631 (
            .O(N__11083),
            .I(N__11074));
    LocalMux I__1630 (
            .O(N__11080),
            .I(N__11071));
    LocalMux I__1629 (
            .O(N__11077),
            .I(\POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71 ));
    LocalMux I__1628 (
            .O(N__11074),
            .I(\POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71 ));
    Odrv4 I__1627 (
            .O(N__11071),
            .I(\POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71 ));
    InMux I__1626 (
            .O(N__11064),
            .I(N__11061));
    LocalMux I__1625 (
            .O(N__11061),
            .I(N__11058));
    Odrv4 I__1624 (
            .O(N__11058),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_4 ));
    InMux I__1623 (
            .O(N__11055),
            .I(N__11051));
    InMux I__1622 (
            .O(N__11054),
            .I(N__11048));
    LocalMux I__1621 (
            .O(N__11051),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    LocalMux I__1620 (
            .O(N__11048),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    InMux I__1619 (
            .O(N__11043),
            .I(N__11039));
    InMux I__1618 (
            .O(N__11042),
            .I(N__11036));
    LocalMux I__1617 (
            .O(N__11039),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    LocalMux I__1616 (
            .O(N__11036),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    InMux I__1615 (
            .O(N__11031),
            .I(\VPP_VDDQ.un1_count_1_cry_0 ));
    InMux I__1614 (
            .O(N__11028),
            .I(N__11024));
    InMux I__1613 (
            .O(N__11027),
            .I(N__11021));
    LocalMux I__1612 (
            .O(N__11024),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    LocalMux I__1611 (
            .O(N__11021),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    InMux I__1610 (
            .O(N__11016),
            .I(\VPP_VDDQ.un1_count_1_cry_1 ));
    InMux I__1609 (
            .O(N__11013),
            .I(\POWERLED.un1_dutycycle_1_cry_6 ));
    InMux I__1608 (
            .O(N__11010),
            .I(bfn_5_11_0_));
    InMux I__1607 (
            .O(N__11007),
            .I(\POWERLED.un1_dutycycle_1_cry_8 ));
    InMux I__1606 (
            .O(N__11004),
            .I(\POWERLED.un1_dutycycle_1_cry_9 ));
    InMux I__1605 (
            .O(N__11001),
            .I(\POWERLED.un1_dutycycle_1_cry_10 ));
    CascadeMux I__1604 (
            .O(N__10998),
            .I(N__10995));
    InMux I__1603 (
            .O(N__10995),
            .I(N__10991));
    InMux I__1602 (
            .O(N__10994),
            .I(N__10988));
    LocalMux I__1601 (
            .O(N__10991),
            .I(N__10985));
    LocalMux I__1600 (
            .O(N__10988),
            .I(\POWERLED.mult1_un61_sum ));
    Odrv4 I__1599 (
            .O(N__10985),
            .I(\POWERLED.mult1_un61_sum ));
    InMux I__1598 (
            .O(N__10980),
            .I(\POWERLED.un1_dutycycle_1_cry_11 ));
    CascadeMux I__1597 (
            .O(N__10977),
            .I(N__10973));
    InMux I__1596 (
            .O(N__10976),
            .I(N__10970));
    InMux I__1595 (
            .O(N__10973),
            .I(N__10967));
    LocalMux I__1594 (
            .O(N__10970),
            .I(N__10962));
    LocalMux I__1593 (
            .O(N__10967),
            .I(N__10962));
    Odrv4 I__1592 (
            .O(N__10962),
            .I(\POWERLED.mult1_un54_sum ));
    InMux I__1591 (
            .O(N__10959),
            .I(\POWERLED.un1_dutycycle_1_cry_12 ));
    CascadeMux I__1590 (
            .O(N__10956),
            .I(N__10953));
    InMux I__1589 (
            .O(N__10953),
            .I(N__10949));
    InMux I__1588 (
            .O(N__10952),
            .I(N__10946));
    LocalMux I__1587 (
            .O(N__10949),
            .I(N__10943));
    LocalMux I__1586 (
            .O(N__10946),
            .I(\POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1 ));
    Odrv4 I__1585 (
            .O(N__10943),
            .I(\POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1 ));
    InMux I__1584 (
            .O(N__10938),
            .I(\POWERLED.un1_dutycycle_1_cry_13 ));
    InMux I__1583 (
            .O(N__10935),
            .I(\POWERLED.un1_dutycycle_1_cry_14 ));
    CascadeMux I__1582 (
            .O(N__10932),
            .I(N__10929));
    InMux I__1581 (
            .O(N__10929),
            .I(N__10926));
    LocalMux I__1580 (
            .O(N__10926),
            .I(\POWERLED.mult1_un68_sum_axb_8 ));
    InMux I__1579 (
            .O(N__10923),
            .I(\POWERLED.mult1_un68_sum_cry_7 ));
    CascadeMux I__1578 (
            .O(N__10920),
            .I(\POWERLED.mult1_un68_sum_s_8_cascade_ ));
    CascadeMux I__1577 (
            .O(N__10917),
            .I(N__10913));
    InMux I__1576 (
            .O(N__10916),
            .I(N__10910));
    InMux I__1575 (
            .O(N__10913),
            .I(N__10907));
    LocalMux I__1574 (
            .O(N__10910),
            .I(N__10902));
    LocalMux I__1573 (
            .O(N__10907),
            .I(N__10902));
    Span12Mux_s9_v I__1572 (
            .O(N__10902),
            .I(N__10899));
    Odrv12 I__1571 (
            .O(N__10899),
            .I(\POWERLED.un1_dutycycle_1_axb_0 ));
    InMux I__1570 (
            .O(N__10896),
            .I(N__10892));
    InMux I__1569 (
            .O(N__10895),
            .I(N__10889));
    LocalMux I__1568 (
            .O(N__10892),
            .I(N__10886));
    LocalMux I__1567 (
            .O(N__10889),
            .I(N__10883));
    Span4Mux_h I__1566 (
            .O(N__10886),
            .I(N__10880));
    Span4Mux_h I__1565 (
            .O(N__10883),
            .I(N__10875));
    Span4Mux_v I__1564 (
            .O(N__10880),
            .I(N__10875));
    Odrv4 I__1563 (
            .O(N__10875),
            .I(\POWERLED.mult1_un138_sum ));
    InMux I__1562 (
            .O(N__10872),
            .I(\POWERLED.un1_dutycycle_1_cry_0 ));
    InMux I__1561 (
            .O(N__10869),
            .I(N__10865));
    InMux I__1560 (
            .O(N__10868),
            .I(N__10862));
    LocalMux I__1559 (
            .O(N__10865),
            .I(N__10859));
    LocalMux I__1558 (
            .O(N__10862),
            .I(N__10856));
    Span4Mux_h I__1557 (
            .O(N__10859),
            .I(N__10853));
    Span4Mux_h I__1556 (
            .O(N__10856),
            .I(N__10850));
    Span4Mux_v I__1555 (
            .O(N__10853),
            .I(N__10847));
    Span4Mux_v I__1554 (
            .O(N__10850),
            .I(N__10844));
    Odrv4 I__1553 (
            .O(N__10847),
            .I(\POWERLED.mult1_un131_sum ));
    Odrv4 I__1552 (
            .O(N__10844),
            .I(\POWERLED.mult1_un131_sum ));
    InMux I__1551 (
            .O(N__10839),
            .I(\POWERLED.un1_dutycycle_1_cry_1 ));
    InMux I__1550 (
            .O(N__10836),
            .I(N__10832));
    InMux I__1549 (
            .O(N__10835),
            .I(N__10829));
    LocalMux I__1548 (
            .O(N__10832),
            .I(N__10826));
    LocalMux I__1547 (
            .O(N__10829),
            .I(N__10823));
    Span4Mux_h I__1546 (
            .O(N__10826),
            .I(N__10820));
    Span4Mux_h I__1545 (
            .O(N__10823),
            .I(N__10817));
    Span4Mux_v I__1544 (
            .O(N__10820),
            .I(N__10814));
    Span4Mux_v I__1543 (
            .O(N__10817),
            .I(N__10811));
    Odrv4 I__1542 (
            .O(N__10814),
            .I(\POWERLED.mult1_un124_sum ));
    Odrv4 I__1541 (
            .O(N__10811),
            .I(\POWERLED.mult1_un124_sum ));
    InMux I__1540 (
            .O(N__10806),
            .I(\POWERLED.un1_dutycycle_1_cry_2 ));
    InMux I__1539 (
            .O(N__10803),
            .I(N__10799));
    InMux I__1538 (
            .O(N__10802),
            .I(N__10796));
    LocalMux I__1537 (
            .O(N__10799),
            .I(N__10793));
    LocalMux I__1536 (
            .O(N__10796),
            .I(N__10790));
    Span4Mux_v I__1535 (
            .O(N__10793),
            .I(N__10787));
    Span4Mux_v I__1534 (
            .O(N__10790),
            .I(N__10784));
    Span4Mux_v I__1533 (
            .O(N__10787),
            .I(N__10781));
    Span4Mux_h I__1532 (
            .O(N__10784),
            .I(N__10778));
    Odrv4 I__1531 (
            .O(N__10781),
            .I(\POWERLED.mult1_un117_sum ));
    Odrv4 I__1530 (
            .O(N__10778),
            .I(\POWERLED.mult1_un117_sum ));
    InMux I__1529 (
            .O(N__10773),
            .I(\POWERLED.un1_dutycycle_1_cry_3 ));
    InMux I__1528 (
            .O(N__10770),
            .I(N__10766));
    InMux I__1527 (
            .O(N__10769),
            .I(N__10763));
    LocalMux I__1526 (
            .O(N__10766),
            .I(N__10758));
    LocalMux I__1525 (
            .O(N__10763),
            .I(N__10758));
    Odrv12 I__1524 (
            .O(N__10758),
            .I(\POWERLED.mult1_un110_sum ));
    InMux I__1523 (
            .O(N__10755),
            .I(\POWERLED.un1_dutycycle_1_cry_4 ));
    InMux I__1522 (
            .O(N__10752),
            .I(\POWERLED.un1_dutycycle_1_cry_5 ));
    CascadeMux I__1521 (
            .O(N__10749),
            .I(N__10745));
    InMux I__1520 (
            .O(N__10748),
            .I(N__10742));
    InMux I__1519 (
            .O(N__10745),
            .I(N__10739));
    LocalMux I__1518 (
            .O(N__10742),
            .I(\POWERLED.mult1_un47_sum_cry_6_s ));
    LocalMux I__1517 (
            .O(N__10739),
            .I(\POWERLED.mult1_un47_sum_cry_6_s ));
    CascadeMux I__1516 (
            .O(N__10734),
            .I(N__10729));
    InMux I__1515 (
            .O(N__10733),
            .I(N__10722));
    InMux I__1514 (
            .O(N__10732),
            .I(N__10722));
    InMux I__1513 (
            .O(N__10729),
            .I(N__10722));
    LocalMux I__1512 (
            .O(N__10722),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    CascadeMux I__1511 (
            .O(N__10719),
            .I(N__10716));
    InMux I__1510 (
            .O(N__10716),
            .I(N__10713));
    LocalMux I__1509 (
            .O(N__10713),
            .I(\POWERLED.mult1_un54_sum_cry_6_THRU_CO ));
    InMux I__1508 (
            .O(N__10710),
            .I(\POWERLED.mult1_un61_sum_cry_7 ));
    CascadeMux I__1507 (
            .O(N__10707),
            .I(\POWERLED.mult1_un61_sum_s_8_cascade_ ));
    InMux I__1506 (
            .O(N__10704),
            .I(N__10701));
    LocalMux I__1505 (
            .O(N__10701),
            .I(N__10698));
    Odrv4 I__1504 (
            .O(N__10698),
            .I(\POWERLED.mult1_un61_sum_i ));
    InMux I__1503 (
            .O(N__10695),
            .I(\POWERLED.mult1_un68_sum_cry_2 ));
    CascadeMux I__1502 (
            .O(N__10692),
            .I(N__10689));
    InMux I__1501 (
            .O(N__10689),
            .I(N__10686));
    LocalMux I__1500 (
            .O(N__10686),
            .I(\POWERLED.mult1_un61_sum_cry_3_s ));
    InMux I__1499 (
            .O(N__10683),
            .I(\POWERLED.mult1_un68_sum_cry_3 ));
    InMux I__1498 (
            .O(N__10680),
            .I(N__10677));
    LocalMux I__1497 (
            .O(N__10677),
            .I(\POWERLED.mult1_un61_sum_cry_4_s ));
    InMux I__1496 (
            .O(N__10674),
            .I(\POWERLED.mult1_un68_sum_cry_4 ));
    CascadeMux I__1495 (
            .O(N__10671),
            .I(N__10666));
    InMux I__1494 (
            .O(N__10670),
            .I(N__10662));
    InMux I__1493 (
            .O(N__10669),
            .I(N__10657));
    InMux I__1492 (
            .O(N__10666),
            .I(N__10657));
    InMux I__1491 (
            .O(N__10665),
            .I(N__10654));
    LocalMux I__1490 (
            .O(N__10662),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__1489 (
            .O(N__10657),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__1488 (
            .O(N__10654),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    CascadeMux I__1487 (
            .O(N__10647),
            .I(N__10644));
    InMux I__1486 (
            .O(N__10644),
            .I(N__10641));
    LocalMux I__1485 (
            .O(N__10641),
            .I(\POWERLED.mult1_un61_sum_cry_5_s ));
    InMux I__1484 (
            .O(N__10638),
            .I(\POWERLED.mult1_un68_sum_cry_5 ));
    InMux I__1483 (
            .O(N__10635),
            .I(N__10632));
    LocalMux I__1482 (
            .O(N__10632),
            .I(\POWERLED.mult1_un61_sum_cry_6_s ));
    CascadeMux I__1481 (
            .O(N__10629),
            .I(N__10625));
    CascadeMux I__1480 (
            .O(N__10628),
            .I(N__10621));
    InMux I__1479 (
            .O(N__10625),
            .I(N__10614));
    InMux I__1478 (
            .O(N__10624),
            .I(N__10614));
    InMux I__1477 (
            .O(N__10621),
            .I(N__10614));
    LocalMux I__1476 (
            .O(N__10614),
            .I(\POWERLED.mult1_un61_sum_i_0_8 ));
    InMux I__1475 (
            .O(N__10611),
            .I(\POWERLED.mult1_un68_sum_cry_6 ));
    InMux I__1474 (
            .O(N__10608),
            .I(\POWERLED.mult1_un96_sum_cry_6 ));
    InMux I__1473 (
            .O(N__10605),
            .I(\POWERLED.mult1_un96_sum_cry_7 ));
    CascadeMux I__1472 (
            .O(N__10602),
            .I(\POWERLED.mult1_un96_sum_s_8_cascade_ ));
    InMux I__1471 (
            .O(N__10599),
            .I(N__10596));
    LocalMux I__1470 (
            .O(N__10596),
            .I(\POWERLED.mult1_un54_sum_i ));
    InMux I__1469 (
            .O(N__10593),
            .I(\POWERLED.mult1_un61_sum_cry_2 ));
    CascadeMux I__1468 (
            .O(N__10590),
            .I(N__10587));
    InMux I__1467 (
            .O(N__10587),
            .I(N__10584));
    LocalMux I__1466 (
            .O(N__10584),
            .I(\POWERLED.mult1_un54_sum_cry_3_s ));
    InMux I__1465 (
            .O(N__10581),
            .I(\POWERLED.mult1_un61_sum_cry_3 ));
    InMux I__1464 (
            .O(N__10578),
            .I(N__10575));
    LocalMux I__1463 (
            .O(N__10575),
            .I(\POWERLED.mult1_un54_sum_cry_4_s ));
    InMux I__1462 (
            .O(N__10572),
            .I(\POWERLED.mult1_un61_sum_cry_4 ));
    CascadeMux I__1461 (
            .O(N__10569),
            .I(N__10566));
    InMux I__1460 (
            .O(N__10566),
            .I(N__10563));
    LocalMux I__1459 (
            .O(N__10563),
            .I(\POWERLED.mult1_un54_sum_cry_5_s ));
    InMux I__1458 (
            .O(N__10560),
            .I(\POWERLED.mult1_un61_sum_cry_5 ));
    InMux I__1457 (
            .O(N__10557),
            .I(N__10554));
    LocalMux I__1456 (
            .O(N__10554),
            .I(\POWERLED.mult1_un54_sum_cry_6_s ));
    CascadeMux I__1455 (
            .O(N__10551),
            .I(N__10547));
    CascadeMux I__1454 (
            .O(N__10550),
            .I(N__10543));
    InMux I__1453 (
            .O(N__10547),
            .I(N__10536));
    InMux I__1452 (
            .O(N__10546),
            .I(N__10536));
    InMux I__1451 (
            .O(N__10543),
            .I(N__10536));
    LocalMux I__1450 (
            .O(N__10536),
            .I(\POWERLED.mult1_un54_sum_i_8 ));
    InMux I__1449 (
            .O(N__10533),
            .I(\POWERLED.mult1_un61_sum_cry_6 ));
    InMux I__1448 (
            .O(N__10530),
            .I(N__10527));
    LocalMux I__1447 (
            .O(N__10527),
            .I(\POWERLED.mult1_un110_sum_cry_6_s ));
    InMux I__1446 (
            .O(N__10524),
            .I(\POWERLED.mult1_un110_sum_cry_5 ));
    InMux I__1445 (
            .O(N__10521),
            .I(N__10518));
    LocalMux I__1444 (
            .O(N__10518),
            .I(\POWERLED.mult1_un117_sum_axb_8 ));
    InMux I__1443 (
            .O(N__10515),
            .I(\POWERLED.mult1_un110_sum_cry_6 ));
    InMux I__1442 (
            .O(N__10512),
            .I(\POWERLED.mult1_un110_sum_cry_7 ));
    CascadeMux I__1441 (
            .O(N__10509),
            .I(N__10505));
    InMux I__1440 (
            .O(N__10508),
            .I(N__10497));
    InMux I__1439 (
            .O(N__10505),
            .I(N__10497));
    InMux I__1438 (
            .O(N__10504),
            .I(N__10494));
    InMux I__1437 (
            .O(N__10503),
            .I(N__10489));
    InMux I__1436 (
            .O(N__10502),
            .I(N__10489));
    LocalMux I__1435 (
            .O(N__10497),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__1434 (
            .O(N__10494),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__1433 (
            .O(N__10489),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    InMux I__1432 (
            .O(N__10482),
            .I(N__10479));
    LocalMux I__1431 (
            .O(N__10479),
            .I(\POWERLED.mult1_un103_sum_i ));
    InMux I__1430 (
            .O(N__10476),
            .I(\POWERLED.mult1_un96_sum_cry_2 ));
    InMux I__1429 (
            .O(N__10473),
            .I(\POWERLED.mult1_un96_sum_cry_3 ));
    InMux I__1428 (
            .O(N__10470),
            .I(\POWERLED.mult1_un96_sum_cry_4 ));
    InMux I__1427 (
            .O(N__10467),
            .I(\POWERLED.mult1_un96_sum_cry_5 ));
    CascadeMux I__1426 (
            .O(N__10464),
            .I(\POWERLED.un1_countlt6_cascade_ ));
    InMux I__1425 (
            .O(N__10461),
            .I(N__10458));
    LocalMux I__1424 (
            .O(N__10458),
            .I(\POWERLED.un1_countlto15_5 ));
    InMux I__1423 (
            .O(N__10455),
            .I(N__10452));
    LocalMux I__1422 (
            .O(N__10452),
            .I(\POWERLED.un1_countlto15_7 ));
    IoInMux I__1421 (
            .O(N__10449),
            .I(N__10445));
    InMux I__1420 (
            .O(N__10448),
            .I(N__10442));
    LocalMux I__1419 (
            .O(N__10445),
            .I(N__10439));
    LocalMux I__1418 (
            .O(N__10442),
            .I(N__10436));
    IoSpan4Mux I__1417 (
            .O(N__10439),
            .I(N__10433));
    Span4Mux_v I__1416 (
            .O(N__10436),
            .I(N__10428));
    Span4Mux_s1_h I__1415 (
            .O(N__10433),
            .I(N__10428));
    Odrv4 I__1414 (
            .O(N__10428),
            .I(tmp_RNIRH3P));
    InMux I__1413 (
            .O(N__10425),
            .I(N__10422));
    LocalMux I__1412 (
            .O(N__10422),
            .I(\POWERLED.mult1_un110_sum_i ));
    InMux I__1411 (
            .O(N__10419),
            .I(N__10413));
    InMux I__1410 (
            .O(N__10418),
            .I(N__10413));
    LocalMux I__1409 (
            .O(N__10413),
            .I(\COUNTER.tmp_i ));
    CascadeMux I__1408 (
            .O(N__10410),
            .I(N__10407));
    InMux I__1407 (
            .O(N__10407),
            .I(N__10404));
    LocalMux I__1406 (
            .O(N__10404),
            .I(\POWERLED.mult1_un110_sum_cry_3_s ));
    InMux I__1405 (
            .O(N__10401),
            .I(\POWERLED.mult1_un110_sum_cry_2 ));
    InMux I__1404 (
            .O(N__10398),
            .I(N__10395));
    LocalMux I__1403 (
            .O(N__10395),
            .I(\POWERLED.mult1_un110_sum_cry_4_s ));
    InMux I__1402 (
            .O(N__10392),
            .I(\POWERLED.mult1_un110_sum_cry_3 ));
    CascadeMux I__1401 (
            .O(N__10389),
            .I(N__10386));
    InMux I__1400 (
            .O(N__10386),
            .I(N__10383));
    LocalMux I__1399 (
            .O(N__10383),
            .I(\POWERLED.mult1_un110_sum_cry_5_s ));
    InMux I__1398 (
            .O(N__10380),
            .I(\POWERLED.mult1_un110_sum_cry_4 ));
    InMux I__1397 (
            .O(N__10377),
            .I(N__10374));
    LocalMux I__1396 (
            .O(N__10374),
            .I(\VPP_VDDQ.un6_count_10 ));
    CascadeMux I__1395 (
            .O(N__10371),
            .I(\VPP_VDDQ.un6_count_9_cascade_ ));
    InMux I__1394 (
            .O(N__10368),
            .I(N__10365));
    LocalMux I__1393 (
            .O(N__10365),
            .I(\VPP_VDDQ.un6_count_8 ));
    InMux I__1392 (
            .O(N__10362),
            .I(N__10359));
    LocalMux I__1391 (
            .O(N__10359),
            .I(\VPP_VDDQ.un6_count_11 ));
    InMux I__1390 (
            .O(N__10356),
            .I(N__10353));
    LocalMux I__1389 (
            .O(N__10353),
            .I(N__10350));
    Span4Mux_s2_h I__1388 (
            .O(N__10350),
            .I(N__10347));
    Span4Mux_v I__1387 (
            .O(N__10347),
            .I(N__10343));
    InMux I__1386 (
            .O(N__10346),
            .I(N__10340));
    Odrv4 I__1385 (
            .O(N__10343),
            .I(\POWERLED.count_RNIOVT24Z0Z_11 ));
    LocalMux I__1384 (
            .O(N__10340),
            .I(\POWERLED.count_RNIOVT24Z0Z_11 ));
    CascadeMux I__1383 (
            .O(N__10335),
            .I(N__10332));
    InMux I__1382 (
            .O(N__10332),
            .I(N__10329));
    LocalMux I__1381 (
            .O(N__10329),
            .I(\POWERLED.un1_countlto15_4 ));
    CascadeMux I__1380 (
            .O(N__10326),
            .I(N__10323));
    InMux I__1379 (
            .O(N__10323),
            .I(N__10320));
    LocalMux I__1378 (
            .O(N__10320),
            .I(\POWERLED.un1_dutycycle_1_i_29 ));
    CascadeMux I__1377 (
            .O(N__10317),
            .I(N__10314));
    InMux I__1376 (
            .O(N__10314),
            .I(N__10311));
    LocalMux I__1375 (
            .O(N__10311),
            .I(N__10308));
    Odrv4 I__1374 (
            .O(N__10308),
            .I(\POWERLED.un1_dutycycle_1_i_28 ));
    CascadeMux I__1373 (
            .O(N__10305),
            .I(N__10302));
    InMux I__1372 (
            .O(N__10302),
            .I(N__10299));
    LocalMux I__1371 (
            .O(N__10299),
            .I(\POWERLED.mult1_un47_sum_axb_4 ));
    CascadeMux I__1370 (
            .O(N__10296),
            .I(vccst_en_cascade_));
    CascadeMux I__1369 (
            .O(N__10293),
            .I(N__10290));
    InMux I__1368 (
            .O(N__10290),
            .I(N__10287));
    LocalMux I__1367 (
            .O(N__10287),
            .I(N__10284));
    Odrv4 I__1366 (
            .O(N__10284),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_5 ));
    InMux I__1365 (
            .O(N__10281),
            .I(N__10278));
    LocalMux I__1364 (
            .O(N__10278),
            .I(N__10271));
    CascadeMux I__1363 (
            .O(N__10277),
            .I(N__10268));
    InMux I__1362 (
            .O(N__10276),
            .I(N__10265));
    InMux I__1361 (
            .O(N__10275),
            .I(N__10262));
    InMux I__1360 (
            .O(N__10274),
            .I(N__10259));
    Span4Mux_h I__1359 (
            .O(N__10271),
            .I(N__10256));
    InMux I__1358 (
            .O(N__10268),
            .I(N__10253));
    LocalMux I__1357 (
            .O(N__10265),
            .I(N__10248));
    LocalMux I__1356 (
            .O(N__10262),
            .I(N__10248));
    LocalMux I__1355 (
            .O(N__10259),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    Odrv4 I__1354 (
            .O(N__10256),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__1353 (
            .O(N__10253),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    Odrv12 I__1352 (
            .O(N__10248),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    InMux I__1351 (
            .O(N__10239),
            .I(N__10235));
    InMux I__1350 (
            .O(N__10238),
            .I(N__10231));
    LocalMux I__1349 (
            .O(N__10235),
            .I(N__10228));
    InMux I__1348 (
            .O(N__10234),
            .I(N__10225));
    LocalMux I__1347 (
            .O(N__10231),
            .I(N__10222));
    Span4Mux_h I__1346 (
            .O(N__10228),
            .I(N__10217));
    LocalMux I__1345 (
            .O(N__10225),
            .I(N__10217));
    Odrv12 I__1344 (
            .O(N__10222),
            .I(\RSMRST_PWRGD.N_240 ));
    Odrv4 I__1343 (
            .O(N__10217),
            .I(\RSMRST_PWRGD.N_240 ));
    InMux I__1342 (
            .O(N__10212),
            .I(N__10209));
    LocalMux I__1341 (
            .O(N__10209),
            .I(N__10206));
    Span4Mux_s3_h I__1340 (
            .O(N__10206),
            .I(N__10203));
    Odrv4 I__1339 (
            .O(N__10203),
            .I(\POWERLED.un1_count_2_15 ));
    CascadeMux I__1338 (
            .O(N__10200),
            .I(N__10197));
    InMux I__1337 (
            .O(N__10197),
            .I(N__10194));
    LocalMux I__1336 (
            .O(N__10194),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    InMux I__1335 (
            .O(N__10191),
            .I(\POWERLED.mult1_un47_sum_cry_2 ));
    CascadeMux I__1334 (
            .O(N__10188),
            .I(N__10185));
    InMux I__1333 (
            .O(N__10185),
            .I(N__10182));
    LocalMux I__1332 (
            .O(N__10182),
            .I(\POWERLED.mult1_un47_sum_cry_4_s ));
    InMux I__1331 (
            .O(N__10179),
            .I(\POWERLED.mult1_un47_sum_cry_3 ));
    CascadeMux I__1330 (
            .O(N__10176),
            .I(N__10173));
    InMux I__1329 (
            .O(N__10173),
            .I(N__10170));
    LocalMux I__1328 (
            .O(N__10170),
            .I(\POWERLED.mult1_un47_sum_cry_5_s ));
    InMux I__1327 (
            .O(N__10167),
            .I(\POWERLED.mult1_un47_sum_cry_4 ));
    InMux I__1326 (
            .O(N__10164),
            .I(\POWERLED.mult1_un47_sum_cry_5 ));
    CascadeMux I__1325 (
            .O(N__10161),
            .I(N__10158));
    InMux I__1324 (
            .O(N__10158),
            .I(N__10155));
    LocalMux I__1323 (
            .O(N__10155),
            .I(\POWERLED.mult1_un54_sum_cry_7_THRU_CO ));
    InMux I__1322 (
            .O(N__10152),
            .I(\POWERLED.mult1_un47_sum_cry_6 ));
    CascadeMux I__1321 (
            .O(N__10149),
            .I(\POWERLED.mult1_un54_sum_s_8_cascade_ ));
    InMux I__1320 (
            .O(N__10146),
            .I(N__10143));
    LocalMux I__1319 (
            .O(N__10143),
            .I(N__10139));
    InMux I__1318 (
            .O(N__10142),
            .I(N__10136));
    Span4Mux_v I__1317 (
            .O(N__10139),
            .I(N__10130));
    LocalMux I__1316 (
            .O(N__10136),
            .I(N__10130));
    CascadeMux I__1315 (
            .O(N__10135),
            .I(N__10126));
    Span4Mux_h I__1314 (
            .O(N__10130),
            .I(N__10123));
    InMux I__1313 (
            .O(N__10129),
            .I(N__10120));
    InMux I__1312 (
            .O(N__10126),
            .I(N__10117));
    Span4Mux_s0_h I__1311 (
            .O(N__10123),
            .I(N__10114));
    LocalMux I__1310 (
            .O(N__10120),
            .I(\POWERLED.curr_state_0_0 ));
    LocalMux I__1309 (
            .O(N__10117),
            .I(\POWERLED.curr_state_0_0 ));
    Odrv4 I__1308 (
            .O(N__10114),
            .I(\POWERLED.curr_state_0_0 ));
    IoInMux I__1307 (
            .O(N__10107),
            .I(N__10104));
    LocalMux I__1306 (
            .O(N__10104),
            .I(N__10101));
    Span4Mux_s1_v I__1305 (
            .O(N__10101),
            .I(N__10098));
    Span4Mux_v I__1304 (
            .O(N__10098),
            .I(N__10095));
    Span4Mux_v I__1303 (
            .O(N__10095),
            .I(N__10092));
    Odrv4 I__1302 (
            .O(N__10092),
            .I(pwrbtn_led));
    CEMux I__1301 (
            .O(N__10089),
            .I(N__10086));
    LocalMux I__1300 (
            .O(N__10086),
            .I(N__10083));
    Span4Mux_v I__1299 (
            .O(N__10083),
            .I(N__10080));
    Odrv4 I__1298 (
            .O(N__10080),
            .I(\POWERLED.pwm_out_RNOZ0 ));
    InMux I__1297 (
            .O(N__10077),
            .I(\POWERLED.mult1_un54_sum_cry_2 ));
    InMux I__1296 (
            .O(N__10074),
            .I(\POWERLED.mult1_un54_sum_cry_3 ));
    InMux I__1295 (
            .O(N__10071),
            .I(\POWERLED.mult1_un54_sum_cry_4 ));
    InMux I__1294 (
            .O(N__10068),
            .I(\POWERLED.mult1_un54_sum_cry_5 ));
    InMux I__1293 (
            .O(N__10065),
            .I(\POWERLED.mult1_un54_sum_cry_6 ));
    InMux I__1292 (
            .O(N__10062),
            .I(\POWERLED.mult1_un54_sum_cry_7 ));
    InMux I__1291 (
            .O(N__10059),
            .I(\POWERLED.mult1_un117_sum_cry_7 ));
    CascadeMux I__1290 (
            .O(N__10056),
            .I(N__10052));
    InMux I__1289 (
            .O(N__10055),
            .I(N__10046));
    InMux I__1288 (
            .O(N__10052),
            .I(N__10046));
    InMux I__1287 (
            .O(N__10051),
            .I(N__10043));
    LocalMux I__1286 (
            .O(N__10046),
            .I(N__10040));
    LocalMux I__1285 (
            .O(N__10043),
            .I(N__10036));
    Span4Mux_s3_h I__1284 (
            .O(N__10040),
            .I(N__10033));
    InMux I__1283 (
            .O(N__10039),
            .I(N__10030));
    Span4Mux_s3_h I__1282 (
            .O(N__10036),
            .I(N__10027));
    Odrv4 I__1281 (
            .O(N__10033),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__1280 (
            .O(N__10030),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    Odrv4 I__1279 (
            .O(N__10027),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    CascadeMux I__1278 (
            .O(N__10020),
            .I(\POWERLED.mult1_un117_sum_s_8_cascade_ ));
    InMux I__1277 (
            .O(N__10017),
            .I(N__10014));
    LocalMux I__1276 (
            .O(N__10014),
            .I(N__10011));
    Odrv4 I__1275 (
            .O(N__10011),
            .I(\POWERLED.un1_count_2_7 ));
    InMux I__1274 (
            .O(N__10008),
            .I(N__10005));
    LocalMux I__1273 (
            .O(N__10005),
            .I(N__10002));
    Odrv4 I__1272 (
            .O(N__10002),
            .I(\POWERLED.un1_count_2_14 ));
    InMux I__1271 (
            .O(N__9999),
            .I(N__9996));
    LocalMux I__1270 (
            .O(N__9996),
            .I(N__9993));
    Odrv4 I__1269 (
            .O(N__9993),
            .I(\POWERLED.un1_count_2_9 ));
    InMux I__1268 (
            .O(N__9990),
            .I(N__9987));
    LocalMux I__1267 (
            .O(N__9987),
            .I(N__9984));
    Odrv4 I__1266 (
            .O(N__9984),
            .I(\POWERLED.un1_count_2_8 ));
    CascadeMux I__1265 (
            .O(N__9981),
            .I(N__9977));
    CascadeMux I__1264 (
            .O(N__9980),
            .I(N__9973));
    InMux I__1263 (
            .O(N__9977),
            .I(N__9966));
    InMux I__1262 (
            .O(N__9976),
            .I(N__9966));
    InMux I__1261 (
            .O(N__9973),
            .I(N__9966));
    LocalMux I__1260 (
            .O(N__9966),
            .I(\POWERLED.mult1_un110_sum_i_0_8 ));
    CascadeMux I__1259 (
            .O(N__9963),
            .I(N__9960));
    InMux I__1258 (
            .O(N__9960),
            .I(N__9957));
    LocalMux I__1257 (
            .O(N__9957),
            .I(N__9954));
    Odrv4 I__1256 (
            .O(N__9954),
            .I(\POWERLED.un1_count_2_13 ));
    InMux I__1255 (
            .O(N__9951),
            .I(N__9948));
    LocalMux I__1254 (
            .O(N__9948),
            .I(N__9945));
    Odrv4 I__1253 (
            .O(N__9945),
            .I(\POWERLED.un1_count_2_10 ));
    InMux I__1252 (
            .O(N__9942),
            .I(N__9939));
    LocalMux I__1251 (
            .O(N__9939),
            .I(N__9936));
    Odrv4 I__1250 (
            .O(N__9936),
            .I(\POWERLED.un1_count_2_11 ));
    InMux I__1249 (
            .O(N__9933),
            .I(N__9930));
    LocalMux I__1248 (
            .O(N__9930),
            .I(\POWERLED.un1_countlt6_0 ));
    CascadeMux I__1247 (
            .O(N__9927),
            .I(\POWERLED.g0_0_5_cascade_ ));
    InMux I__1246 (
            .O(N__9924),
            .I(N__9921));
    LocalMux I__1245 (
            .O(N__9921),
            .I(\POWERLED.g0_0_7 ));
    CascadeMux I__1244 (
            .O(N__9918),
            .I(N__9915));
    InMux I__1243 (
            .O(N__9915),
            .I(N__9912));
    LocalMux I__1242 (
            .O(N__9912),
            .I(N__9909));
    Span4Mux_s3_h I__1241 (
            .O(N__9909),
            .I(N__9906));
    Odrv4 I__1240 (
            .O(N__9906),
            .I(\POWERLED.mult1_un117_sum_cry_3_s ));
    InMux I__1239 (
            .O(N__9903),
            .I(\POWERLED.mult1_un117_sum_cry_2 ));
    InMux I__1238 (
            .O(N__9900),
            .I(N__9897));
    LocalMux I__1237 (
            .O(N__9897),
            .I(N__9894));
    Span4Mux_s3_h I__1236 (
            .O(N__9894),
            .I(N__9891));
    Odrv4 I__1235 (
            .O(N__9891),
            .I(\POWERLED.mult1_un117_sum_cry_4_s ));
    InMux I__1234 (
            .O(N__9888),
            .I(\POWERLED.mult1_un117_sum_cry_3 ));
    CascadeMux I__1233 (
            .O(N__9885),
            .I(N__9882));
    InMux I__1232 (
            .O(N__9882),
            .I(N__9879));
    LocalMux I__1231 (
            .O(N__9879),
            .I(N__9876));
    Span4Mux_s3_h I__1230 (
            .O(N__9876),
            .I(N__9873));
    Odrv4 I__1229 (
            .O(N__9873),
            .I(\POWERLED.mult1_un117_sum_cry_5_s ));
    InMux I__1228 (
            .O(N__9870),
            .I(\POWERLED.mult1_un117_sum_cry_4 ));
    InMux I__1227 (
            .O(N__9867),
            .I(N__9864));
    LocalMux I__1226 (
            .O(N__9864),
            .I(N__9861));
    Span4Mux_v I__1225 (
            .O(N__9861),
            .I(N__9858));
    Odrv4 I__1224 (
            .O(N__9858),
            .I(\POWERLED.mult1_un117_sum_cry_6_s ));
    InMux I__1223 (
            .O(N__9855),
            .I(\POWERLED.mult1_un117_sum_cry_5 ));
    CascadeMux I__1222 (
            .O(N__9852),
            .I(N__9849));
    InMux I__1221 (
            .O(N__9849),
            .I(N__9846));
    LocalMux I__1220 (
            .O(N__9846),
            .I(N__9843));
    Span4Mux_v I__1219 (
            .O(N__9843),
            .I(N__9840));
    Odrv4 I__1218 (
            .O(N__9840),
            .I(\POWERLED.mult1_un124_sum_axb_8 ));
    InMux I__1217 (
            .O(N__9837),
            .I(\POWERLED.mult1_un117_sum_cry_6 ));
    InMux I__1216 (
            .O(N__9834),
            .I(N__9831));
    LocalMux I__1215 (
            .O(N__9831),
            .I(\RSMRST_PWRGD.m4_i_i_a2_0_10 ));
    InMux I__1214 (
            .O(N__9828),
            .I(N__9825));
    LocalMux I__1213 (
            .O(N__9825),
            .I(\RSMRST_PWRGD.m4_i_i_a2_0_11 ));
    CascadeMux I__1212 (
            .O(N__9822),
            .I(\RSMRST_PWRGD.m4_i_i_a2_0_9_cascade_ ));
    InMux I__1211 (
            .O(N__9819),
            .I(N__9816));
    LocalMux I__1210 (
            .O(N__9816),
            .I(\RSMRST_PWRGD.m4_i_i_a2_0_12 ));
    SRMux I__1209 (
            .O(N__9813),
            .I(N__9809));
    SRMux I__1208 (
            .O(N__9812),
            .I(N__9806));
    LocalMux I__1207 (
            .O(N__9809),
            .I(N__9802));
    LocalMux I__1206 (
            .O(N__9806),
            .I(N__9799));
    SRMux I__1205 (
            .O(N__9805),
            .I(N__9796));
    Span4Mux_v I__1204 (
            .O(N__9802),
            .I(N__9793));
    Span4Mux_s1_h I__1203 (
            .O(N__9799),
            .I(N__9790));
    LocalMux I__1202 (
            .O(N__9796),
            .I(N__9787));
    Odrv4 I__1201 (
            .O(N__9793),
            .I(\RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0 ));
    Odrv4 I__1200 (
            .O(N__9790),
            .I(\RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0 ));
    Odrv12 I__1199 (
            .O(N__9787),
            .I(\RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0 ));
    CascadeMux I__1198 (
            .O(N__9780),
            .I(\RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0_cascade_ ));
    CEMux I__1197 (
            .O(N__9777),
            .I(N__9774));
    LocalMux I__1196 (
            .O(N__9774),
            .I(N__9771));
    Span4Mux_s2_h I__1195 (
            .O(N__9771),
            .I(N__9768));
    Odrv4 I__1194 (
            .O(N__9768),
            .I(\RSMRST_PWRGD.N_49_2 ));
    IoInMux I__1193 (
            .O(N__9765),
            .I(N__9762));
    LocalMux I__1192 (
            .O(N__9762),
            .I(N__9758));
    IoInMux I__1191 (
            .O(N__9761),
            .I(N__9755));
    Span4Mux_s1_h I__1190 (
            .O(N__9758),
            .I(N__9752));
    LocalMux I__1189 (
            .O(N__9755),
            .I(N__9749));
    Odrv4 I__1188 (
            .O(N__9752),
            .I(v5s_enn));
    Odrv4 I__1187 (
            .O(N__9749),
            .I(v5s_enn));
    InMux I__1186 (
            .O(N__9744),
            .I(N__9740));
    InMux I__1185 (
            .O(N__9743),
            .I(N__9737));
    LocalMux I__1184 (
            .O(N__9740),
            .I(N__9733));
    LocalMux I__1183 (
            .O(N__9737),
            .I(N__9730));
    InMux I__1182 (
            .O(N__9736),
            .I(N__9727));
    Odrv4 I__1181 (
            .O(N__9733),
            .I(\RSMRST_PWRGD.N_241 ));
    Odrv4 I__1180 (
            .O(N__9730),
            .I(\RSMRST_PWRGD.N_241 ));
    LocalMux I__1179 (
            .O(N__9727),
            .I(\RSMRST_PWRGD.N_241 ));
    CascadeMux I__1178 (
            .O(N__9720),
            .I(\POWERLED.g0_0_4_cascade_ ));
    InMux I__1177 (
            .O(N__9717),
            .I(N__9714));
    LocalMux I__1176 (
            .O(N__9714),
            .I(N__9711));
    Span4Mux_s3_h I__1175 (
            .O(N__9711),
            .I(N__9708));
    Odrv4 I__1174 (
            .O(N__9708),
            .I(\POWERLED.un1_count_0 ));
    CascadeMux I__1173 (
            .O(N__9705),
            .I(N__9701));
    InMux I__1172 (
            .O(N__9704),
            .I(N__9698));
    InMux I__1171 (
            .O(N__9701),
            .I(N__9695));
    LocalMux I__1170 (
            .O(N__9698),
            .I(\RSMRST_PWRGD.N_37 ));
    LocalMux I__1169 (
            .O(N__9695),
            .I(\RSMRST_PWRGD.N_37 ));
    InMux I__1168 (
            .O(N__9690),
            .I(N__9686));
    InMux I__1167 (
            .O(N__9689),
            .I(N__9683));
    LocalMux I__1166 (
            .O(N__9686),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    LocalMux I__1165 (
            .O(N__9683),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    InMux I__1164 (
            .O(N__9678),
            .I(N__9674));
    InMux I__1163 (
            .O(N__9677),
            .I(N__9671));
    LocalMux I__1162 (
            .O(N__9674),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    LocalMux I__1161 (
            .O(N__9671),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    CascadeMux I__1160 (
            .O(N__9666),
            .I(N__9662));
    CascadeMux I__1159 (
            .O(N__9665),
            .I(N__9657));
    InMux I__1158 (
            .O(N__9662),
            .I(N__9654));
    InMux I__1157 (
            .O(N__9661),
            .I(N__9647));
    InMux I__1156 (
            .O(N__9660),
            .I(N__9647));
    InMux I__1155 (
            .O(N__9657),
            .I(N__9647));
    LocalMux I__1154 (
            .O(N__9654),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__1153 (
            .O(N__9647),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    InMux I__1152 (
            .O(N__9642),
            .I(N__9638));
    InMux I__1151 (
            .O(N__9641),
            .I(N__9635));
    LocalMux I__1150 (
            .O(N__9638),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    LocalMux I__1149 (
            .O(N__9635),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    InMux I__1148 (
            .O(N__9630),
            .I(N__9626));
    InMux I__1147 (
            .O(N__9629),
            .I(N__9623));
    LocalMux I__1146 (
            .O(N__9626),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    LocalMux I__1145 (
            .O(N__9623),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    CascadeMux I__1144 (
            .O(N__9618),
            .I(N__9614));
    InMux I__1143 (
            .O(N__9617),
            .I(N__9611));
    InMux I__1142 (
            .O(N__9614),
            .I(N__9608));
    LocalMux I__1141 (
            .O(N__9611),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    LocalMux I__1140 (
            .O(N__9608),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    InMux I__1139 (
            .O(N__9603),
            .I(N__9599));
    InMux I__1138 (
            .O(N__9602),
            .I(N__9596));
    LocalMux I__1137 (
            .O(N__9599),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    LocalMux I__1136 (
            .O(N__9596),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    InMux I__1135 (
            .O(N__9591),
            .I(N__9587));
    InMux I__1134 (
            .O(N__9590),
            .I(N__9584));
    LocalMux I__1133 (
            .O(N__9587),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    LocalMux I__1132 (
            .O(N__9584),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    InMux I__1131 (
            .O(N__9579),
            .I(N__9575));
    InMux I__1130 (
            .O(N__9578),
            .I(N__9572));
    LocalMux I__1129 (
            .O(N__9575),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    LocalMux I__1128 (
            .O(N__9572),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    CascadeMux I__1127 (
            .O(N__9567),
            .I(N__9563));
    InMux I__1126 (
            .O(N__9566),
            .I(N__9560));
    InMux I__1125 (
            .O(N__9563),
            .I(N__9557));
    LocalMux I__1124 (
            .O(N__9560),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    LocalMux I__1123 (
            .O(N__9557),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    InMux I__1122 (
            .O(N__9552),
            .I(N__9548));
    InMux I__1121 (
            .O(N__9551),
            .I(N__9545));
    LocalMux I__1120 (
            .O(N__9548),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    LocalMux I__1119 (
            .O(N__9545),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    InMux I__1118 (
            .O(N__9540),
            .I(N__9536));
    InMux I__1117 (
            .O(N__9539),
            .I(N__9533));
    LocalMux I__1116 (
            .O(N__9536),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    LocalMux I__1115 (
            .O(N__9533),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    InMux I__1114 (
            .O(N__9528),
            .I(N__9524));
    InMux I__1113 (
            .O(N__9527),
            .I(N__9521));
    LocalMux I__1112 (
            .O(N__9524),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    LocalMux I__1111 (
            .O(N__9521),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    InMux I__1110 (
            .O(N__9516),
            .I(N__9513));
    LocalMux I__1109 (
            .O(N__9513),
            .I(\RSMRST_PWRGD.m4_i_i_a2_0_7 ));
    InMux I__1108 (
            .O(N__9510),
            .I(N__9506));
    InMux I__1107 (
            .O(N__9509),
            .I(N__9503));
    LocalMux I__1106 (
            .O(N__9506),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    LocalMux I__1105 (
            .O(N__9503),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    InMux I__1104 (
            .O(N__9498),
            .I(N__9494));
    InMux I__1103 (
            .O(N__9497),
            .I(N__9491));
    LocalMux I__1102 (
            .O(N__9494),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    LocalMux I__1101 (
            .O(N__9491),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    CascadeMux I__1100 (
            .O(N__9486),
            .I(N__9482));
    InMux I__1099 (
            .O(N__9485),
            .I(N__9479));
    InMux I__1098 (
            .O(N__9482),
            .I(N__9476));
    LocalMux I__1097 (
            .O(N__9479),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    LocalMux I__1096 (
            .O(N__9476),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    InMux I__1095 (
            .O(N__9471),
            .I(N__9467));
    InMux I__1094 (
            .O(N__9470),
            .I(N__9464));
    LocalMux I__1093 (
            .O(N__9467),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    LocalMux I__1092 (
            .O(N__9464),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    CascadeMux I__1091 (
            .O(N__9459),
            .I(N__9456));
    InMux I__1090 (
            .O(N__9456),
            .I(N__9452));
    InMux I__1089 (
            .O(N__9455),
            .I(N__9449));
    LocalMux I__1088 (
            .O(N__9452),
            .I(\POWERLED.un1_count_2_cry_15_THRU_CO ));
    LocalMux I__1087 (
            .O(N__9449),
            .I(\POWERLED.un1_count_2_cry_15_THRU_CO ));
    CascadeMux I__1086 (
            .O(N__9444),
            .I(N__9441));
    InMux I__1085 (
            .O(N__9441),
            .I(N__9438));
    LocalMux I__1084 (
            .O(N__9438),
            .I(\POWERLED.mult1_un159_sum_cry_2_s ));
    CascadeMux I__1083 (
            .O(N__9435),
            .I(N__9432));
    InMux I__1082 (
            .O(N__9432),
            .I(N__9429));
    LocalMux I__1081 (
            .O(N__9429),
            .I(\POWERLED.mult1_un159_sum_cry_3_s ));
    InMux I__1080 (
            .O(N__9426),
            .I(N__9423));
    LocalMux I__1079 (
            .O(N__9423),
            .I(\POWERLED.mult1_un159_sum_cry_4_s ));
    CascadeMux I__1078 (
            .O(N__9420),
            .I(N__9416));
    InMux I__1077 (
            .O(N__9419),
            .I(N__9411));
    InMux I__1076 (
            .O(N__9416),
            .I(N__9404));
    InMux I__1075 (
            .O(N__9415),
            .I(N__9404));
    InMux I__1074 (
            .O(N__9414),
            .I(N__9404));
    LocalMux I__1073 (
            .O(N__9411),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__1072 (
            .O(N__9404),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    InMux I__1071 (
            .O(N__9399),
            .I(N__9396));
    LocalMux I__1070 (
            .O(N__9396),
            .I(\POWERLED.mult1_un159_sum_cry_5_s ));
    CascadeMux I__1069 (
            .O(N__9393),
            .I(N__9389));
    CascadeMux I__1068 (
            .O(N__9392),
            .I(N__9385));
    InMux I__1067 (
            .O(N__9389),
            .I(N__9378));
    InMux I__1066 (
            .O(N__9388),
            .I(N__9378));
    InMux I__1065 (
            .O(N__9385),
            .I(N__9378));
    LocalMux I__1064 (
            .O(N__9378),
            .I(G_385));
    CascadeMux I__1063 (
            .O(N__9375),
            .I(N__9372));
    InMux I__1062 (
            .O(N__9372),
            .I(N__9369));
    LocalMux I__1061 (
            .O(N__9369),
            .I(\POWERLED.mult1_un166_sum_axb_6 ));
    InMux I__1060 (
            .O(N__9366),
            .I(\POWERLED.mult1_un166_sum_cry_5 ));
    CascadeMux I__1059 (
            .O(N__9363),
            .I(N__9360));
    InMux I__1058 (
            .O(N__9360),
            .I(N__9357));
    LocalMux I__1057 (
            .O(N__9357),
            .I(N__9354));
    Odrv12 I__1056 (
            .O(N__9354),
            .I(\POWERLED.un1_count_2_0 ));
    InMux I__1055 (
            .O(N__9351),
            .I(N__9348));
    LocalMux I__1054 (
            .O(N__9348),
            .I(\POWERLED.mult1_un159_sum_i ));
    CascadeMux I__1053 (
            .O(N__9345),
            .I(N__9342));
    InMux I__1052 (
            .O(N__9342),
            .I(N__9339));
    LocalMux I__1051 (
            .O(N__9339),
            .I(\POWERLED.count_i_14 ));
    CascadeMux I__1050 (
            .O(N__9336),
            .I(N__9333));
    InMux I__1049 (
            .O(N__9333),
            .I(N__9330));
    LocalMux I__1048 (
            .O(N__9330),
            .I(\POWERLED.count_i_15 ));
    InMux I__1047 (
            .O(N__9327),
            .I(bfn_2_7_0_));
    InMux I__1046 (
            .O(N__9324),
            .I(N__9321));
    LocalMux I__1045 (
            .O(N__9321),
            .I(N__9318));
    Odrv4 I__1044 (
            .O(N__9318),
            .I(\POWERLED.mult1_un138_sum_i ));
    InMux I__1043 (
            .O(N__9315),
            .I(N__9312));
    LocalMux I__1042 (
            .O(N__9312),
            .I(N__9307));
    IoInMux I__1041 (
            .O(N__9311),
            .I(N__9304));
    IoInMux I__1040 (
            .O(N__9310),
            .I(N__9301));
    Span4Mux_h I__1039 (
            .O(N__9307),
            .I(N__9298));
    LocalMux I__1038 (
            .O(N__9304),
            .I(N__9295));
    LocalMux I__1037 (
            .O(N__9301),
            .I(N__9292));
    Span4Mux_h I__1036 (
            .O(N__9298),
            .I(N__9289));
    IoSpan4Mux I__1035 (
            .O(N__9295),
            .I(N__9286));
    Span12Mux_s8_h I__1034 (
            .O(N__9292),
            .I(N__9283));
    Sp12to4 I__1033 (
            .O(N__9289),
            .I(N__9280));
    IoSpan4Mux I__1032 (
            .O(N__9286),
            .I(N__9277));
    Odrv12 I__1031 (
            .O(N__9283),
            .I(slp_susn));
    Odrv12 I__1030 (
            .O(N__9280),
            .I(slp_susn));
    Odrv4 I__1029 (
            .O(N__9277),
            .I(slp_susn));
    InMux I__1028 (
            .O(N__9270),
            .I(N__9267));
    LocalMux I__1027 (
            .O(N__9267),
            .I(N__9264));
    Span4Mux_v I__1026 (
            .O(N__9264),
            .I(N__9261));
    Odrv4 I__1025 (
            .O(N__9261),
            .I(v5a_ok));
    CascadeMux I__1024 (
            .O(N__9258),
            .I(N__9255));
    InMux I__1023 (
            .O(N__9255),
            .I(N__9252));
    LocalMux I__1022 (
            .O(N__9252),
            .I(N__9249));
    Span4Mux_s3_h I__1021 (
            .O(N__9249),
            .I(N__9246));
    Sp12to4 I__1020 (
            .O(N__9246),
            .I(N__9243));
    Span12Mux_v I__1019 (
            .O(N__9243),
            .I(N__9240));
    Odrv12 I__1018 (
            .O(N__9240),
            .I(v33a_ok));
    IoInMux I__1017 (
            .O(N__9237),
            .I(N__9234));
    LocalMux I__1016 (
            .O(N__9234),
            .I(N__9231));
    Span4Mux_s2_h I__1015 (
            .O(N__9231),
            .I(N__9227));
    InMux I__1014 (
            .O(N__9230),
            .I(N__9224));
    Sp12to4 I__1013 (
            .O(N__9227),
            .I(N__9221));
    LocalMux I__1012 (
            .O(N__9224),
            .I(N__9218));
    Span12Mux_s11_v I__1011 (
            .O(N__9221),
            .I(N__9215));
    Span12Mux_s11_v I__1010 (
            .O(N__9218),
            .I(N__9212));
    Odrv12 I__1009 (
            .O(N__9215),
            .I(v1p8a_ok));
    Odrv12 I__1008 (
            .O(N__9212),
            .I(v1p8a_ok));
    InMux I__1007 (
            .O(N__9207),
            .I(N__9204));
    LocalMux I__1006 (
            .O(N__9204),
            .I(\POWERLED.mult1_un152_sum_i ));
    CascadeMux I__1005 (
            .O(N__9201),
            .I(N__9196));
    InMux I__1004 (
            .O(N__9200),
            .I(N__9192));
    InMux I__1003 (
            .O(N__9199),
            .I(N__9187));
    InMux I__1002 (
            .O(N__9196),
            .I(N__9187));
    InMux I__1001 (
            .O(N__9195),
            .I(N__9184));
    LocalMux I__1000 (
            .O(N__9192),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__999 (
            .O(N__9187),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__998 (
            .O(N__9184),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    InMux I__997 (
            .O(N__9177),
            .I(N__9174));
    LocalMux I__996 (
            .O(N__9174),
            .I(N__9171));
    Odrv4 I__995 (
            .O(N__9171),
            .I(\POWERLED.un1_count_2_2 ));
    InMux I__994 (
            .O(N__9168),
            .I(N__9165));
    LocalMux I__993 (
            .O(N__9165),
            .I(\POWERLED.un1_count_2_12 ));
    CascadeMux I__992 (
            .O(N__9162),
            .I(N__9159));
    InMux I__991 (
            .O(N__9159),
            .I(N__9156));
    LocalMux I__990 (
            .O(N__9156),
            .I(\POWERLED.un1_count_2_5 ));
    InMux I__989 (
            .O(N__9153),
            .I(N__9150));
    LocalMux I__988 (
            .O(N__9150),
            .I(\POWERLED.count_i_5 ));
    InMux I__987 (
            .O(N__9147),
            .I(N__9144));
    LocalMux I__986 (
            .O(N__9144),
            .I(\POWERLED.un1_count_2_6 ));
    CascadeMux I__985 (
            .O(N__9141),
            .I(N__9138));
    InMux I__984 (
            .O(N__9138),
            .I(N__9135));
    LocalMux I__983 (
            .O(N__9135),
            .I(\POWERLED.count_i_6 ));
    CascadeMux I__982 (
            .O(N__9132),
            .I(N__9129));
    InMux I__981 (
            .O(N__9129),
            .I(N__9126));
    LocalMux I__980 (
            .O(N__9126),
            .I(\POWERLED.count_i_7 ));
    CascadeMux I__979 (
            .O(N__9123),
            .I(N__9120));
    InMux I__978 (
            .O(N__9120),
            .I(N__9117));
    LocalMux I__977 (
            .O(N__9117),
            .I(\POWERLED.count_i_8 ));
    CascadeMux I__976 (
            .O(N__9114),
            .I(N__9111));
    InMux I__975 (
            .O(N__9111),
            .I(N__9108));
    LocalMux I__974 (
            .O(N__9108),
            .I(\POWERLED.count_i_9 ));
    CascadeMux I__973 (
            .O(N__9105),
            .I(N__9102));
    InMux I__972 (
            .O(N__9102),
            .I(N__9099));
    LocalMux I__971 (
            .O(N__9099),
            .I(\POWERLED.count_i_10 ));
    CascadeMux I__970 (
            .O(N__9096),
            .I(N__9093));
    InMux I__969 (
            .O(N__9093),
            .I(N__9090));
    LocalMux I__968 (
            .O(N__9090),
            .I(\POWERLED.count_i_11 ));
    CascadeMux I__967 (
            .O(N__9087),
            .I(N__9084));
    InMux I__966 (
            .O(N__9084),
            .I(N__9081));
    LocalMux I__965 (
            .O(N__9081),
            .I(\POWERLED.count_i_12 ));
    InMux I__964 (
            .O(N__9078),
            .I(N__9075));
    LocalMux I__963 (
            .O(N__9075),
            .I(\POWERLED.count_i_13 ));
    InMux I__962 (
            .O(N__9072),
            .I(N__9068));
    CascadeMux I__961 (
            .O(N__9071),
            .I(N__9064));
    LocalMux I__960 (
            .O(N__9068),
            .I(N__9059));
    InMux I__959 (
            .O(N__9067),
            .I(N__9054));
    InMux I__958 (
            .O(N__9064),
            .I(N__9054));
    InMux I__957 (
            .O(N__9063),
            .I(N__9051));
    InMux I__956 (
            .O(N__9062),
            .I(N__9048));
    Odrv4 I__955 (
            .O(N__9059),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__954 (
            .O(N__9054),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__953 (
            .O(N__9051),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__952 (
            .O(N__9048),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    CascadeMux I__951 (
            .O(N__9039),
            .I(N__9035));
    InMux I__950 (
            .O(N__9038),
            .I(N__9029));
    InMux I__949 (
            .O(N__9035),
            .I(N__9029));
    InMux I__948 (
            .O(N__9034),
            .I(N__9022));
    LocalMux I__947 (
            .O(N__9029),
            .I(N__9019));
    InMux I__946 (
            .O(N__9028),
            .I(N__9016));
    InMux I__945 (
            .O(N__9027),
            .I(N__9009));
    InMux I__944 (
            .O(N__9026),
            .I(N__9009));
    InMux I__943 (
            .O(N__9025),
            .I(N__9009));
    LocalMux I__942 (
            .O(N__9022),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    Odrv4 I__941 (
            .O(N__9019),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__940 (
            .O(N__9016),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__939 (
            .O(N__9009),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    CascadeMux I__938 (
            .O(N__9000),
            .I(N__8995));
    InMux I__937 (
            .O(N__8999),
            .I(N__8990));
    InMux I__936 (
            .O(N__8998),
            .I(N__8985));
    InMux I__935 (
            .O(N__8995),
            .I(N__8985));
    InMux I__934 (
            .O(N__8994),
            .I(N__8982));
    InMux I__933 (
            .O(N__8993),
            .I(N__8979));
    LocalMux I__932 (
            .O(N__8990),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__931 (
            .O(N__8985),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__930 (
            .O(N__8982),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__929 (
            .O(N__8979),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    InMux I__928 (
            .O(N__8970),
            .I(N__8967));
    LocalMux I__927 (
            .O(N__8967),
            .I(N__8964));
    Span4Mux_s2_h I__926 (
            .O(N__8964),
            .I(N__8961));
    Odrv4 I__925 (
            .O(N__8961),
            .I(\POWERLED.count_i_0_0 ));
    CascadeMux I__924 (
            .O(N__8958),
            .I(N__8955));
    InMux I__923 (
            .O(N__8955),
            .I(N__8952));
    LocalMux I__922 (
            .O(N__8952),
            .I(N__8949));
    Odrv4 I__921 (
            .O(N__8949),
            .I(\POWERLED.un1_count_2_1 ));
    InMux I__920 (
            .O(N__8946),
            .I(N__8943));
    LocalMux I__919 (
            .O(N__8943),
            .I(\POWERLED.count_i_1 ));
    CascadeMux I__918 (
            .O(N__8940),
            .I(N__8937));
    InMux I__917 (
            .O(N__8937),
            .I(N__8934));
    LocalMux I__916 (
            .O(N__8934),
            .I(\POWERLED.count_i_2 ));
    InMux I__915 (
            .O(N__8931),
            .I(N__8928));
    LocalMux I__914 (
            .O(N__8928),
            .I(\POWERLED.un1_count_2_3 ));
    CascadeMux I__913 (
            .O(N__8925),
            .I(N__8922));
    InMux I__912 (
            .O(N__8922),
            .I(N__8919));
    LocalMux I__911 (
            .O(N__8919),
            .I(N__8916));
    Odrv4 I__910 (
            .O(N__8916),
            .I(\POWERLED.count_i_3 ));
    InMux I__909 (
            .O(N__8913),
            .I(N__8910));
    LocalMux I__908 (
            .O(N__8910),
            .I(\POWERLED.un1_count_2_4 ));
    CascadeMux I__907 (
            .O(N__8907),
            .I(N__8904));
    InMux I__906 (
            .O(N__8904),
            .I(N__8901));
    LocalMux I__905 (
            .O(N__8901),
            .I(\POWERLED.count_i_4 ));
    CascadeMux I__904 (
            .O(N__8898),
            .I(N__8895));
    InMux I__903 (
            .O(N__8895),
            .I(N__8892));
    LocalMux I__902 (
            .O(N__8892),
            .I(\POWERLED.mult1_un124_sum_cry_5_s ));
    InMux I__901 (
            .O(N__8889),
            .I(\POWERLED.mult1_un124_sum_cry_4 ));
    InMux I__900 (
            .O(N__8886),
            .I(N__8883));
    LocalMux I__899 (
            .O(N__8883),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    InMux I__898 (
            .O(N__8880),
            .I(\POWERLED.mult1_un124_sum_cry_5 ));
    InMux I__897 (
            .O(N__8877),
            .I(N__8874));
    LocalMux I__896 (
            .O(N__8874),
            .I(\POWERLED.mult1_un131_sum_axb_8 ));
    InMux I__895 (
            .O(N__8871),
            .I(\POWERLED.mult1_un124_sum_cry_6 ));
    InMux I__894 (
            .O(N__8868),
            .I(\POWERLED.mult1_un124_sum_cry_7 ));
    CascadeMux I__893 (
            .O(N__8865),
            .I(N__8861));
    CascadeMux I__892 (
            .O(N__8864),
            .I(N__8857));
    InMux I__891 (
            .O(N__8861),
            .I(N__8850));
    InMux I__890 (
            .O(N__8860),
            .I(N__8850));
    InMux I__889 (
            .O(N__8857),
            .I(N__8850));
    LocalMux I__888 (
            .O(N__8850),
            .I(\POWERLED.mult1_un124_sum_i_0_8 ));
    InMux I__887 (
            .O(N__8847),
            .I(N__8844));
    LocalMux I__886 (
            .O(N__8844),
            .I(\POWERLED.mult1_un131_sum_i ));
    InMux I__885 (
            .O(N__8841),
            .I(N__8838));
    LocalMux I__884 (
            .O(N__8838),
            .I(\POWERLED.mult1_un124_sum_i ));
    CascadeMux I__883 (
            .O(N__8835),
            .I(N__8831));
    CascadeMux I__882 (
            .O(N__8834),
            .I(N__8827));
    InMux I__881 (
            .O(N__8831),
            .I(N__8820));
    InMux I__880 (
            .O(N__8830),
            .I(N__8820));
    InMux I__879 (
            .O(N__8827),
            .I(N__8820));
    LocalMux I__878 (
            .O(N__8820),
            .I(\POWERLED.mult1_un117_sum_i_0_8 ));
    InMux I__877 (
            .O(N__8817),
            .I(N__8814));
    LocalMux I__876 (
            .O(N__8814),
            .I(\POWERLED.mult1_un117_sum_i ));
    InMux I__875 (
            .O(N__8811),
            .I(\RSMRST_PWRGD.un1_count_1_cry_11 ));
    InMux I__874 (
            .O(N__8808),
            .I(\RSMRST_PWRGD.un1_count_1_cry_12 ));
    InMux I__873 (
            .O(N__8805),
            .I(\RSMRST_PWRGD.un1_count_1_cry_13 ));
    InMux I__872 (
            .O(N__8802),
            .I(bfn_1_12_0_));
    InMux I__871 (
            .O(N__8799),
            .I(N__8796));
    LocalMux I__870 (
            .O(N__8796),
            .I(vpp_ok));
    IoInMux I__869 (
            .O(N__8793),
            .I(N__8790));
    LocalMux I__868 (
            .O(N__8790),
            .I(N__8787));
    Odrv12 I__867 (
            .O(N__8787),
            .I(vddq_en));
    CascadeMux I__866 (
            .O(N__8784),
            .I(N__8781));
    InMux I__865 (
            .O(N__8781),
            .I(N__8778));
    LocalMux I__864 (
            .O(N__8778),
            .I(\POWERLED.mult1_un124_sum_cry_3_s ));
    InMux I__863 (
            .O(N__8775),
            .I(\POWERLED.mult1_un124_sum_cry_2 ));
    InMux I__862 (
            .O(N__8772),
            .I(N__8769));
    LocalMux I__861 (
            .O(N__8769),
            .I(\POWERLED.mult1_un124_sum_cry_4_s ));
    InMux I__860 (
            .O(N__8766),
            .I(\POWERLED.mult1_un124_sum_cry_3 ));
    InMux I__859 (
            .O(N__8763),
            .I(\RSMRST_PWRGD.un1_count_1_cry_2 ));
    InMux I__858 (
            .O(N__8760),
            .I(\RSMRST_PWRGD.un1_count_1_cry_3 ));
    InMux I__857 (
            .O(N__8757),
            .I(\RSMRST_PWRGD.un1_count_1_cry_4 ));
    InMux I__856 (
            .O(N__8754),
            .I(\RSMRST_PWRGD.un1_count_1_cry_5 ));
    InMux I__855 (
            .O(N__8751),
            .I(\RSMRST_PWRGD.un1_count_1_cry_6 ));
    InMux I__854 (
            .O(N__8748),
            .I(bfn_1_11_0_));
    InMux I__853 (
            .O(N__8745),
            .I(\RSMRST_PWRGD.un1_count_1_cry_8 ));
    InMux I__852 (
            .O(N__8742),
            .I(\RSMRST_PWRGD.un1_count_1_cry_9 ));
    InMux I__851 (
            .O(N__8739),
            .I(\RSMRST_PWRGD.un1_count_1_cry_10 ));
    CascadeMux I__850 (
            .O(N__8736),
            .I(N__8733));
    InMux I__849 (
            .O(N__8733),
            .I(N__8730));
    LocalMux I__848 (
            .O(N__8730),
            .I(\POWERLED.mult1_un152_sum_cry_5_s ));
    InMux I__847 (
            .O(N__8727),
            .I(\POWERLED.mult1_un159_sum_cry_4 ));
    InMux I__846 (
            .O(N__8724),
            .I(N__8721));
    LocalMux I__845 (
            .O(N__8721),
            .I(\POWERLED.mult1_un152_sum_cry_6_s ));
    CascadeMux I__844 (
            .O(N__8718),
            .I(N__8714));
    CascadeMux I__843 (
            .O(N__8717),
            .I(N__8710));
    InMux I__842 (
            .O(N__8714),
            .I(N__8703));
    InMux I__841 (
            .O(N__8713),
            .I(N__8703));
    InMux I__840 (
            .O(N__8710),
            .I(N__8703));
    LocalMux I__839 (
            .O(N__8703),
            .I(\POWERLED.mult1_un152_sum_i_0_8 ));
    InMux I__838 (
            .O(N__8700),
            .I(\POWERLED.mult1_un159_sum_cry_5 ));
    CascadeMux I__837 (
            .O(N__8697),
            .I(N__8694));
    InMux I__836 (
            .O(N__8694),
            .I(N__8691));
    LocalMux I__835 (
            .O(N__8691),
            .I(\POWERLED.mult1_un159_sum_axb_7 ));
    InMux I__834 (
            .O(N__8688),
            .I(\POWERLED.mult1_un159_sum_cry_6 ));
    CascadeMux I__833 (
            .O(N__8685),
            .I(\POWERLED.mult1_un159_sum_s_7_cascade_ ));
    InMux I__832 (
            .O(N__8682),
            .I(N__8679));
    LocalMux I__831 (
            .O(N__8679),
            .I(N__8676));
    Odrv12 I__830 (
            .O(N__8676),
            .I(\POWERLED.mult1_un145_sum_i ));
    InMux I__829 (
            .O(N__8673),
            .I(\RSMRST_PWRGD.un1_count_1_cry_0 ));
    InMux I__828 (
            .O(N__8670),
            .I(\RSMRST_PWRGD.un1_count_1_cry_1 ));
    CascadeMux I__827 (
            .O(N__8667),
            .I(N__8664));
    InMux I__826 (
            .O(N__8664),
            .I(N__8661));
    LocalMux I__825 (
            .O(N__8661),
            .I(\POWERLED.mult1_un145_sum_cry_5_s ));
    InMux I__824 (
            .O(N__8658),
            .I(\POWERLED.mult1_un152_sum_cry_5 ));
    InMux I__823 (
            .O(N__8655),
            .I(N__8652));
    LocalMux I__822 (
            .O(N__8652),
            .I(\POWERLED.mult1_un145_sum_cry_6_s ));
    CascadeMux I__821 (
            .O(N__8649),
            .I(N__8645));
    CascadeMux I__820 (
            .O(N__8648),
            .I(N__8641));
    InMux I__819 (
            .O(N__8645),
            .I(N__8634));
    InMux I__818 (
            .O(N__8644),
            .I(N__8634));
    InMux I__817 (
            .O(N__8641),
            .I(N__8634));
    LocalMux I__816 (
            .O(N__8634),
            .I(\POWERLED.mult1_un145_sum_i_0_8 ));
    InMux I__815 (
            .O(N__8631),
            .I(\POWERLED.mult1_un152_sum_cry_6 ));
    CascadeMux I__814 (
            .O(N__8628),
            .I(N__8625));
    InMux I__813 (
            .O(N__8625),
            .I(N__8622));
    LocalMux I__812 (
            .O(N__8622),
            .I(\POWERLED.mult1_un152_sum_axb_8 ));
    InMux I__811 (
            .O(N__8619),
            .I(\POWERLED.mult1_un152_sum_cry_7 ));
    CascadeMux I__810 (
            .O(N__8616),
            .I(\POWERLED.mult1_un152_sum_s_8_cascade_ ));
    InMux I__809 (
            .O(N__8613),
            .I(\POWERLED.mult1_un159_sum_cry_1 ));
    CascadeMux I__808 (
            .O(N__8610),
            .I(N__8607));
    InMux I__807 (
            .O(N__8607),
            .I(N__8604));
    LocalMux I__806 (
            .O(N__8604),
            .I(\POWERLED.mult1_un152_sum_cry_3_s ));
    InMux I__805 (
            .O(N__8601),
            .I(\POWERLED.mult1_un159_sum_cry_2 ));
    InMux I__804 (
            .O(N__8598),
            .I(N__8595));
    LocalMux I__803 (
            .O(N__8595),
            .I(\POWERLED.mult1_un152_sum_cry_4_s ));
    InMux I__802 (
            .O(N__8592),
            .I(\POWERLED.mult1_un159_sum_cry_3 ));
    InMux I__801 (
            .O(N__8589),
            .I(N__8586));
    LocalMux I__800 (
            .O(N__8586),
            .I(N__8583));
    Odrv4 I__799 (
            .O(N__8583),
            .I(\POWERLED.mult1_un138_sum_cry_4_s ));
    InMux I__798 (
            .O(N__8580),
            .I(\POWERLED.mult1_un145_sum_cry_4 ));
    CascadeMux I__797 (
            .O(N__8577),
            .I(N__8574));
    InMux I__796 (
            .O(N__8574),
            .I(N__8571));
    LocalMux I__795 (
            .O(N__8571),
            .I(N__8568));
    Odrv4 I__794 (
            .O(N__8568),
            .I(\POWERLED.mult1_un138_sum_cry_5_s ));
    InMux I__793 (
            .O(N__8565),
            .I(\POWERLED.mult1_un145_sum_cry_5 ));
    InMux I__792 (
            .O(N__8562),
            .I(N__8558));
    InMux I__791 (
            .O(N__8561),
            .I(N__8555));
    LocalMux I__790 (
            .O(N__8558),
            .I(N__8552));
    LocalMux I__789 (
            .O(N__8555),
            .I(\POWERLED.mult1_un138_sum_cry_6_s ));
    Odrv4 I__788 (
            .O(N__8552),
            .I(\POWERLED.mult1_un138_sum_cry_6_s ));
    CascadeMux I__787 (
            .O(N__8547),
            .I(N__8544));
    InMux I__786 (
            .O(N__8544),
            .I(N__8541));
    LocalMux I__785 (
            .O(N__8541),
            .I(\POWERLED.mult1_un145_sum_axb_7_l_fx ));
    InMux I__784 (
            .O(N__8538),
            .I(\POWERLED.mult1_un145_sum_cry_6 ));
    CascadeMux I__783 (
            .O(N__8535),
            .I(N__8532));
    InMux I__782 (
            .O(N__8532),
            .I(N__8529));
    LocalMux I__781 (
            .O(N__8529),
            .I(N__8526));
    Odrv4 I__780 (
            .O(N__8526),
            .I(\POWERLED.mult1_un145_sum_axb_8 ));
    InMux I__779 (
            .O(N__8523),
            .I(\POWERLED.mult1_un145_sum_cry_7 ));
    InMux I__778 (
            .O(N__8520),
            .I(\POWERLED.mult1_un152_sum_cry_2 ));
    CascadeMux I__777 (
            .O(N__8517),
            .I(N__8514));
    InMux I__776 (
            .O(N__8514),
            .I(N__8511));
    LocalMux I__775 (
            .O(N__8511),
            .I(\POWERLED.mult1_un145_sum_cry_3_s ));
    InMux I__774 (
            .O(N__8508),
            .I(\POWERLED.mult1_un152_sum_cry_3 ));
    InMux I__773 (
            .O(N__8505),
            .I(N__8502));
    LocalMux I__772 (
            .O(N__8502),
            .I(\POWERLED.mult1_un145_sum_cry_4_s ));
    InMux I__771 (
            .O(N__8499),
            .I(\POWERLED.mult1_un152_sum_cry_4 ));
    InMux I__770 (
            .O(N__8496),
            .I(N__8493));
    LocalMux I__769 (
            .O(N__8493),
            .I(\POWERLED.mult1_un131_sum_cry_6_s ));
    CascadeMux I__768 (
            .O(N__8490),
            .I(N__8486));
    CascadeMux I__767 (
            .O(N__8489),
            .I(N__8482));
    InMux I__766 (
            .O(N__8486),
            .I(N__8475));
    InMux I__765 (
            .O(N__8485),
            .I(N__8475));
    InMux I__764 (
            .O(N__8482),
            .I(N__8475));
    LocalMux I__763 (
            .O(N__8475),
            .I(\POWERLED.mult1_un131_sum_i_0_8 ));
    InMux I__762 (
            .O(N__8472),
            .I(\POWERLED.mult1_un138_sum_cry_6 ));
    CascadeMux I__761 (
            .O(N__8469),
            .I(N__8466));
    InMux I__760 (
            .O(N__8466),
            .I(N__8463));
    LocalMux I__759 (
            .O(N__8463),
            .I(\POWERLED.mult1_un138_sum_axb_8 ));
    InMux I__758 (
            .O(N__8460),
            .I(\POWERLED.mult1_un138_sum_cry_7 ));
    InMux I__757 (
            .O(N__8457),
            .I(N__8453));
    CascadeMux I__756 (
            .O(N__8456),
            .I(N__8449));
    LocalMux I__755 (
            .O(N__8453),
            .I(N__8445));
    InMux I__754 (
            .O(N__8452),
            .I(N__8440));
    InMux I__753 (
            .O(N__8449),
            .I(N__8440));
    InMux I__752 (
            .O(N__8448),
            .I(N__8437));
    Odrv4 I__751 (
            .O(N__8445),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__750 (
            .O(N__8440),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__749 (
            .O(N__8437),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    CascadeMux I__748 (
            .O(N__8430),
            .I(N__8427));
    InMux I__747 (
            .O(N__8427),
            .I(N__8424));
    LocalMux I__746 (
            .O(N__8424),
            .I(\POWERLED.mult1_un138_sum_i_0_8 ));
    InMux I__745 (
            .O(N__8421),
            .I(\POWERLED.mult1_un145_sum_cry_2 ));
    InMux I__744 (
            .O(N__8418),
            .I(N__8414));
    InMux I__743 (
            .O(N__8417),
            .I(N__8411));
    LocalMux I__742 (
            .O(N__8414),
            .I(N__8408));
    LocalMux I__741 (
            .O(N__8411),
            .I(\POWERLED.mult1_un138_sum_cry_3_s ));
    Odrv4 I__740 (
            .O(N__8408),
            .I(\POWERLED.mult1_un138_sum_cry_3_s ));
    CascadeMux I__739 (
            .O(N__8403),
            .I(N__8400));
    InMux I__738 (
            .O(N__8400),
            .I(N__8397));
    LocalMux I__737 (
            .O(N__8397),
            .I(\POWERLED.mult1_un145_sum_axb_4_l_fx ));
    InMux I__736 (
            .O(N__8394),
            .I(\POWERLED.mult1_un145_sum_cry_3 ));
    InMux I__735 (
            .O(N__8391),
            .I(\POWERLED.mult1_un131_sum_cry_5 ));
    InMux I__734 (
            .O(N__8388),
            .I(\POWERLED.mult1_un131_sum_cry_6 ));
    InMux I__733 (
            .O(N__8385),
            .I(\POWERLED.mult1_un131_sum_cry_7 ));
    CascadeMux I__732 (
            .O(N__8382),
            .I(\POWERLED.mult1_un131_sum_s_8_cascade_ ));
    InMux I__731 (
            .O(N__8379),
            .I(\POWERLED.mult1_un138_sum_cry_2 ));
    CascadeMux I__730 (
            .O(N__8376),
            .I(N__8373));
    InMux I__729 (
            .O(N__8373),
            .I(N__8370));
    LocalMux I__728 (
            .O(N__8370),
            .I(\POWERLED.mult1_un131_sum_cry_3_s ));
    InMux I__727 (
            .O(N__8367),
            .I(\POWERLED.mult1_un138_sum_cry_3 ));
    InMux I__726 (
            .O(N__8364),
            .I(N__8361));
    LocalMux I__725 (
            .O(N__8361),
            .I(\POWERLED.mult1_un131_sum_cry_4_s ));
    InMux I__724 (
            .O(N__8358),
            .I(\POWERLED.mult1_un138_sum_cry_4 ));
    CascadeMux I__723 (
            .O(N__8355),
            .I(N__8352));
    InMux I__722 (
            .O(N__8352),
            .I(N__8349));
    LocalMux I__721 (
            .O(N__8349),
            .I(\POWERLED.mult1_un131_sum_cry_5_s ));
    InMux I__720 (
            .O(N__8346),
            .I(\POWERLED.mult1_un138_sum_cry_5 ));
    InMux I__719 (
            .O(N__8343),
            .I(\POWERLED.mult1_un131_sum_cry_2 ));
    InMux I__718 (
            .O(N__8340),
            .I(\POWERLED.mult1_un131_sum_cry_3 ));
    InMux I__717 (
            .O(N__8337),
            .I(\POWERLED.mult1_un131_sum_cry_4 ));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(\POWERLED.dutycycle_cry_6 ),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(\POWERLED.dutycycle_cry_14 ),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_6_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_8_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_4_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_8_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_9_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_5_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_3_0_));
    defparam IN_MUX_bfv_1_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_2_0_));
    defparam IN_MUX_bfv_2_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_2_0_));
    defparam IN_MUX_bfv_4_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_5_0_));
    defparam IN_MUX_bfv_5_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_6_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\POWERLED.un1_count_off_1_cry_7 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(\POWERLED.un1_count_1_cry_8 ),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(\POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO ),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_9_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_4_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(\COUNTER.un4_counter_7 ),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(\COUNTER.counter_1_cry_8 ),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(\COUNTER.counter_1_cry_16 ),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(\COUNTER.counter_1_cry_24 ),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_7 ),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_2_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_5_0_));
    defparam IN_MUX_bfv_2_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_6_0_ (
            .carryinitin(\POWERLED.un1_count_2_cry_7 ),
            .carryinitout(bfn_2_6_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(\POWERLED.un1_count_2_cry_15 ),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_1_cry_7 ),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_1_cry_15 ),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\POWERLED.un1_count_clk_1_cry_7 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(\POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_1_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(\PCH_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(\PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(\ALL_SYS_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_11_9_0_));
    ICE_GB \COUNTER.tmp_RNIRH3P_0  (
            .USERSIGNALTOGLOBALBUFFER(N__10449),
            .GLOBALBUFFEROUTPUT(N_49_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_2_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_2_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_2_0  (
            .in0(_gnd_net_),
            .in1(N__10868),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_2_0_),
            .carryout(\POWERLED.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_2_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_2_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_2_1  (
            .in0(_gnd_net_),
            .in1(N__8841),
            .in2(N__8864),
            .in3(N__8343),
            .lcout(\POWERLED.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_2_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_2_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_2_2  (
            .in0(_gnd_net_),
            .in1(N__8860),
            .in2(N__8784),
            .in3(N__8340),
            .lcout(\POWERLED.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_2_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_2_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_2_3  (
            .in0(_gnd_net_),
            .in1(N__8772),
            .in2(N__9071),
            .in3(N__8337),
            .lcout(\POWERLED.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_2_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_2_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_2_4  (
            .in0(_gnd_net_),
            .in1(N__9067),
            .in2(N__8898),
            .in3(N__8391),
            .lcout(\POWERLED.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_2_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_2_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_2_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_2_5  (
            .in0(N__8448),
            .in1(N__8886),
            .in2(N__8865),
            .in3(N__8388),
            .lcout(\POWERLED.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_2_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_2_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_2_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_2_6  (
            .in0(_gnd_net_),
            .in1(N__8877),
            .in2(_gnd_net_),
            .in3(N__8385),
            .lcout(\POWERLED.mult1_un131_sum_s_8 ),
            .ltout(\POWERLED.mult1_un131_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_2_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_2_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_2_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8382),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_3_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_3_0  (
            .in0(_gnd_net_),
            .in1(N__10896),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(\POWERLED.mult1_un138_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_3_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_3_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_3_1  (
            .in0(_gnd_net_),
            .in1(N__8847),
            .in2(N__8489),
            .in3(N__8379),
            .lcout(\POWERLED.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_3_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_3_2  (
            .in0(_gnd_net_),
            .in1(N__8485),
            .in2(N__8376),
            .in3(N__8367),
            .lcout(\POWERLED.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_3_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_3_3  (
            .in0(_gnd_net_),
            .in1(N__8364),
            .in2(N__8456),
            .in3(N__8358),
            .lcout(\POWERLED.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_3_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_3_4  (
            .in0(_gnd_net_),
            .in1(N__8452),
            .in2(N__8355),
            .in3(N__8346),
            .lcout(\POWERLED.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_3_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_3_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_3_5  (
            .in0(N__9028),
            .in1(N__8496),
            .in2(N__8490),
            .in3(N__8472),
            .lcout(\POWERLED.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_3_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_3_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8469),
            .in3(N__8460),
            .lcout(\POWERLED.mult1_un138_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_4_l_fx_LC_1_4_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_4_l_fx_LC_1_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_4_l_fx_LC_1_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_4_l_fx_LC_1_4_1  (
            .in0(N__8417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9026),
            .lcout(\POWERLED.mult1_un145_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_1_4_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_1_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_1_4_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_1_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8457),
            .lcout(\POWERLED.un1_count_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_4_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_4_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9025),
            .lcout(\POWERLED.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_7_l_fx_LC_1_4_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_7_l_fx_LC_1_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_7_l_fx_LC_1_4_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_7_l_fx_LC_1_4_7  (
            .in0(N__8561),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9027),
            .lcout(\POWERLED.mult1_un145_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_1_5_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_1_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10917),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_5_0_),
            .carryout(\POWERLED.mult1_un145_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_1_5_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_1_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_1_5_1  (
            .in0(_gnd_net_),
            .in1(N__9324),
            .in2(N__8430),
            .in3(N__8421),
            .lcout(\POWERLED.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_1_5_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_1_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_1_5_2  (
            .in0(_gnd_net_),
            .in1(N__8418),
            .in2(N__8403),
            .in3(N__8394),
            .lcout(\POWERLED.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_1_5_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_1_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_1_5_3  (
            .in0(_gnd_net_),
            .in1(N__8589),
            .in2(N__9039),
            .in3(N__8580),
            .lcout(\POWERLED.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_1_5_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_1_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(N__9038),
            .in2(N__8577),
            .in3(N__8565),
            .lcout(\POWERLED.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_1_5_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_1_5_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_1_5_5  (
            .in0(N__8994),
            .in1(N__8562),
            .in2(N__8547),
            .in3(N__8538),
            .lcout(\POWERLED.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_1_5_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_1_5_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_1_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8535),
            .in3(N__8523),
            .lcout(\POWERLED.mult1_un145_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_1_5_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_1_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_1_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8993),
            .lcout(\POWERLED.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_1_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_1_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__14102),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(\POWERLED.mult1_un152_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_1_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_1_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__8682),
            .in2(N__8648),
            .in3(N__8520),
            .lcout(\POWERLED.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_1_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_1_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(N__8644),
            .in2(N__8517),
            .in3(N__8508),
            .lcout(\POWERLED.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_1_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_1_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(N__8505),
            .in2(N__9000),
            .in3(N__8499),
            .lcout(\POWERLED.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_1_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_1_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(N__8998),
            .in2(N__8667),
            .in3(N__8658),
            .lcout(\POWERLED.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_1_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_1_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_1_6_5  (
            .in0(N__9195),
            .in1(N__8655),
            .in2(N__8649),
            .in3(N__8631),
            .lcout(\POWERLED.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_1_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_1_6_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8628),
            .in3(N__8619),
            .lcout(\POWERLED.mult1_un152_sum_s_8 ),
            .ltout(\POWERLED.mult1_un152_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_1_6_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_1_6_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8616),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_1_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_1_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__14652),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(\POWERLED.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_1_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_1_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(N__9207),
            .in2(N__8717),
            .in3(N__8613),
            .lcout(\POWERLED.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_1_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_1_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_1_7_2  (
            .in0(_gnd_net_),
            .in1(N__8713),
            .in2(N__8610),
            .in3(N__8601),
            .lcout(\POWERLED.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_1_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_1_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_1_7_3  (
            .in0(_gnd_net_),
            .in1(N__8598),
            .in2(N__9201),
            .in3(N__8592),
            .lcout(\POWERLED.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_1_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_1_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_1_7_4  (
            .in0(_gnd_net_),
            .in1(N__9199),
            .in2(N__8736),
            .in3(N__8727),
            .lcout(\POWERLED.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_1_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_1_7_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_1_7_5  (
            .in0(N__9419),
            .in1(N__8724),
            .in2(N__8718),
            .in3(N__8700),
            .lcout(\POWERLED.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_1_7_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_1_7_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_1_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8697),
            .in3(N__8688),
            .lcout(\POWERLED.mult1_un159_sum_s_7 ),
            .ltout(\POWERLED.mult1_un159_sum_s_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_1_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_1_7_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_1_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8685),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_0_LC_1_8_3 .C_ON=1'b0;
    defparam \POWERLED.curr_state_0_LC_1_8_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.curr_state_0_LC_1_8_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \POWERLED.curr_state_0_LC_1_8_3  (
            .in0(_gnd_net_),
            .in1(N__10129),
            .in2(N__9459),
            .in3(N__10356),
            .lcout(\POWERLED.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19243),
            .ce(N__18491),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_1_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_1_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10916),
            .lcout(\POWERLED.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_0_LC_1_10_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_0_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_0_LC_1_10_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_0_LC_1_10_0  (
            .in0(N__18837),
            .in1(N__9471),
            .in2(N__9705),
            .in3(N__9704),
            .lcout(\RSMRST_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .clk(N__19244),
            .ce(),
            .sr(N__9813));
    defparam \RSMRST_PWRGD.count_1_LC_1_10_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_1_LC_1_10_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_1_LC_1_10_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_1_LC_1_10_1  (
            .in0(N__18833),
            .in1(N__9630),
            .in2(_gnd_net_),
            .in3(N__8673),
            .lcout(\RSMRST_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .clk(N__19244),
            .ce(),
            .sr(N__9813));
    defparam \RSMRST_PWRGD.count_2_LC_1_10_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_2_LC_1_10_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_2_LC_1_10_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_2_LC_1_10_2  (
            .in0(N__18838),
            .in1(N__9603),
            .in2(_gnd_net_),
            .in3(N__8670),
            .lcout(\RSMRST_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .clk(N__19244),
            .ce(),
            .sr(N__9813));
    defparam \RSMRST_PWRGD.count_3_LC_1_10_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_3_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_3_LC_1_10_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_3_LC_1_10_3  (
            .in0(N__18834),
            .in1(N__9678),
            .in2(_gnd_net_),
            .in3(N__8763),
            .lcout(\RSMRST_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .clk(N__19244),
            .ce(),
            .sr(N__9813));
    defparam \RSMRST_PWRGD.count_4_LC_1_10_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_4_LC_1_10_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_4_LC_1_10_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_4_LC_1_10_4  (
            .in0(N__18839),
            .in1(N__9642),
            .in2(_gnd_net_),
            .in3(N__8760),
            .lcout(\RSMRST_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .clk(N__19244),
            .ce(),
            .sr(N__9813));
    defparam \RSMRST_PWRGD.count_5_LC_1_10_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_5_LC_1_10_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_5_LC_1_10_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_5_LC_1_10_5  (
            .in0(N__18835),
            .in1(N__9617),
            .in2(_gnd_net_),
            .in3(N__8757),
            .lcout(\RSMRST_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .clk(N__19244),
            .ce(),
            .sr(N__9813));
    defparam \RSMRST_PWRGD.count_6_LC_1_10_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_6_LC_1_10_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_6_LC_1_10_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_6_LC_1_10_6  (
            .in0(N__18840),
            .in1(N__9552),
            .in2(_gnd_net_),
            .in3(N__8754),
            .lcout(\RSMRST_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .clk(N__19244),
            .ce(),
            .sr(N__9813));
    defparam \RSMRST_PWRGD.count_7_LC_1_10_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_7_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_7_LC_1_10_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_7_LC_1_10_7  (
            .in0(N__18836),
            .in1(N__9690),
            .in2(_gnd_net_),
            .in3(N__8751),
            .lcout(\RSMRST_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .clk(N__19244),
            .ce(),
            .sr(N__9813));
    defparam \RSMRST_PWRGD.count_8_LC_1_11_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_8_LC_1_11_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_8_LC_1_11_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_8_LC_1_11_0  (
            .in0(N__18832),
            .in1(N__9498),
            .in2(_gnd_net_),
            .in3(N__8748),
            .lcout(\RSMRST_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .clk(N__19231),
            .ce(),
            .sr(N__9812));
    defparam \RSMRST_PWRGD.count_9_LC_1_11_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_9_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_9_LC_1_11_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_9_LC_1_11_1  (
            .in0(N__18798),
            .in1(N__9510),
            .in2(_gnd_net_),
            .in3(N__8745),
            .lcout(\RSMRST_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .clk(N__19231),
            .ce(),
            .sr(N__9812));
    defparam \RSMRST_PWRGD.count_10_LC_1_11_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_10_LC_1_11_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_10_LC_1_11_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_10_LC_1_11_2  (
            .in0(N__18829),
            .in1(N__9591),
            .in2(_gnd_net_),
            .in3(N__8742),
            .lcout(\RSMRST_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .clk(N__19231),
            .ce(),
            .sr(N__9812));
    defparam \RSMRST_PWRGD.count_11_LC_1_11_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_11_LC_1_11_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_11_LC_1_11_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_11_LC_1_11_3  (
            .in0(N__18796),
            .in1(N__9579),
            .in2(_gnd_net_),
            .in3(N__8739),
            .lcout(\RSMRST_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .clk(N__19231),
            .ce(),
            .sr(N__9812));
    defparam \RSMRST_PWRGD.count_12_LC_1_11_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_12_LC_1_11_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_12_LC_1_11_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_12_LC_1_11_4  (
            .in0(N__18830),
            .in1(N__9485),
            .in2(_gnd_net_),
            .in3(N__8811),
            .lcout(\RSMRST_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .clk(N__19231),
            .ce(),
            .sr(N__9812));
    defparam \RSMRST_PWRGD.count_13_LC_1_11_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_13_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_13_LC_1_11_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_13_LC_1_11_5  (
            .in0(N__18797),
            .in1(N__9566),
            .in2(_gnd_net_),
            .in3(N__8808),
            .lcout(\RSMRST_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .clk(N__19231),
            .ce(),
            .sr(N__9812));
    defparam \RSMRST_PWRGD.count_14_LC_1_11_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_14_LC_1_11_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_14_LC_1_11_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_14_LC_1_11_6  (
            .in0(N__18831),
            .in1(N__9528),
            .in2(_gnd_net_),
            .in3(N__8805),
            .lcout(\RSMRST_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .clk(N__19231),
            .ce(),
            .sr(N__9812));
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_11_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__17298),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_15_LC_1_12_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_15_LC_1_12_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_esr_15_LC_1_12_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \RSMRST_PWRGD.count_esr_15_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__9540),
            .in2(_gnd_net_),
            .in3(N__8802),
            .lcout(\RSMRST_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19248),
            .ce(N__9777),
            .sr(N__9805));
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_13_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_13_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \VPP_VDDQ.un1_vddq_en_LC_1_13_7  (
            .in0(N__17674),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8799),
            .lcout(vddq_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_2_2_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_2_2_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_2_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_2_2_0  (
            .in0(_gnd_net_),
            .in1(N__10835),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_2_0_),
            .carryout(\POWERLED.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_2_2_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_2_2_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_2_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_2_2_1  (
            .in0(_gnd_net_),
            .in1(N__8817),
            .in2(N__8834),
            .in3(N__8775),
            .lcout(\POWERLED.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_2_2_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_2_2_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_2_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_2_2_2  (
            .in0(_gnd_net_),
            .in1(N__8830),
            .in2(N__9918),
            .in3(N__8766),
            .lcout(\POWERLED.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_2_2_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_2_2_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_2_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_2_2_3  (
            .in0(_gnd_net_),
            .in1(N__9900),
            .in2(N__10056),
            .in3(N__8889),
            .lcout(\POWERLED.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_2_2_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_2_2_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_2_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_2_2_4  (
            .in0(_gnd_net_),
            .in1(N__10055),
            .in2(N__9885),
            .in3(N__8880),
            .lcout(\POWERLED.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_2_2_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_2_2_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_2_2_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_2_2_5  (
            .in0(N__9063),
            .in1(N__9867),
            .in2(N__8835),
            .in3(N__8871),
            .lcout(\POWERLED.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_2_2_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_2_2_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_2_2_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_2_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9852),
            .in3(N__8868),
            .lcout(\POWERLED.mult1_un124_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_2_2_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_2_2_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_2_2_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_2_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9062),
            .lcout(\POWERLED.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_3_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_3_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_3_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10869),
            .lcout(\POWERLED.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_2_3_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_2_3_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_2_3_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_2_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10836),
            .lcout(\POWERLED.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_2_3_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_2_3_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_2_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10051),
            .lcout(\POWERLED.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_2_3_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_2_3_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_2_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10803),
            .lcout(\POWERLED.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_2_4_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_2_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_2_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9072),
            .lcout(\POWERLED.un1_count_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_2_4_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_2_4_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_2_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9034),
            .lcout(\POWERLED.un1_count_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_2_4_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_2_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_2_4_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_2_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8999),
            .lcout(\POWERLED.un1_count_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_0_c_inv_LC_2_5_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_0_c_inv_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_0_c_inv_LC_2_5_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_0_c_inv_LC_2_5_0  (
            .in0(_gnd_net_),
            .in1(N__8970),
            .in2(N__9363),
            .in3(N__11384),
            .lcout(\POWERLED.count_i_0_0 ),
            .ltout(),
            .carryin(bfn_2_5_0_),
            .carryout(\POWERLED.un1_count_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_1_c_inv_LC_2_5_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_1_c_inv_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_1_c_inv_LC_2_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_1_c_inv_LC_2_5_1  (
            .in0(_gnd_net_),
            .in1(N__8946),
            .in2(N__8958),
            .in3(N__11412),
            .lcout(\POWERLED.count_i_1 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_0 ),
            .carryout(\POWERLED.un1_count_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_2_c_inv_LC_2_5_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_2_c_inv_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_2_c_inv_LC_2_5_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_2_c_inv_LC_2_5_2  (
            .in0(_gnd_net_),
            .in1(N__9177),
            .in2(N__8940),
            .in3(N__11348),
            .lcout(\POWERLED.count_i_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_1 ),
            .carryout(\POWERLED.un1_count_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_3_c_inv_LC_2_5_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_3_c_inv_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_3_c_inv_LC_2_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_3_c_inv_LC_2_5_3  (
            .in0(_gnd_net_),
            .in1(N__8931),
            .in2(N__8925),
            .in3(N__11309),
            .lcout(\POWERLED.count_i_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_2 ),
            .carryout(\POWERLED.un1_count_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_4_c_inv_LC_2_5_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_4_c_inv_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_4_c_inv_LC_2_5_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_4_c_inv_LC_2_5_4  (
            .in0(_gnd_net_),
            .in1(N__8913),
            .in2(N__8907),
            .in3(N__11783),
            .lcout(\POWERLED.count_i_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_3 ),
            .carryout(\POWERLED.un1_count_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_5_c_inv_LC_2_5_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_5_c_inv_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_5_c_inv_LC_2_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_5_c_inv_LC_2_5_5  (
            .in0(_gnd_net_),
            .in1(N__9153),
            .in2(N__9162),
            .in3(N__11744),
            .lcout(\POWERLED.count_i_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_4 ),
            .carryout(\POWERLED.un1_count_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_6_c_inv_LC_2_5_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_6_c_inv_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_6_c_inv_LC_2_5_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_6_c_inv_LC_2_5_6  (
            .in0(_gnd_net_),
            .in1(N__9147),
            .in2(N__9141),
            .in3(N__11706),
            .lcout(\POWERLED.count_i_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_5 ),
            .carryout(\POWERLED.un1_count_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_7_c_inv_LC_2_5_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_7_c_inv_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_7_c_inv_LC_2_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_7_c_inv_LC_2_5_7  (
            .in0(_gnd_net_),
            .in1(N__10017),
            .in2(N__9132),
            .in3(N__11663),
            .lcout(\POWERLED.count_i_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_6 ),
            .carryout(\POWERLED.un1_count_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_8_c_inv_LC_2_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_8_c_inv_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_8_c_inv_LC_2_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_8_c_inv_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(N__9990),
            .in2(N__9123),
            .in3(N__11624),
            .lcout(\POWERLED.count_i_8 ),
            .ltout(),
            .carryin(bfn_2_6_0_),
            .carryout(\POWERLED.un1_count_2_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_9_c_inv_LC_2_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_9_c_inv_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_9_c_inv_LC_2_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_9_c_inv_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(N__9999),
            .in2(N__9114),
            .in3(N__11586),
            .lcout(\POWERLED.count_i_9 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_8 ),
            .carryout(\POWERLED.un1_count_2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_10_c_inv_LC_2_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_10_c_inv_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_10_c_inv_LC_2_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_10_c_inv_LC_2_6_2  (
            .in0(_gnd_net_),
            .in1(N__9951),
            .in2(N__9105),
            .in3(N__11550),
            .lcout(\POWERLED.count_i_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_9 ),
            .carryout(\POWERLED.un1_count_2_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_11_c_inv_LC_2_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_11_c_inv_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_11_c_inv_LC_2_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_11_c_inv_LC_2_6_3  (
            .in0(_gnd_net_),
            .in1(N__9942),
            .in2(N__9096),
            .in3(N__11508),
            .lcout(\POWERLED.count_i_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_10 ),
            .carryout(\POWERLED.un1_count_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_12_c_inv_LC_2_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_12_c_inv_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_12_c_inv_LC_2_6_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_count_2_cry_12_c_inv_LC_2_6_4  (
            .in0(N__12045),
            .in1(N__9168),
            .in2(N__9087),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_i_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_11 ),
            .carryout(\POWERLED.un1_count_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_13_c_inv_LC_2_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_13_c_inv_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_13_c_inv_LC_2_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_13_c_inv_LC_2_6_5  (
            .in0(_gnd_net_),
            .in1(N__9078),
            .in2(N__9963),
            .in3(N__12012),
            .lcout(\POWERLED.count_i_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_12 ),
            .carryout(\POWERLED.un1_count_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_14_c_inv_LC_2_6_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_14_c_inv_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_14_c_inv_LC_2_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_14_c_inv_LC_2_6_6  (
            .in0(_gnd_net_),
            .in1(N__10008),
            .in2(N__9345),
            .in3(N__11976),
            .lcout(\POWERLED.count_i_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_13 ),
            .carryout(\POWERLED.un1_count_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_15_c_inv_LC_2_6_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_15_c_inv_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_15_c_inv_LC_2_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_15_c_inv_LC_2_6_7  (
            .in0(_gnd_net_),
            .in1(N__10212),
            .in2(N__9336),
            .in3(N__11933),
            .lcout(\POWERLED.count_i_15 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_14 ),
            .carryout(\POWERLED.un1_count_2_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_2_7_0 .C_ON=1'b0;
    defparam \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_2_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_2_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9327),
            .lcout(\POWERLED.un1_count_2_cry_15_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_2_7_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_2_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10895),
            .lcout(\POWERLED.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_2_7_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_2_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_2_7_2  (
            .in0(N__9315),
            .in1(N__9270),
            .in2(N__9258),
            .in3(N__9230),
            .lcout(rsmrst_pwrgd_signal),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_2_7_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_2_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_2_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14103),
            .lcout(\POWERLED.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_2_7_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_2_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_2_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9200),
            .lcout(\POWERLED.un1_count_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_7_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12456),
            .lcout(\POWERLED.un1_count_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_LC_2_7_6 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_LC_2_7_6 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \POWERLED.pwm_out_RNO_LC_2_7_6  (
            .in0(N__9717),
            .in1(N__10448),
            .in2(N__10135),
            .in3(N__9455),
            .lcout(\POWERLED.pwm_out_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_2_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_2_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(N__14547),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(\POWERLED.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_2_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_2_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_2_8_1  (
            .in0(_gnd_net_),
            .in1(N__9351),
            .in2(N__9392),
            .in3(N__9414),
            .lcout(G_385),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_0 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_2_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_2_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(N__9388),
            .in2(N__9444),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_2_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_2_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_2_8_3  (
            .in0(_gnd_net_),
            .in1(N__9415),
            .in2(N__9435),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_2_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_2_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__9426),
            .in2(N__9420),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_2_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_2_8_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(N__9399),
            .in2(N__9393),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_2_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_2_8_6 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9375),
            .in3(N__9366),
            .lcout(\POWERLED.un1_count_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_2_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_2_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_2_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14651),
            .lcout(\POWERLED.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_1_LC_2_9_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_1_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_1_LC_2_9_0 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \RSMRST_PWRGD.curr_state_1_LC_2_9_0  (
            .in0(N__10276),
            .in1(N__18069),
            .in2(N__9666),
            .in3(N__9743),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19170),
            .ce(N__18475),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_2_10_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_2_10_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_2_10_0  (
            .in0(N__9661),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18070),
            .lcout(\RSMRST_PWRGD.N_240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_2_10_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_2_10_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_2_10_1  (
            .in0(N__18071),
            .in1(N__9660),
            .in2(_gnd_net_),
            .in3(N__10275),
            .lcout(\RSMRST_PWRGD.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_12_LC_2_10_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_12_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_12_LC_2_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_12_LC_2_10_2  (
            .in0(N__9689),
            .in1(N__9677),
            .in2(N__9665),
            .in3(N__9516),
            .lcout(\RSMRST_PWRGD.m4_i_i_a2_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_10_LC_2_10_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_10_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_10_LC_2_10_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_10_LC_2_10_6  (
            .in0(N__9641),
            .in1(N__9629),
            .in2(N__9618),
            .in3(N__9602),
            .lcout(\RSMRST_PWRGD.m4_i_i_a2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_11_LC_2_11_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_11_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_11_LC_2_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_11_LC_2_11_2  (
            .in0(N__9590),
            .in1(N__9578),
            .in2(N__9567),
            .in3(N__9551),
            .lcout(\RSMRST_PWRGD.m4_i_i_a2_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_7_LC_2_11_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_7_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_7_LC_2_11_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_7_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__9539),
            .in2(_gnd_net_),
            .in3(N__9527),
            .lcout(\RSMRST_PWRGD.m4_i_i_a2_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_9_LC_2_11_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_9_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_9_LC_2_11_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_9_LC_2_11_5  (
            .in0(N__9509),
            .in1(N__9497),
            .in2(N__9486),
            .in3(N__9470),
            .lcout(),
            .ltout(\RSMRST_PWRGD.m4_i_i_a2_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_LC_2_11_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_LC_2_11_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_LC_2_11_6  (
            .in0(N__9834),
            .in1(N__9828),
            .in2(N__9822),
            .in3(N__9819),
            .lcout(\RSMRST_PWRGD.N_241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNIJULM7_0_LC_2_12_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNIJULM7_0_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNIJULM7_0_LC_2_12_3 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNIJULM7_0_LC_2_12_3  (
            .in0(N__10234),
            .in1(N__9736),
            .in2(N__10277),
            .in3(N__18755),
            .lcout(\RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0 ),
            .ltout(\RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_2_12_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_2_12_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \RSMRST_PWRGD.count_esr_RNO_0_15_LC_2_12_4  (
            .in0(N__18756),
            .in1(_gnd_net_),
            .in2(N__9780),
            .in3(_gnd_net_),
            .lcout(\RSMRST_PWRGD.N_49_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_EN_i_i_i_LC_2_12_5 .C_ON=1'b0;
    defparam \POWERLED.VCCST_EN_i_i_i_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_EN_i_i_i_LC_2_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.VCCST_EN_i_i_i_LC_2_12_5  (
            .in0(N__16782),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(v5s_enn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_0_LC_2_13_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_0_LC_2_13_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_0_LC_2_13_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \RSMRST_PWRGD.curr_state_0_LC_2_13_6  (
            .in0(N__10274),
            .in1(N__10238),
            .in2(_gnd_net_),
            .in3(N__9744),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19213),
            .ce(N__18487),
            .sr(_gnd_net_));
    defparam \POWERLED.count_0_LC_4_3_1 .C_ON=1'b0;
    defparam \POWERLED.count_0_LC_4_3_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_0_LC_4_3_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.count_0_LC_4_3_1  (
            .in0(_gnd_net_),
            .in1(N__11382),
            .in2(_gnd_net_),
            .in3(N__18779),
            .lcout(\POWERLED.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19067),
            .ce(),
            .sr(N__11867));
    defparam \POWERLED.pwm_out_RNO_4_LC_4_4_0 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_4_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_4_LC_4_4_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.pwm_out_RNO_4_LC_4_4_0  (
            .in0(N__11784),
            .in1(N__11310),
            .in2(_gnd_net_),
            .in3(N__11349),
            .lcout(\POWERLED.un1_countlt6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_1_LC_4_4_1 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_1_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_1_LC_4_4_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.pwm_out_RNO_1_LC_4_4_1  (
            .in0(N__12044),
            .in1(N__11507),
            .in2(_gnd_net_),
            .in3(N__11625),
            .lcout(),
            .ltout(\POWERLED.g0_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_0_LC_4_4_2 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_0_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_0_LC_4_4_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \POWERLED.pwm_out_RNO_0_LC_4_4_2  (
            .in0(N__9924),
            .in1(N__11546),
            .in2(N__9720),
            .in3(N__11664),
            .lcout(\POWERLED.un1_count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNI75RB5_0_LC_4_4_4 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI75RB5_0_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI75RB5_0_LC_4_4_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \POWERLED.curr_state_RNI75RB5_0_LC_4_4_4  (
            .in0(N__10142),
            .in1(N__10346),
            .in2(_gnd_net_),
            .in3(N__18739),
            .lcout(\POWERLED.curr_state_RNI75RB5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_3_LC_4_4_5 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_3_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_3_LC_4_4_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.pwm_out_RNO_3_LC_4_4_5  (
            .in0(N__12011),
            .in1(N__11585),
            .in2(N__11934),
            .in3(N__11972),
            .lcout(),
            .ltout(\POWERLED.g0_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_2_LC_4_4_6 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_2_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_2_LC_4_4_6 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \POWERLED.pwm_out_RNO_2_LC_4_4_6  (
            .in0(N__9933),
            .in1(N__11705),
            .in2(N__9927),
            .in3(N__11745),
            .lcout(\POWERLED.g0_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_5_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_5_0  (
            .in0(_gnd_net_),
            .in1(N__10802),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_5_0_),
            .carryout(\POWERLED.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_5_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_5_1  (
            .in0(_gnd_net_),
            .in1(N__10425),
            .in2(N__9980),
            .in3(N__9903),
            .lcout(\POWERLED.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_5_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_5_2  (
            .in0(_gnd_net_),
            .in1(N__9976),
            .in2(N__10410),
            .in3(N__9888),
            .lcout(\POWERLED.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_5_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(N__10398),
            .in2(N__10509),
            .in3(N__9870),
            .lcout(\POWERLED.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_5_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(N__10508),
            .in2(N__10389),
            .in3(N__9855),
            .lcout(\POWERLED.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_5_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_5_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_5_5  (
            .in0(N__10039),
            .in1(N__10530),
            .in2(N__9981),
            .in3(N__9837),
            .lcout(\POWERLED.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_5_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_5_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_5_6  (
            .in0(_gnd_net_),
            .in1(N__10521),
            .in2(_gnd_net_),
            .in3(N__10059),
            .lcout(\POWERLED.mult1_un117_sum_s_8 ),
            .ltout(\POWERLED.mult1_un117_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_5_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_5_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10020),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_6_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12666),
            .lcout(\POWERLED.un1_count_2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_4_6_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_4_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12114),
            .lcout(\POWERLED.un1_count_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_6_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_6_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_6_3  (
            .in0(N__10503),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_6_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10502),
            .lcout(\POWERLED.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_4_6_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_4_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_4_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12570),
            .lcout(\POWERLED.un1_count_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_4_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_4_6_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_4_6_6  (
            .in0(N__12200),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_6_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12303),
            .lcout(\POWERLED.un1_count_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_7_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12405),
            .lcout(\POWERLED.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_LC_4_7_7 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_LC_4_7_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.pwm_out_LC_4_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.pwm_out_LC_4_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10146),
            .lcout(pwrbtn_led),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19138),
            .ce(N__10089),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10977),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_8_0_),
            .carryout(\POWERLED.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_8_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10317),
            .in3(N__10077),
            .lcout(\POWERLED.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_8_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10200),
            .in3(N__10074),
            .lcout(\POWERLED.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_8_3  (
            .in0(_gnd_net_),
            .in1(N__17260),
            .in2(N__10188),
            .in3(N__10071),
            .lcout(\POWERLED.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(N__17266),
            .in2(N__10176),
            .in3(N__10068),
            .lcout(\POWERLED.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_4_8_5 .C_ON=1'b1;
    defparam \POWERLED.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_4_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10749),
            .in3(N__10065),
            .lcout(\POWERLED.mult1_un54_sum_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_4_8_6 .C_ON=1'b0;
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_4_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_4_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10062),
            .lcout(\POWERLED.mult1_un54_sum_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10670),
            .lcout(\POWERLED.un1_count_2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10956),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(\POWERLED.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_9_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10326),
            .in3(N__10191),
            .lcout(\POWERLED.mult1_un47_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_9_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10305),
            .in3(N__10179),
            .lcout(\POWERLED.mult1_un47_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__11064),
            .in2(N__17299),
            .in3(N__10167),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_4_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_4_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(N__17288),
            .in2(N__10293),
            .in3(N__10164),
            .lcout(\POWERLED.mult1_un47_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_9_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_9_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10161),
            .in3(N__10152),
            .lcout(\POWERLED.mult1_un54_sum_s_8 ),
            .ltout(\POWERLED.mult1_un54_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_9_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10149),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_9_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_9_7  (
            .in0(N__10976),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un54_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_4_10_0 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_4_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_4_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11109),
            .lcout(\POWERLED.un1_dutycycle_1_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_4_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_4_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_4_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10952),
            .lcout(\POWERLED.un1_dutycycle_1_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_4_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_4_10_7 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_4_10_7  (
            .in0(N__11110),
            .in1(_gnd_net_),
            .in2(N__11088),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_EN_i_i_0_a2_LC_4_11_2 .C_ON=1'b0;
    defparam \POWERLED.VCCST_EN_i_i_0_a2_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_EN_i_i_0_a2_LC_4_11_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.VCCST_EN_i_i_0_a2_LC_4_11_2  (
            .in0(N__16536),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14683),
            .lcout(vccst_en),
            .ltout(vccst_en_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_1_sqmuxa_5_0_a2_LC_4_11_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_1_sqmuxa_5_0_a2_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_1_sqmuxa_5_0_a2_LC_4_11_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \POWERLED.count_clk_1_sqmuxa_5_0_a2_LC_4_11_3  (
            .in0(N__16435),
            .in1(_gnd_net_),
            .in2(N__10296),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_4_11_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_4_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10994),
            .lcout(\POWERLED.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_4_11_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_4_11_5 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(N__11121),
            .in2(N__11115),
            .in3(N__11084),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_LC_4_12_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_LC_4_12_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_LC_4_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(N__10281),
            .in2(_gnd_net_),
            .in3(N__10239),
            .lcout(rsmrstn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19224),
            .ce(N__18486),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI63141_10_LC_4_13_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_4_13_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_RNI63141_10_LC_4_13_5  (
            .in0(N__11225),
            .in1(N__11027),
            .in2(N__11163),
            .in3(N__11042),
            .lcout(\VPP_VDDQ.un6_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_4_13_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_4_13_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_RNIVJP51_3_LC_4_13_7  (
            .in0(N__11240),
            .in1(N__11255),
            .in2(N__11211),
            .in3(N__11270),
            .lcout(\VPP_VDDQ.un6_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_4_14_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_4_14_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \VPP_VDDQ.count_RNIFC141_11_LC_4_14_3  (
            .in0(N__11177),
            .in1(N__11054),
            .in2(N__11145),
            .in3(N__11192),
            .lcout(),
            .ltout(\VPP_VDDQ.un6_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_4_14_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_4_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_esr_RNIRFM64_15_LC_4_14_4  (
            .in0(N__10362),
            .in1(N__10377),
            .in2(N__10371),
            .in3(N__10368),
            .lcout(\VPP_VDDQ.count_esr_RNIRFM64Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_4_14_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_4_14_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_esr_RNI7CQO_15_LC_4_14_5  (
            .in0(N__11444),
            .in1(N__11459),
            .in2(N__11427),
            .in3(N__11474),
            .lcout(\VPP_VDDQ.un6_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_1_LC_5_3_3 .C_ON=1'b0;
    defparam \POWERLED.count_1_LC_5_3_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_1_LC_5_3_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \POWERLED.count_1_LC_5_3_3  (
            .in0(N__11405),
            .in1(N__11383),
            .in2(_gnd_net_),
            .in3(N__18780),
            .lcout(\POWERLED.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19066),
            .ce(),
            .sr(N__11871));
    defparam \POWERLED.count_RNIOVT24_11_LC_5_4_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNIOVT24_11_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIOVT24_11_LC_5_4_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.count_RNIOVT24_11_LC_5_4_1  (
            .in0(N__12039),
            .in1(N__11502),
            .in2(N__10335),
            .in3(N__10455),
            .lcout(\POWERLED.count_RNIOVT24Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNID4E61_7_LC_5_4_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNID4E61_7_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNID4E61_7_LC_5_4_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_RNID4E61_7_LC_5_4_2  (
            .in0(N__11574),
            .in1(N__11610),
            .in2(N__11542),
            .in3(N__11649),
            .lcout(\POWERLED.un1_countlto15_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_esr_RNIBHMO_15_LC_5_4_4 .C_ON=1'b0;
    defparam \POWERLED.count_esr_RNIBHMO_15_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_esr_RNIBHMO_15_LC_5_4_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.count_esr_RNIBHMO_15_LC_5_4_4  (
            .in0(N__11932),
            .in1(N__11964),
            .in2(_gnd_net_),
            .in3(N__12003),
            .lcout(\POWERLED.un1_countlto15_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNICO6R_2_LC_5_4_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNICO6R_2_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNICO6R_2_LC_5_4_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.count_RNICO6R_2_LC_5_4_6  (
            .in0(N__11769),
            .in1(N__11334),
            .in2(_gnd_net_),
            .in3(N__11295),
            .lcout(),
            .ltout(\POWERLED.un1_countlt6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI6IPJ2_5_LC_5_4_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNI6IPJ2_5_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI6IPJ2_5_LC_5_4_7 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \POWERLED.count_RNI6IPJ2_5_LC_5_4_7  (
            .in0(N__11694),
            .in1(N__11733),
            .in2(N__10464),
            .in3(N__10461),
            .lcout(\POWERLED.un1_countlto15_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_esr_RNO_0_15_LC_5_5_1 .C_ON=1'b0;
    defparam \POWERLED.count_esr_RNO_0_15_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_esr_RNO_0_15_LC_5_5_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.count_esr_RNO_0_15_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(N__18742),
            .in2(_gnd_net_),
            .in3(N__11866),
            .lcout(\POWERLED.N_49_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_RNIRH3P_LC_5_5_2 .C_ON=1'b0;
    defparam \COUNTER.tmp_RNIRH3P_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_RNIRH3P_LC_5_5_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \COUNTER.tmp_RNIRH3P_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(N__10418),
            .in2(_gnd_net_),
            .in3(N__15779),
            .lcout(tmp_RNIRH3P),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_5_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10770),
            .lcout(\POWERLED.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_LC_5_5_6 .C_ON=1'b0;
    defparam \COUNTER.tmp_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_LC_5_5_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.tmp_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(N__10419),
            .in2(_gnd_net_),
            .in3(N__15780),
            .lcout(\COUNTER.tmp_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19137),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(N__10769),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_6_0_),
            .carryout(\POWERLED.mult1_un110_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_6_1  (
            .in0(_gnd_net_),
            .in1(N__10482),
            .in2(N__12083),
            .in3(N__10401),
            .lcout(\POWERLED.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__12079),
            .in2(N__11814),
            .in3(N__10392),
            .lcout(\POWERLED.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(N__11793),
            .in2(N__12113),
            .in3(N__10380),
            .lcout(\POWERLED.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_6_4  (
            .in0(_gnd_net_),
            .in1(N__12109),
            .in2(N__12213),
            .in3(N__10524),
            .lcout(\POWERLED.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_6_5  (
            .in0(N__10504),
            .in1(N__12168),
            .in2(N__12084),
            .in3(N__10515),
            .lcout(\POWERLED.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_6_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_6_6  (
            .in0(_gnd_net_),
            .in1(N__12135),
            .in2(_gnd_net_),
            .in3(N__10512),
            .lcout(\POWERLED.mult1_un110_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_6_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11835),
            .lcout(\POWERLED.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13019),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(\POWERLED.mult1_un96_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_7_1  (
            .in0(_gnd_net_),
            .in1(N__12972),
            .in2(N__12269),
            .in3(N__10476),
            .lcout(\POWERLED.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(N__12265),
            .in2(N__12066),
            .in3(N__10473),
            .lcout(\POWERLED.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(N__12054),
            .in2(N__12299),
            .in3(N__10470),
            .lcout(\POWERLED.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_7_4  (
            .in0(_gnd_net_),
            .in1(N__12295),
            .in2(N__12336),
            .in3(N__10467),
            .lcout(\POWERLED.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_7_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_7_5  (
            .in0(N__12195),
            .in1(N__12324),
            .in2(N__12270),
            .in3(N__10608),
            .lcout(\POWERLED.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_7_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_7_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_7_6  (
            .in0(_gnd_net_),
            .in1(N__12315),
            .in2(_gnd_net_),
            .in3(N__10605),
            .lcout(\POWERLED.mult1_un96_sum_s_8 ),
            .ltout(\POWERLED.mult1_un96_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_5_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_5_7_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_5_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10602),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10998),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(\POWERLED.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__10599),
            .in2(N__10550),
            .in3(N__10593),
            .lcout(\POWERLED.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_8_2  (
            .in0(_gnd_net_),
            .in1(N__10546),
            .in2(N__10590),
            .in3(N__10581),
            .lcout(\POWERLED.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_8_3  (
            .in0(_gnd_net_),
            .in1(N__10578),
            .in2(N__10734),
            .in3(N__10572),
            .lcout(\POWERLED.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_8_4  (
            .in0(_gnd_net_),
            .in1(N__10732),
            .in2(N__10569),
            .in3(N__10560),
            .lcout(\POWERLED.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_8_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_8_5  (
            .in0(N__10665),
            .in1(N__10557),
            .in2(N__10551),
            .in3(N__10533),
            .lcout(\POWERLED.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_8_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_8_6  (
            .in0(N__10748),
            .in1(N__10733),
            .in2(N__10719),
            .in3(N__10710),
            .lcout(\POWERLED.mult1_un61_sum_s_8 ),
            .ltout(\POWERLED.mult1_un61_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_5_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_5_8_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_5_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10707),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12726),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\POWERLED.mult1_un68_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(N__10704),
            .in2(N__10628),
            .in3(N__10695),
            .lcout(\POWERLED.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__10624),
            .in2(N__10692),
            .in3(N__10683),
            .lcout(\POWERLED.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(N__10680),
            .in2(N__10671),
            .in3(N__10674),
            .lcout(\POWERLED.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(N__10669),
            .in2(N__10647),
            .in3(N__10638),
            .lcout(\POWERLED.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_9_5  (
            .in0(N__12654),
            .in1(N__10635),
            .in2(N__10629),
            .in3(N__10611),
            .lcout(\POWERLED.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_9_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10932),
            .in3(N__10923),
            .lcout(\POWERLED.mult1_un68_sum_s_8 ),
            .ltout(\POWERLED.mult1_un68_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_9_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10920),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIVL3D_0_LC_5_10_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNIVL3D_0_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIVL3D_0_LC_5_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \POWERLED.dutycycle_RNIVL3D_0_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__14535),
            .in2(N__14163),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_dutycycle_1_axb_0 ),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\POWERLED.un1_dutycycle_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_5_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_5_10_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14577),
            .in3(N__10872),
            .lcout(\POWERLED.mult1_un138_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_0 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_5_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_5_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__13767),
            .in2(N__13713),
            .in3(N__10839),
            .lcout(\POWERLED.mult1_un131_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_1 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_5_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_5_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__13140),
            .in2(N__13157),
            .in3(N__10806),
            .lcout(\POWERLED.mult1_un124_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_2 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_5_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_5_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__12498),
            .in2(N__13131),
            .in3(N__10773),
            .lcout(\POWERLED.mult1_un117_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_3 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_5_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_5_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(N__12687),
            .in2(N__12507),
            .in3(N__10755),
            .lcout(\POWERLED.mult1_un110_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_4 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_5_10_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_5_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(N__13167),
            .in2(N__13182),
            .in3(N__10752),
            .lcout(\POWERLED.mult1_un103_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_5 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_5_10_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_5_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(N__12693),
            .in2(N__13326),
            .in3(N__11013),
            .lcout(\POWERLED.mult1_un96_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_6 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_5_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_5_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__12797),
            .in2(N__12519),
            .in3(N__11010),
            .lcout(\POWERLED.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\POWERLED.un1_dutycycle_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_5_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_5_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__12672),
            .in2(N__12765),
            .in3(N__11007),
            .lcout(\POWERLED.mult1_un82_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_8 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_5_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_5_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__12750),
            .in2(N__13851),
            .in3(N__11004),
            .lcout(\POWERLED.mult1_un75_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_5_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_5_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__12774),
            .in2(N__12876),
            .in3(N__11001),
            .lcout(\POWERLED.mult1_un68_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_5_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_5_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__12744),
            .in2(N__12735),
            .in3(N__10980),
            .lcout(\POWERLED.mult1_un61_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_5_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_5_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(N__12756),
            .in2(N__12843),
            .in3(N__10959),
            .lcout(\POWERLED.mult1_un54_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_5_11_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_5_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__12852),
            .in2(N__12783),
            .in3(N__10938),
            .lcout(\POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_5_11_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_5_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__12699),
            .in2(N__12861),
            .in3(N__10935),
            .lcout(\POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_14 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_5_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_5_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(N__14284),
            .in2(N__12828),
            .in3(N__11127),
            .lcout(\POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71 ),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(\POWERLED.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_5_12_1 .C_ON=1'b0;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_5_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.CO2_THRU_LUT4_0_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11124),
            .lcout(\POWERLED.CO2_THRU_CO ),
            .ltout(\POWERLED.CO2_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_12_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_12_2 .LUT_INIT=16'b1111000011000011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__11111),
            .in2(N__11091),
            .in3(N__11083),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_ns_0_i_0_0_a2_0_0_LC_5_12_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_ns_0_i_0_0_a2_0_0_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_ns_0_i_0_0_a2_0_0_LC_5_12_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \POWERLED.func_state_ns_0_i_0_0_a2_0_0_LC_5_12_4  (
            .in0(N__14682),
            .in1(N__16460),
            .in2(_gnd_net_),
            .in3(N__16535),
            .lcout(\POWERLED.N_222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.N_55_i_i_o6_LC_5_12_5 .C_ON=1'b0;
    defparam \POWERLED.N_55_i_i_o6_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.N_55_i_i_o6_LC_5_12_5 .LUT_INIT=16'b0111011101110111;
    LogicCell40 \POWERLED.N_55_i_i_o6_LC_5_12_5  (
            .in0(N__16459),
            .in1(N__14681),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_55),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_0_LC_5_13_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_0_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_0_LC_5_13_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_0_LC_5_13_0  (
            .in0(N__18813),
            .in1(N__11055),
            .in2(N__12818),
            .in3(N__12819),
            .lcout(\VPP_VDDQ.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_0 ),
            .clk(N__19229),
            .ce(),
            .sr(N__12935));
    defparam \VPP_VDDQ.count_1_LC_5_13_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_1_LC_5_13_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_1_LC_5_13_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_1_LC_5_13_1  (
            .in0(N__18799),
            .in1(N__11043),
            .in2(_gnd_net_),
            .in3(N__11031),
            .lcout(\VPP_VDDQ.countZ0Z_1 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_0 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_1 ),
            .clk(N__19229),
            .ce(),
            .sr(N__12935));
    defparam \VPP_VDDQ.count_2_LC_5_13_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_2_LC_5_13_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_LC_5_13_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_2_LC_5_13_2  (
            .in0(N__18814),
            .in1(N__11028),
            .in2(_gnd_net_),
            .in3(N__11016),
            .lcout(\VPP_VDDQ.countZ0Z_2 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_2 ),
            .clk(N__19229),
            .ce(),
            .sr(N__12935));
    defparam \VPP_VDDQ.count_3_LC_5_13_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_3_LC_5_13_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_3_LC_5_13_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_3_LC_5_13_3  (
            .in0(N__18800),
            .in1(N__11271),
            .in2(_gnd_net_),
            .in3(N__11259),
            .lcout(\VPP_VDDQ.countZ0Z_3 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_3 ),
            .clk(N__19229),
            .ce(),
            .sr(N__12935));
    defparam \VPP_VDDQ.count_4_LC_5_13_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_4_LC_5_13_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_4_LC_5_13_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_4_LC_5_13_4  (
            .in0(N__18815),
            .in1(N__11256),
            .in2(_gnd_net_),
            .in3(N__11244),
            .lcout(\VPP_VDDQ.countZ0Z_4 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_4 ),
            .clk(N__19229),
            .ce(),
            .sr(N__12935));
    defparam \VPP_VDDQ.count_5_LC_5_13_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_5_LC_5_13_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_5_LC_5_13_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_5_LC_5_13_5  (
            .in0(N__18801),
            .in1(N__11241),
            .in2(_gnd_net_),
            .in3(N__11229),
            .lcout(\VPP_VDDQ.countZ0Z_5 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_5 ),
            .clk(N__19229),
            .ce(),
            .sr(N__12935));
    defparam \VPP_VDDQ.count_6_LC_5_13_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_6_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_6_LC_5_13_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_6_LC_5_13_6  (
            .in0(N__18816),
            .in1(N__11226),
            .in2(_gnd_net_),
            .in3(N__11214),
            .lcout(\VPP_VDDQ.countZ0Z_6 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_6 ),
            .clk(N__19229),
            .ce(),
            .sr(N__12935));
    defparam \VPP_VDDQ.count_7_LC_5_13_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_7_LC_5_13_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_7_LC_5_13_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_7_LC_5_13_7  (
            .in0(N__18802),
            .in1(N__11210),
            .in2(_gnd_net_),
            .in3(N__11196),
            .lcout(\VPP_VDDQ.countZ0Z_7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_7 ),
            .clk(N__19229),
            .ce(),
            .sr(N__12935));
    defparam \VPP_VDDQ.count_8_LC_5_14_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_8_LC_5_14_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_8_LC_5_14_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_8_LC_5_14_0  (
            .in0(N__18820),
            .in1(N__11193),
            .in2(_gnd_net_),
            .in3(N__11181),
            .lcout(\VPP_VDDQ.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_8 ),
            .clk(N__19225),
            .ce(),
            .sr(N__12934));
    defparam \VPP_VDDQ.count_9_LC_5_14_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_9_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_9_LC_5_14_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_9_LC_5_14_1  (
            .in0(N__18805),
            .in1(N__11178),
            .in2(_gnd_net_),
            .in3(N__11166),
            .lcout(\VPP_VDDQ.countZ0Z_9 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_8 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_9 ),
            .clk(N__19225),
            .ce(),
            .sr(N__12934));
    defparam \VPP_VDDQ.count_10_LC_5_14_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_10_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_10_LC_5_14_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_10_LC_5_14_2  (
            .in0(N__18817),
            .in1(N__11162),
            .in2(_gnd_net_),
            .in3(N__11148),
            .lcout(\VPP_VDDQ.countZ0Z_10 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_10 ),
            .clk(N__19225),
            .ce(),
            .sr(N__12934));
    defparam \VPP_VDDQ.count_11_LC_5_14_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_11_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_11_LC_5_14_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_11_LC_5_14_3  (
            .in0(N__18803),
            .in1(N__11144),
            .in2(_gnd_net_),
            .in3(N__11130),
            .lcout(\VPP_VDDQ.countZ0Z_11 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_11 ),
            .clk(N__19225),
            .ce(),
            .sr(N__12934));
    defparam \VPP_VDDQ.count_12_LC_5_14_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_12_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_12_LC_5_14_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_12_LC_5_14_4  (
            .in0(N__18818),
            .in1(N__11475),
            .in2(_gnd_net_),
            .in3(N__11463),
            .lcout(\VPP_VDDQ.countZ0Z_12 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_12 ),
            .clk(N__19225),
            .ce(),
            .sr(N__12934));
    defparam \VPP_VDDQ.count_13_LC_5_14_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_13_LC_5_14_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_13_LC_5_14_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_13_LC_5_14_5  (
            .in0(N__18804),
            .in1(N__11460),
            .in2(_gnd_net_),
            .in3(N__11448),
            .lcout(\VPP_VDDQ.countZ0Z_13 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_13 ),
            .clk(N__19225),
            .ce(),
            .sr(N__12934));
    defparam \VPP_VDDQ.count_14_LC_5_14_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_14_LC_5_14_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_14_LC_5_14_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_14_LC_5_14_6  (
            .in0(N__18819),
            .in1(N__11445),
            .in2(_gnd_net_),
            .in3(N__11433),
            .lcout(\VPP_VDDQ.countZ0Z_14 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14 ),
            .clk(N__19225),
            .ce(),
            .sr(N__12934));
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_14_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(N__17297),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_14 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_15_LC_5_15_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_15_LC_5_15_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_esr_15_LC_5_15_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \VPP_VDDQ.count_esr_15_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__11426),
            .in2(_gnd_net_),
            .in3(N__11430),
            .lcout(\VPP_VDDQ.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19230),
            .ce(N__12912),
            .sr(N__12936));
    defparam \POWERLED.un1_count_1_cry_1_c_LC_6_3_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_1_cry_1_c_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_1_cry_1_c_LC_6_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_1_cry_1_c_LC_6_3_0  (
            .in0(_gnd_net_),
            .in1(N__11404),
            .in2(N__11385),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(\POWERLED.un1_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_2_LC_6_3_1 .C_ON=1'b1;
    defparam \POWERLED.count_2_LC_6_3_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_2_LC_6_3_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_2_LC_6_3_1  (
            .in0(N__18760),
            .in1(N__11341),
            .in2(_gnd_net_),
            .in3(N__11313),
            .lcout(\POWERLED.countZ0Z_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_1 ),
            .carryout(\POWERLED.un1_count_1_cry_2 ),
            .clk(N__18958),
            .ce(),
            .sr(N__11885));
    defparam \POWERLED.count_3_LC_6_3_2 .C_ON=1'b1;
    defparam \POWERLED.count_3_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_3_LC_6_3_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_3_LC_6_3_2  (
            .in0(N__18757),
            .in1(N__11302),
            .in2(_gnd_net_),
            .in3(N__11274),
            .lcout(\POWERLED.countZ0Z_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_2 ),
            .carryout(\POWERLED.un1_count_1_cry_3 ),
            .clk(N__18958),
            .ce(),
            .sr(N__11885));
    defparam \POWERLED.count_4_LC_6_3_3 .C_ON=1'b1;
    defparam \POWERLED.count_4_LC_6_3_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_4_LC_6_3_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_4_LC_6_3_3  (
            .in0(N__18761),
            .in1(N__11776),
            .in2(_gnd_net_),
            .in3(N__11748),
            .lcout(\POWERLED.countZ0Z_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_3 ),
            .carryout(\POWERLED.un1_count_1_cry_4 ),
            .clk(N__18958),
            .ce(),
            .sr(N__11885));
    defparam \POWERLED.count_5_LC_6_3_4 .C_ON=1'b1;
    defparam \POWERLED.count_5_LC_6_3_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_5_LC_6_3_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_5_LC_6_3_4  (
            .in0(N__18758),
            .in1(N__11737),
            .in2(_gnd_net_),
            .in3(N__11709),
            .lcout(\POWERLED.countZ0Z_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_4 ),
            .carryout(\POWERLED.un1_count_1_cry_5 ),
            .clk(N__18958),
            .ce(),
            .sr(N__11885));
    defparam \POWERLED.count_6_LC_6_3_5 .C_ON=1'b1;
    defparam \POWERLED.count_6_LC_6_3_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_6_LC_6_3_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_6_LC_6_3_5  (
            .in0(N__18762),
            .in1(N__11695),
            .in2(_gnd_net_),
            .in3(N__11667),
            .lcout(\POWERLED.countZ0Z_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_5 ),
            .carryout(\POWERLED.un1_count_1_cry_6 ),
            .clk(N__18958),
            .ce(),
            .sr(N__11885));
    defparam \POWERLED.count_7_LC_6_3_6 .C_ON=1'b1;
    defparam \POWERLED.count_7_LC_6_3_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_7_LC_6_3_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_7_LC_6_3_6  (
            .in0(N__18759),
            .in1(N__11656),
            .in2(_gnd_net_),
            .in3(N__11628),
            .lcout(\POWERLED.countZ0Z_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_6 ),
            .carryout(\POWERLED.un1_count_1_cry_7 ),
            .clk(N__18958),
            .ce(),
            .sr(N__11885));
    defparam \POWERLED.count_8_LC_6_3_7 .C_ON=1'b1;
    defparam \POWERLED.count_8_LC_6_3_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_8_LC_6_3_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_8_LC_6_3_7  (
            .in0(N__18763),
            .in1(N__11617),
            .in2(_gnd_net_),
            .in3(N__11589),
            .lcout(\POWERLED.countZ0Z_8 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_7 ),
            .carryout(\POWERLED.un1_count_1_cry_8 ),
            .clk(N__18958),
            .ce(),
            .sr(N__11885));
    defparam \POWERLED.count_9_LC_6_4_0 .C_ON=1'b1;
    defparam \POWERLED.count_9_LC_6_4_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_9_LC_6_4_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_9_LC_6_4_0  (
            .in0(N__18774),
            .in1(N__11581),
            .in2(_gnd_net_),
            .in3(N__11553),
            .lcout(\POWERLED.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(\POWERLED.un1_count_1_cry_9 ),
            .clk(N__19022),
            .ce(),
            .sr(N__11878));
    defparam \POWERLED.count_10_LC_6_4_1 .C_ON=1'b1;
    defparam \POWERLED.count_10_LC_6_4_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_10_LC_6_4_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_10_LC_6_4_1  (
            .in0(N__18775),
            .in1(N__11541),
            .in2(_gnd_net_),
            .in3(N__11511),
            .lcout(\POWERLED.countZ0Z_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_9 ),
            .carryout(\POWERLED.un1_count_1_cry_10 ),
            .clk(N__19022),
            .ce(),
            .sr(N__11878));
    defparam \POWERLED.count_11_LC_6_4_2 .C_ON=1'b1;
    defparam \POWERLED.count_11_LC_6_4_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_11_LC_6_4_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_11_LC_6_4_2  (
            .in0(N__18772),
            .in1(N__11503),
            .in2(_gnd_net_),
            .in3(N__11478),
            .lcout(\POWERLED.countZ0Z_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_10 ),
            .carryout(\POWERLED.un1_count_1_cry_11 ),
            .clk(N__19022),
            .ce(),
            .sr(N__11878));
    defparam \POWERLED.count_12_LC_6_4_3 .C_ON=1'b1;
    defparam \POWERLED.count_12_LC_6_4_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_12_LC_6_4_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_12_LC_6_4_3  (
            .in0(N__18776),
            .in1(N__12040),
            .in2(_gnd_net_),
            .in3(N__12015),
            .lcout(\POWERLED.countZ0Z_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_11 ),
            .carryout(\POWERLED.un1_count_1_cry_12 ),
            .clk(N__19022),
            .ce(),
            .sr(N__11878));
    defparam \POWERLED.count_13_LC_6_4_4 .C_ON=1'b1;
    defparam \POWERLED.count_13_LC_6_4_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_13_LC_6_4_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_13_LC_6_4_4  (
            .in0(N__18773),
            .in1(N__12007),
            .in2(_gnd_net_),
            .in3(N__11979),
            .lcout(\POWERLED.countZ0Z_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_12 ),
            .carryout(\POWERLED.un1_count_1_cry_13 ),
            .clk(N__19022),
            .ce(),
            .sr(N__11878));
    defparam \POWERLED.count_14_LC_6_4_5 .C_ON=1'b1;
    defparam \POWERLED.count_14_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_14_LC_6_4_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_14_LC_6_4_5  (
            .in0(N__18777),
            .in1(N__11968),
            .in2(_gnd_net_),
            .in3(N__11940),
            .lcout(\POWERLED.countZ0Z_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_13 ),
            .carryout(\POWERLED.un1_count_1_cry_14 ),
            .clk(N__19022),
            .ce(),
            .sr(N__11878));
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_6  (
            .in0(_gnd_net_),
            .in1(N__17293),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_14 ),
            .carryout(\POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_6_4_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_6_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_6_4_7  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__17301),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryout(\POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_esr_15_LC_6_5_0 .C_ON=1'b0;
    defparam \POWERLED.count_esr_15_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_esr_15_LC_6_5_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.count_esr_15_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(N__11925),
            .in2(_gnd_net_),
            .in3(N__11937),
            .lcout(\POWERLED.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19023),
            .ce(N__11895),
            .sr(N__11886));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_6_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_6_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__11834),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(\POWERLED.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_6_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_6_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__12999),
            .in2(N__12152),
            .in3(N__11805),
            .lcout(\POWERLED.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_6_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_6_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__12148),
            .in2(N__11802),
            .in3(N__11787),
            .lcout(\POWERLED.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_6_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_6_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__12219),
            .in2(N__12201),
            .in3(N__12204),
            .lcout(\POWERLED.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_6_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_6_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(N__12199),
            .in2(N__12177),
            .in3(N__12162),
            .lcout(\POWERLED.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_6_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_6_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_6_6_5  (
            .in0(N__12105),
            .in1(N__12159),
            .in2(N__12153),
            .in3(N__12129),
            .lcout(\POWERLED.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_6_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_6_6_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12126),
            .in3(N__12117),
            .lcout(\POWERLED.mult1_un103_sum_s_8 ),
            .ltout(\POWERLED.mult1_un103_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_6_6_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_6_6_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_6_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12087),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_6_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_6_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(N__12989),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(\POWERLED.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_6_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_6_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_6_7_1  (
            .in0(_gnd_net_),
            .in1(N__13188),
            .in2(N__12422),
            .in3(N__12057),
            .lcout(\POWERLED.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_6_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_6_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(N__12418),
            .in2(N__12240),
            .in3(N__12048),
            .lcout(\POWERLED.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_6_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_6_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_6_7_3  (
            .in0(_gnd_net_),
            .in1(N__12228),
            .in2(N__12452),
            .in3(N__12327),
            .lcout(\POWERLED.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_6_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_6_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(N__12448),
            .in2(N__12492),
            .in3(N__12318),
            .lcout(\POWERLED.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_6_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_6_7_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_6_7_5  (
            .in0(N__12291),
            .in1(N__12480),
            .in2(N__12423),
            .in3(N__12309),
            .lcout(\POWERLED.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_6_7_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_6_7_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_6_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12471),
            .in3(N__12306),
            .lcout(\POWERLED.mult1_un89_sum_s_8 ),
            .ltout(\POWERLED.mult1_un89_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_6_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_6_7_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_6_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12273),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13211),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_8_0_),
            .carryout(\POWERLED.mult1_un82_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_8_1  (
            .in0(_gnd_net_),
            .in1(N__12252),
            .in2(N__12536),
            .in3(N__12231),
            .lcout(\POWERLED.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_8_2  (
            .in0(_gnd_net_),
            .in1(N__12532),
            .in2(N__12384),
            .in3(N__12222),
            .lcout(\POWERLED.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_8_3  (
            .in0(_gnd_net_),
            .in1(N__12363),
            .in2(N__12566),
            .in3(N__12483),
            .lcout(\POWERLED.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_8_4  (
            .in0(_gnd_net_),
            .in1(N__12562),
            .in2(N__12348),
            .in3(N__12474),
            .lcout(\POWERLED.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_8_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_8_5  (
            .in0(N__12444),
            .in1(N__12627),
            .in2(N__12537),
            .in3(N__12462),
            .lcout(\POWERLED.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_8_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12594),
            .in3(N__12459),
            .lcout(\POWERLED.mult1_un82_sum_s_8 ),
            .ltout(\POWERLED.mult1_un82_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_6_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_6_8_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_6_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12426),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_9_0  (
            .in0(_gnd_net_),
            .in1(N__12401),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(\POWERLED.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__12708),
            .in2(N__12611),
            .in3(N__12375),
            .lcout(\POWERLED.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_9_2  (
            .in0(_gnd_net_),
            .in1(N__12607),
            .in2(N__12372),
            .in3(N__12357),
            .lcout(\POWERLED.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(N__12354),
            .in2(N__12662),
            .in3(N__12339),
            .lcout(\POWERLED.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_9_4  (
            .in0(_gnd_net_),
            .in1(N__12658),
            .in2(N__12636),
            .in3(N__12621),
            .lcout(\POWERLED.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_9_5  (
            .in0(N__12558),
            .in1(N__12618),
            .in2(N__12612),
            .in3(N__12585),
            .lcout(\POWERLED.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_9_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12582),
            .in3(N__12573),
            .lcout(\POWERLED.mult1_un75_sum_s_8 ),
            .ltout(\POWERLED.mult1_un75_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_9_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12540),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJL1R1_6_LC_6_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJL1R1_6_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJL1R1_6_LC_6_10_0 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNIJL1R1_6_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12798),
            .in3(N__12678),
            .lcout(\POWERLED.dutycycle_RNIJL1R1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNIMOAE_5_LC_6_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNIMOAE_5_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNIMOAE_5_LC_6_10_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_fast_RNIMOAE_5_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14348),
            .in3(N__14897),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_1_19_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIEJ021_4_LC_6_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIEJ021_4_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIEJ021_4_LC_6_10_2 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \POWERLED.dutycycle_RNIEJ021_4_LC_6_10_2  (
            .in0(N__14321),
            .in1(N__14162),
            .in2(N__12510),
            .in3(N__14223),
            .lcout(\POWERLED.dutycycle_RNIEJ021Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQAI81_4_LC_6_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQAI81_4_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQAI81_4_LC_6_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNIQAI81_4_LC_6_10_3  (
            .in0(N__13127),
            .in1(N__14149),
            .in2(N__14226),
            .in3(N__14320),
            .lcout(\POWERLED.dutycycle_RNIQAI81Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_10_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12722),
            .lcout(\POWERLED.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI53MG_14_LC_6_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI53MG_14_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI53MG_14_LC_6_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI53MG_14_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(N__14036),
            .in2(_gnd_net_),
            .in3(N__13977),
            .lcout(\POWERLED.dutycycle_RNI53MGZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNIVCSK_5_LC_6_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNIVCSK_5_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNIVCSK_5_LC_6_10_6 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_fast_RNIVCSK_5_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(N__14344),
            .in2(N__14647),
            .in3(N__14077),
            .lcout(\POWERLED.dutycycle_fast_RNIVCSKZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNI8MSK_5_LC_6_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNI8MSK_5_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNI8MSK_5_LC_6_10_7 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_fast_RNI8MSK_5_LC_6_10_7  (
            .in0(_gnd_net_),
            .in1(N__14898),
            .in2(N__14349),
            .in3(N__14322),
            .lcout(\POWERLED.dutycycle_fast_RNI8MSKZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJNBA1_6_LC_6_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJNBA1_6_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJNBA1_6_LC_6_11_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNIJNBA1_6_LC_6_11_0  (
            .in0(N__13252),
            .in1(N__13322),
            .in2(N__14218),
            .in3(N__15029),
            .lcout(\POWERLED.dutycycle_RNIJNBA1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOQLJ_4_LC_6_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOQLJ_4_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOQLJ_4_LC_6_11_1 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_RNIOQLJ_4_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(N__14323),
            .in2(N__14152),
            .in3(N__14199),
            .lcout(\POWERLED.dutycycle_RNIOQLJZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIM0TE_8_LC_6_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIM0TE_8_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIM0TE_8_LC_6_11_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNIM0TE_8_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14990),
            .in3(N__14885),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_1_34_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIUUB41_6_LC_6_11_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIUUB41_6_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIUUB41_6_LC_6_11_3 .LUT_INIT=16'b1110000101111000;
    LogicCell40 \POWERLED.dutycycle_RNIUUB41_6_LC_6_11_3  (
            .in0(N__15028),
            .in1(N__13251),
            .in2(N__12681),
            .in3(N__14198),
            .lcout(\POWERLED.un1_dutycycle_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIB1FL_8_LC_6_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIB1FL_8_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIB1FL_8_LC_6_11_4 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \POWERLED.dutycycle_RNIB1FL_8_LC_6_11_4  (
            .in0(N__14980),
            .in1(_gnd_net_),
            .in2(N__14219),
            .in3(N__14886),
            .lcout(\POWERLED.dutycycle_RNIB1FLZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNILMLM_6_LC_6_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNILMLM_6_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNILMLM_6_LC_6_11_5 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_fast_RNILMLM_6_LC_6_11_5  (
            .in0(_gnd_net_),
            .in1(N__13341),
            .in2(N__15038),
            .in3(N__14197),
            .lcout(\POWERLED.dutycycle_fast_RNILMLMZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI84C11_14_LC_6_11_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI84C11_14_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI84C11_14_LC_6_11_6 .LUT_INIT=16'b0100101101111000;
    LogicCell40 \POWERLED.dutycycle_RNI84C11_14_LC_6_11_6  (
            .in0(N__13965),
            .in1(N__13900),
            .in2(N__14034),
            .in3(N__13966),
            .lcout(\POWERLED.dutycycle_RNI84C11Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQ09G1_10_LC_6_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQ09G1_10_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQ09G1_10_LC_6_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNIQ09G1_10_LC_6_11_7  (
            .in0(N__12875),
            .in1(N__14981),
            .in2(N__15039),
            .in3(N__14017),
            .lcout(\POWERLED.dutycycle_RNIQ09G1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIO2TE_9_LC_6_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIO2TE_9_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIO2TE_9_LC_6_12_0 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNIO2TE_9_LC_6_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13904),
            .in3(N__14930),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_1_39_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI34C41_8_LC_6_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI34C41_8_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI34C41_8_LC_6_12_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI34C41_8_LC_6_12_1  (
            .in0(N__14985),
            .in1(N__14225),
            .in2(N__12768),
            .in3(N__14892),
            .lcout(\POWERLED.dutycycle_RNI34C41Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI73C11_15_LC_6_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI73C11_15_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI73C11_15_LC_6_12_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \POWERLED.dutycycle_RNI73C11_15_LC_6_12_2  (
            .in0(N__13895),
            .in1(N__13970),
            .in2(N__14273),
            .in3(N__14984),
            .lcout(\POWERLED.dutycycle_RNI73C11Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIE4FL_9_LC_6_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIE4FL_9_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIE4FL_9_LC_6_12_3 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_RNIE4FL_9_LC_6_12_3  (
            .in0(_gnd_net_),
            .in1(N__13893),
            .in2(N__14944),
            .in3(N__14893),
            .lcout(\POWERLED.dutycycle_RNIE4FLZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2V0P_10_LC_6_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2V0P_10_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2V0P_10_LC_6_12_4 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_RNI2V0P_10_LC_6_12_4  (
            .in0(_gnd_net_),
            .in1(N__15035),
            .in2(N__14035),
            .in3(N__14982),
            .lcout(\POWERLED.dutycycle_RNI2V0PZ0Z_10 ),
            .ltout(\POWERLED.dutycycle_RNI2V0PZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI712I1_15_LC_6_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI712I1_15_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI712I1_15_LC_6_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNI712I1_15_LC_6_12_5  (
            .in0(N__14983),
            .in1(N__13894),
            .in2(N__12738),
            .in3(N__14256),
            .lcout(\POWERLED.dutycycle_RNI712I1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIO18N_9_LC_6_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIO18N_9_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIO18N_9_LC_6_12_6 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_RNIO18N_9_LC_6_12_6  (
            .in0(_gnd_net_),
            .in1(N__15034),
            .in2(N__13975),
            .in3(N__14934),
            .lcout(\POWERLED.dutycycle_RNIO18NZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIC8C11_15_LC_6_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIC8C11_15_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIC8C11_15_LC_6_12_7 .LUT_INIT=16'b0100101101111000;
    LogicCell40 \POWERLED.dutycycle_RNIC8C11_15_LC_6_12_7  (
            .in0(N__14028),
            .in1(N__13964),
            .in2(N__14274),
            .in3(N__14024),
            .lcout(\POWERLED.dutycycle_RNIC8C11Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI31MG_12_LC_6_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI31MG_12_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI31MG_12_LC_6_13_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI31MG_12_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13905),
            .in3(N__13960),
            .lcout(\POWERLED.dutycycle_RNI31MGZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI31MG_0_12_LC_6_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI31MG_0_12_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI31MG_0_12_LC_6_13_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI31MG_0_12_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13974),
            .in3(N__13896),
            .lcout(\POWERLED.dutycycle_RNI31MG_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI7LE01_0_LC_6_13_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI7LE01_0_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI7LE01_0_LC_6_13_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \POWERLED.func_state_RNI7LE01_0_LC_6_13_2  (
            .in0(N__16706),
            .in1(N__16527),
            .in2(_gnd_net_),
            .in3(N__16084),
            .lcout(),
            .ltout(\POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI446AD_0_LC_6_13_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI446AD_0_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI446AD_0_LC_6_13_3 .LUT_INIT=16'b1111111111010101;
    LogicCell40 \POWERLED.func_state_RNI446AD_0_LC_6_13_3  (
            .in0(N__14709),
            .in1(N__16725),
            .in2(N__12831),
            .in3(N__16007),
            .lcout(\POWERLED.dutycycle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI75MG_15_LC_6_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI75MG_15_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI75MG_15_LC_6_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI75MG_15_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(N__14263),
            .in2(_gnd_net_),
            .in3(N__14029),
            .lcout(\POWERLED.dutycycle_RNI75MGZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNIDNTT1_0_LC_6_14_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNIDNTT1_0_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNIDNTT1_0_LC_6_14_0 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \VPP_VDDQ.curr_state_RNIDNTT1_0_LC_6_14_0  (
            .in0(N__13423),
            .in1(N__13449),
            .in2(_gnd_net_),
            .in3(N__16556),
            .lcout(\VPP_VDDQ.N_108_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_6_14_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_6_14_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_6_14_2  (
            .in0(_gnd_net_),
            .in1(N__13427),
            .in2(_gnd_net_),
            .in3(N__13450),
            .lcout(),
            .ltout(\VPP_VDDQ.N_242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_6_14_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_6_14_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_6_14_3 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_LC_6_14_3  (
            .in0(N__16558),
            .in1(N__12942),
            .in2(N__12801),
            .in3(N__18745),
            .lcout(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19085),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNI8I855_0_LC_6_14_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNI8I855_0_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNI8I855_0_LC_6_14_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.curr_state_RNI8I855_0_LC_6_14_4  (
            .in0(N__13424),
            .in1(N__13448),
            .in2(_gnd_net_),
            .in3(N__13466),
            .lcout(),
            .ltout(N_154_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_111_LC_6_14_5 .C_ON=1'b0;
    defparam \POWERLED.G_111_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_111_LC_6_14_5 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \POWERLED.G_111_LC_6_14_5  (
            .in0(N__13425),
            .in1(N__12951),
            .in2(N__12954),
            .in3(N__18743),
            .lcout(G_111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNINMKE1_1_LC_6_14_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNINMKE1_1_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNINMKE1_1_LC_6_14_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \VPP_VDDQ.curr_state_RNINMKE1_1_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(N__13447),
            .in2(_gnd_net_),
            .in3(N__16557),
            .lcout(N_128),
            .ltout(N_128_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_6_14_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_6_14_7 .LUT_INIT=16'b0101100011001100;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_6_14_7  (
            .in0(N__13426),
            .in1(N__17687),
            .in2(N__12945),
            .in3(N__18744),
            .lcout(\VPP_VDDQ.delayed_vddq_pwrgd_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_6_15_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_6_15_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \VPP_VDDQ.count_esr_RNO_0_15_LC_6_15_7  (
            .in0(_gnd_net_),
            .in1(N__12933),
            .in2(_gnd_net_),
            .in3(N__18764),
            .lcout(\VPP_VDDQ.N_49_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_sys_pwrok_LC_7_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_sys_pwrok_LC_7_1_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_sys_pwrok_LC_7_1_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PCH_PWRGD.un2_sys_pwrok_LC_7_1_0  (
            .in0(_gnd_net_),
            .in1(N__12897),
            .in2(_gnd_net_),
            .in3(N__16968),
            .lcout(\PCH_PWRGD.N_3_i ),
            .ltout(\PCH_PWRGD.N_3_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIC5474_0_LC_7_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIC5474_0_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIC5474_0_LC_7_1_1 .LUT_INIT=16'b1010101111101111;
    LogicCell40 \PCH_PWRGD.curr_state_RNIC5474_0_LC_7_1_1  (
            .in0(N__13073),
            .in1(N__13109),
            .in2(N__12903),
            .in3(N__15385),
            .lcout(),
            .ltout(\PCH_PWRGD.un1_curr_state_0_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI7N705_0_LC_7_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI7N705_0_LC_7_1_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI7N705_0_LC_7_1_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI7N705_0_LC_7_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12900),
            .in3(N__18738),
            .lcout(\PCH_PWRGD.curr_state_RNI7N705Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIHKNI1_0_LC_7_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIHKNI1_0_LC_7_1_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIHKNI1_0_LC_7_1_6 .LUT_INIT=16'b1010111010101010;
    LogicCell40 \PCH_PWRGD.curr_state_RNIHKNI1_0_LC_7_1_6  (
            .in0(N__13110),
            .in1(N__12896),
            .in2(N__13077),
            .in3(N__16969),
            .lcout(\PCH_PWRGD.un1_curr_state10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_0_LC_7_2_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_0_LC_7_2_4 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_0_LC_7_2_4 .LUT_INIT=16'b0100010010100000;
    LogicCell40 \PCH_PWRGD.curr_state_0_LC_7_2_4  (
            .in0(N__13111),
            .in1(N__13091),
            .in2(N__15399),
            .in3(N__13075),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19001),
            .ce(N__18468),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_1_LC_7_2_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_1_LC_7_2_5 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_1_LC_7_2_5 .LUT_INIT=16'b0000010101000100;
    LogicCell40 \PCH_PWRGD.curr_state_1_LC_7_2_5  (
            .in0(N__13074),
            .in1(N__13092),
            .in2(N__15398),
            .in3(N__13112),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19001),
            .ce(N__18468),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.pch_pwrok_LC_7_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.pch_pwrok_LC_7_2_6 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.pch_pwrok_LC_7_2_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \PCH_PWRGD.pch_pwrok_LC_7_2_6  (
            .in0(N__13113),
            .in1(N__13090),
            .in2(_gnd_net_),
            .in3(N__13076),
            .lcout(pch_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19001),
            .ce(N__18468),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_esr_RNO_0_15_LC_7_3_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_esr_RNO_0_15_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_esr_RNO_0_15_LC_7_3_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \PCH_PWRGD.count_esr_RNO_0_15_LC_7_3_6  (
            .in0(_gnd_net_),
            .in1(N__18741),
            .in2(_gnd_net_),
            .in3(N__13575),
            .lcout(\PCH_PWRGD.N_49_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_6_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13023),
            .lcout(\POWERLED.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_7_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12990),
            .lcout(\POWERLED.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIAA8L4_0_LC_7_8_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIAA8L4_0_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIAA8L4_0_LC_7_8_0 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \POWERLED.func_state_RNIAA8L4_0_LC_7_8_0  (
            .in0(N__13790),
            .in1(N__12963),
            .in2(N__16086),
            .in3(N__14833),
            .lcout(\POWERLED.N_200_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI4I7Q_5_LC_7_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI4I7Q_5_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI4I7Q_5_LC_7_8_1 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \POWERLED.dutycycle_RNI4I7Q_5_LC_7_8_1  (
            .in0(N__14644),
            .in1(N__14539),
            .in2(N__13757),
            .in3(N__13262),
            .lcout(\POWERLED.N_117 ),
            .ltout(\POWERLED.N_117_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2GLJ3_5_LC_7_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2GLJ3_5_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2GLJ3_5_LC_7_8_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI2GLJ3_5_LC_7_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12957),
            .in3(N__14834),
            .lcout(\POWERLED.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_8_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13212),
            .lcout(\POWERLED.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI4I7Q_0_5_LC_7_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI4I7Q_0_5_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI4I7Q_0_5_LC_7_8_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \POWERLED.dutycycle_RNI4I7Q_0_5_LC_7_8_6  (
            .in0(N__13261),
            .in1(N__13748),
            .in2(N__14543),
            .in3(N__14645),
            .lcout(\POWERLED.N_234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_5_LC_7_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_5_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_5_LC_7_9_6 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \POWERLED.dutycycle_5_LC_7_9_6  (
            .in0(N__14473),
            .in1(N__15856),
            .in2(N__14374),
            .in3(N__14493),
            .lcout(\POWERLED.dutycycleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18937),
            .ce(N__18433),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6NI81_5_LC_7_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6NI81_5_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6NI81_5_LC_7_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI6NI81_5_LC_7_10_1  (
            .in0(N__13181),
            .in1(N__13250),
            .in2(N__13755),
            .in3(N__14942),
            .lcout(\POWERLED.dutycycle_RNI6NI81Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_6_LC_7_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_6_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_6_LC_7_10_2 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \POWERLED.dutycycle_6_LC_7_10_2  (
            .in0(N__13223),
            .in1(N__15860),
            .in2(N__14477),
            .in3(N__14381),
            .lcout(\POWERLED.dutycycleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19159),
            .ce(N__18476),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIK4I81_6_LC_7_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIK4I81_6_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIK4I81_6_LC_7_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNIK4I81_6_LC_7_10_3  (
            .in0(N__13158),
            .in1(N__13249),
            .in2(N__14087),
            .in3(N__14138),
            .lcout(\POWERLED.dutycycle_RNIK4I81Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_2_LC_7_10_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_2_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_2_LC_7_10_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \POWERLED.dutycycle_2_LC_7_10_4  (
            .in0(N__14466),
            .in1(N__16410),
            .in2(N__13284),
            .in3(N__14717),
            .lcout(\POWERLED.dutycycleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19159),
            .ce(N__18476),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNI2GSK_6_LC_7_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNI2GSK_6_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNI2GSK_6_LC_7_10_5 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_fast_RNI2GSK_6_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(N__13339),
            .in2(N__14088),
            .in3(N__14139),
            .lcout(\POWERLED.dutycycle_fast_RNI2GSKZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_6_LC_7_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_6_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_fast_6_LC_7_10_6 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \POWERLED.dutycycle_fast_6_LC_7_10_6  (
            .in0(N__13224),
            .in1(N__15861),
            .in2(N__14478),
            .in3(N__14382),
            .lcout(\POWERLED.dutycycle_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19159),
            .ce(N__18476),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNIBPSK_6_LC_7_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNIBPSK_6_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNIBPSK_6_LC_7_10_7 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_fast_RNIBPSK_6_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(N__13340),
            .in2(N__13756),
            .in3(N__14943),
            .lcout(\POWERLED.dutycycle_fast_RNIBPSKZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_7_11_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_7_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__13304),
            .in2(N__13308),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\POWERLED.dutycycle_cry_c_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_0_0_LC_7_11_1 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNO_0_0_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_0_0_LC_7_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNO_0_0_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__14534),
            .in2(N__14796),
            .in3(N__13290),
            .lcout(\POWERLED.dutycycle_s_0 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_c_0_THRU_CO ),
            .carryout(\POWERLED.dutycycle_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_0_1_LC_7_11_2 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNO_0_1_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_0_1_LC_7_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNO_0_1_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__14769),
            .in2(N__14646),
            .in3(N__13287),
            .lcout(\POWERLED.dutycycle_s_1 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_0 ),
            .carryout(\POWERLED.dutycycle_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_1_2_LC_7_11_3 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNO_1_2_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_1_2_LC_7_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNO_1_2_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__14770),
            .in2(N__14095),
            .in3(N__13275),
            .lcout(\POWERLED.dutycycle_s_2 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_1 ),
            .carryout(\POWERLED.dutycycle_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_3_LC_7_11_4 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_3_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_3_LC_7_11_4 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_3_LC_7_11_4  (
            .in0(N__14457),
            .in1(N__14151),
            .in2(N__14797),
            .in3(N__13272),
            .lcout(\POWERLED.dutycycleZ0Z_3 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_2 ),
            .carryout(\POWERLED.dutycycle_cry_3 ),
            .clk(N__19214),
            .ce(N__18485),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_4_LC_7_11_5 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_4_LC_7_11_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_4_LC_7_11_5 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_4_LC_7_11_5  (
            .in0(N__14458),
            .in1(N__14774),
            .in2(N__14328),
            .in3(N__13269),
            .lcout(\POWERLED.dutycycleZ0Z_4 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_3 ),
            .carryout(\POWERLED.dutycycle_cry_4 ),
            .clk(N__19214),
            .ce(N__18485),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_cry_c_RNIV95M9_4_LC_7_11_6 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_cry_c_RNIV95M9_4_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_cry_c_RNIV95M9_4_LC_7_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_cry_c_RNIV95M9_4_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__13758),
            .in2(N__14798),
            .in3(N__13266),
            .lcout(\POWERLED.dutycycle_s_5 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_4 ),
            .carryout(\POWERLED.dutycycle_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_cry_c_RNI1C5M9_5_LC_7_11_7 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_cry_c_RNI1C5M9_5_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_cry_c_RNI1C5M9_5_LC_7_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_cry_c_RNI1C5M9_5_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__14778),
            .in2(N__13263),
            .in3(N__13215),
            .lcout(\POWERLED.dutycycle_s_6 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_5 ),
            .carryout(\POWERLED.dutycycle_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_7_LC_7_12_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_7_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_7_LC_7_12_0 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_7_LC_7_12_0  (
            .in0(N__14435),
            .in1(N__14779),
            .in2(N__14224),
            .in3(N__13368),
            .lcout(\POWERLED.dutycycleZ0Z_7 ),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\POWERLED.dutycycle_cry_7 ),
            .clk(N__19210),
            .ce(N__18488),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_8_LC_7_12_1 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_8_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_8_LC_7_12_1 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_8_LC_7_12_1  (
            .in0(N__14432),
            .in1(N__14896),
            .in2(N__14799),
            .in3(N__13365),
            .lcout(\POWERLED.dutycycleZ0Z_8 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_7 ),
            .carryout(\POWERLED.dutycycle_cry_8 ),
            .clk(N__19210),
            .ce(N__18488),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_9_LC_7_12_2 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_9_LC_7_12_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_9_LC_7_12_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_9_LC_7_12_2  (
            .in0(N__14436),
            .in1(N__14783),
            .in2(N__14946),
            .in3(N__13362),
            .lcout(\POWERLED.dutycycleZ0Z_9 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_8 ),
            .carryout(\POWERLED.dutycycle_cry_9 ),
            .clk(N__19210),
            .ce(N__18488),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_10_LC_7_12_3 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_10_LC_7_12_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_10_LC_7_12_3 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_10_LC_7_12_3  (
            .in0(N__14429),
            .in1(N__15037),
            .in2(N__14800),
            .in3(N__13359),
            .lcout(\POWERLED.dutycycleZ0Z_10 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_9 ),
            .carryout(\POWERLED.dutycycle_cry_10 ),
            .clk(N__19210),
            .ce(N__18488),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_11_LC_7_12_4 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_11_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_11_LC_7_12_4 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_11_LC_7_12_4  (
            .in0(N__14433),
            .in1(N__14787),
            .in2(N__14991),
            .in3(N__13356),
            .lcout(\POWERLED.dutycycleZ0Z_11 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_10 ),
            .carryout(\POWERLED.dutycycle_cry_11 ),
            .clk(N__19210),
            .ce(N__18488),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_12_LC_7_12_5 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_12_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_12_LC_7_12_5 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_12_LC_7_12_5  (
            .in0(N__14430),
            .in1(N__13903),
            .in2(N__14801),
            .in3(N__13353),
            .lcout(\POWERLED.dutycycleZ0Z_12 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_11 ),
            .carryout(\POWERLED.dutycycle_cry_12 ),
            .clk(N__19210),
            .ce(N__18488),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_13_LC_7_12_6 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_13_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_13_LC_7_12_6 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_13_LC_7_12_6  (
            .in0(N__14434),
            .in1(N__14791),
            .in2(N__13976),
            .in3(N__13350),
            .lcout(\POWERLED.dutycycleZ0Z_13 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_12 ),
            .carryout(\POWERLED.dutycycle_cry_13 ),
            .clk(N__19210),
            .ce(N__18488),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_14_LC_7_12_7 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_14_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_14_LC_7_12_7 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_14_LC_7_12_7  (
            .in0(N__14431),
            .in1(N__14033),
            .in2(N__14802),
            .in3(N__13347),
            .lcout(\POWERLED.dutycycleZ0Z_14 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_13 ),
            .carryout(\POWERLED.dutycycle_cry_14 ),
            .clk(N__19210),
            .ce(N__18488),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_15_LC_7_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_15_LC_7_13_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_15_LC_7_13_0 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_15_LC_7_13_0  (
            .in0(N__14446),
            .in1(N__14795),
            .in2(N__14285),
            .in3(N__13344),
            .lcout(\POWERLED.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19008),
            .ce(N__18443),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIROMF7_0_LC_7_13_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIROMF7_0_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIROMF7_0_LC_7_13_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \POWERLED.func_state_RNIROMF7_0_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__14710),
            .in2(_gnd_net_),
            .in3(N__16008),
            .lcout(\POWERLED.un1_dutycycle_4_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_1_LC_7_14_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_1_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_1_LC_7_14_3 .LUT_INIT=16'b0000010010101110;
    LogicCell40 \VPP_VDDQ.curr_state_1_LC_7_14_3  (
            .in0(N__13452),
            .in1(N__13428),
            .in2(N__16563),
            .in3(N__13467),
            .lcout(\VPP_VDDQ.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19211),
            .ce(N__18489),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_0_LC_7_14_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_0_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_0_LC_7_14_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \VPP_VDDQ.curr_state_0_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__13451),
            .in2(_gnd_net_),
            .in3(N__16562),
            .lcout(VPP_VDDQ_curr_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19211),
            .ce(N__18489),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_0_LC_8_1_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_0_LC_8_1_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_0_LC_8_1_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_0_LC_8_1_0  (
            .in0(N__18751),
            .in1(N__15273),
            .in2(N__13400),
            .in3(N__13401),
            .lcout(\PCH_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_1_0_),
            .carryout(\PCH_PWRGD.un1_count_1_cry_0 ),
            .clk(N__18894),
            .ce(),
            .sr(N__13576));
    defparam \PCH_PWRGD.count_1_LC_8_1_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_1_LC_8_1_1 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_1_LC_8_1_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_1_LC_8_1_1  (
            .in0(N__18747),
            .in1(N__15441),
            .in2(_gnd_net_),
            .in3(N__13383),
            .lcout(\PCH_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_0 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_1 ),
            .clk(N__18894),
            .ce(),
            .sr(N__13576));
    defparam \PCH_PWRGD.count_2_LC_8_1_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_2_LC_8_1_2 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_2_LC_8_1_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_2_LC_8_1_2  (
            .in0(N__18752),
            .in1(N__15414),
            .in2(_gnd_net_),
            .in3(N__13380),
            .lcout(\PCH_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_1 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_2 ),
            .clk(N__18894),
            .ce(),
            .sr(N__13576));
    defparam \PCH_PWRGD.count_3_LC_8_1_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_3_LC_8_1_3 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_3_LC_8_1_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_3_LC_8_1_3  (
            .in0(N__18748),
            .in1(N__15330),
            .in2(_gnd_net_),
            .in3(N__13377),
            .lcout(\PCH_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_2 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_3 ),
            .clk(N__18894),
            .ce(),
            .sr(N__13576));
    defparam \PCH_PWRGD.count_4_LC_8_1_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_4_LC_8_1_4 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_4_LC_8_1_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_4_LC_8_1_4  (
            .in0(N__18753),
            .in1(N__15357),
            .in2(_gnd_net_),
            .in3(N__13374),
            .lcout(\PCH_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_3 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_4 ),
            .clk(N__18894),
            .ce(),
            .sr(N__13576));
    defparam \PCH_PWRGD.count_5_LC_8_1_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_5_LC_8_1_5 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_5_LC_8_1_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_5_LC_8_1_5  (
            .in0(N__18749),
            .in1(N__15369),
            .in2(_gnd_net_),
            .in3(N__13371),
            .lcout(\PCH_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_4 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_5 ),
            .clk(N__18894),
            .ce(),
            .sr(N__13576));
    defparam \PCH_PWRGD.count_6_LC_8_1_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_6_LC_8_1_6 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_6_LC_8_1_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_6_LC_8_1_6  (
            .in0(N__18754),
            .in1(N__15453),
            .in2(_gnd_net_),
            .in3(N__13494),
            .lcout(\PCH_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_5 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_6 ),
            .clk(N__18894),
            .ce(),
            .sr(N__13576));
    defparam \PCH_PWRGD.count_7_LC_8_1_7 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_7_LC_8_1_7 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_7_LC_8_1_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_7_LC_8_1_7  (
            .in0(N__18750),
            .in1(N__15344),
            .in2(_gnd_net_),
            .in3(N__13491),
            .lcout(\PCH_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_6 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_7 ),
            .clk(N__18894),
            .ce(),
            .sr(N__13576));
    defparam \PCH_PWRGD.count_8_LC_8_2_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_8_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_8_LC_8_2_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_8_LC_8_2_0  (
            .in0(N__18771),
            .in1(N__15300),
            .in2(_gnd_net_),
            .in3(N__13488),
            .lcout(\PCH_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(\PCH_PWRGD.un1_count_1_cry_8 ),
            .clk(N__19013),
            .ce(),
            .sr(N__13581));
    defparam \PCH_PWRGD.count_9_LC_8_2_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_9_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_9_LC_8_2_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_9_LC_8_2_1  (
            .in0(N__18767),
            .in1(N__15312),
            .in2(_gnd_net_),
            .in3(N__13485),
            .lcout(\PCH_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_8 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_9 ),
            .clk(N__19013),
            .ce(),
            .sr(N__13581));
    defparam \PCH_PWRGD.count_10_LC_8_2_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_10_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_10_LC_8_2_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_10_LC_8_2_2  (
            .in0(N__18768),
            .in1(N__15428),
            .in2(_gnd_net_),
            .in3(N__13482),
            .lcout(\PCH_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_9 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_10 ),
            .clk(N__19013),
            .ce(),
            .sr(N__13581));
    defparam \PCH_PWRGD.count_11_LC_8_2_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_11_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_11_LC_8_2_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_11_LC_8_2_3  (
            .in0(N__18765),
            .in1(N__15287),
            .in2(_gnd_net_),
            .in3(N__13479),
            .lcout(\PCH_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_10 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_11 ),
            .clk(N__19013),
            .ce(),
            .sr(N__13581));
    defparam \PCH_PWRGD.count_12_LC_8_2_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_12_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_12_LC_8_2_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_12_LC_8_2_4  (
            .in0(N__18769),
            .in1(N__15230),
            .in2(_gnd_net_),
            .in3(N__13476),
            .lcout(\PCH_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_11 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_12 ),
            .clk(N__19013),
            .ce(),
            .sr(N__13581));
    defparam \PCH_PWRGD.count_13_LC_8_2_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_13_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_13_LC_8_2_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_13_LC_8_2_5  (
            .in0(N__18766),
            .in1(N__15243),
            .in2(_gnd_net_),
            .in3(N__13473),
            .lcout(\PCH_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_12 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_13 ),
            .clk(N__19013),
            .ce(),
            .sr(N__13581));
    defparam \PCH_PWRGD.count_14_LC_8_2_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_14_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_14_LC_8_2_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_14_LC_8_2_6  (
            .in0(N__18770),
            .in1(N__15255),
            .in2(_gnd_net_),
            .in3(N__13470),
            .lcout(\PCH_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_13 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_14 ),
            .clk(N__19013),
            .ce(),
            .sr(N__13581));
    defparam \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_2_7 .C_ON=1'b1;
    defparam \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_2_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_2_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_2_7  (
            .in0(_gnd_net_),
            .in1(N__17292),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_14 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_esr_15_LC_8_3_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_esr_15_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_esr_15_LC_8_3_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \PCH_PWRGD.count_esr_15_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__15216),
            .in2(_gnd_net_),
            .in3(N__13596),
            .lcout(\PCH_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19042),
            .ce(N__13593),
            .sr(N__13580));
    defparam \COUNTER.counter_2_LC_8_4_2 .C_ON=1'b0;
    defparam \COUNTER.counter_2_LC_8_4_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_2_LC_8_4_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_2_LC_8_4_2  (
            .in0(N__13527),
            .in1(N__13541),
            .in2(_gnd_net_),
            .in3(N__15776),
            .lcout(\COUNTER.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19114),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_RNO_LC_8_4_4 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_8_4_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_RNO_LC_8_4_4  (
            .in0(N__13516),
            .in1(N__13540),
            .in2(N__13647),
            .in3(N__15738),
            .lcout(\COUNTER.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_4_LC_8_4_5 .C_ON=1'b0;
    defparam \COUNTER.counter_4_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_4_LC_8_4_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \COUNTER.counter_4_LC_8_4_5  (
            .in0(N__15778),
            .in1(N__13629),
            .in2(_gnd_net_),
            .in3(N__13645),
            .lcout(\COUNTER.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19114),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_3_LC_8_4_7 .C_ON=1'b0;
    defparam \COUNTER.counter_3_LC_8_4_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_3_LC_8_4_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \COUNTER.counter_3_LC_8_4_7  (
            .in0(N__15777),
            .in1(N__13503),
            .in2(_gnd_net_),
            .in3(N__13517),
            .lcout(\COUNTER.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19114),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_c_LC_8_5_0 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_c_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_c_LC_8_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.counter_1_cry_1_c_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__15675),
            .in2(N__15744),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_5_0_),
            .carryout(\COUNTER.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_8_5_1 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_8_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_8_5_1  (
            .in0(_gnd_net_),
            .in1(N__13542),
            .in2(_gnd_net_),
            .in3(N__13521),
            .lcout(\COUNTER.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_1 ),
            .carryout(\COUNTER.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_8_5_2 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_8_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(N__13518),
            .in2(_gnd_net_),
            .in3(N__13497),
            .lcout(\COUNTER.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_2 ),
            .carryout(\COUNTER.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_8_5_3 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_8_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(N__13646),
            .in2(_gnd_net_),
            .in3(N__13623),
            .lcout(\COUNTER.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_3 ),
            .carryout(\COUNTER.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_8_5_4 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_8_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_8_5_4  (
            .in0(_gnd_net_),
            .in1(N__15705),
            .in2(_gnd_net_),
            .in3(N__13620),
            .lcout(\COUNTER.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_4 ),
            .carryout(\COUNTER.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_8_5_5 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_8_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(N__15720),
            .in2(_gnd_net_),
            .in3(N__13617),
            .lcout(\COUNTER.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_5 ),
            .carryout(\COUNTER.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_7_LC_8_5_6 .C_ON=1'b1;
    defparam \COUNTER.counter_7_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_7_LC_8_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_7_LC_8_5_6  (
            .in0(_gnd_net_),
            .in1(N__15689),
            .in2(_gnd_net_),
            .in3(N__13614),
            .lcout(\COUNTER.counterZ0Z_7 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_6 ),
            .carryout(\COUNTER.counter_1_cry_7 ),
            .clk(N__19081),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_8_LC_8_5_7 .C_ON=1'b1;
    defparam \COUNTER.counter_8_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_8_LC_8_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_8_LC_8_5_7  (
            .in0(_gnd_net_),
            .in1(N__15555),
            .in2(_gnd_net_),
            .in3(N__13611),
            .lcout(\COUNTER.counterZ0Z_8 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_7 ),
            .carryout(\COUNTER.counter_1_cry_8 ),
            .clk(N__19081),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_9_LC_8_6_0 .C_ON=1'b1;
    defparam \COUNTER.counter_9_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_9_LC_8_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_9_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__15582),
            .in2(_gnd_net_),
            .in3(N__13608),
            .lcout(\COUNTER.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\COUNTER.counter_1_cry_9 ),
            .clk(N__19115),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_10_LC_8_6_1 .C_ON=1'b1;
    defparam \COUNTER.counter_10_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_10_LC_8_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_10_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__15594),
            .in2(_gnd_net_),
            .in3(N__13605),
            .lcout(\COUNTER.counterZ0Z_10 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_9 ),
            .carryout(\COUNTER.counter_1_cry_10 ),
            .clk(N__19115),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_11_LC_8_6_2 .C_ON=1'b1;
    defparam \COUNTER.counter_11_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_11_LC_8_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_11_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(N__15569),
            .in2(_gnd_net_),
            .in3(N__13602),
            .lcout(\COUNTER.counterZ0Z_11 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_10 ),
            .carryout(\COUNTER.counter_1_cry_11 ),
            .clk(N__19115),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_12_LC_8_6_3 .C_ON=1'b1;
    defparam \COUNTER.counter_12_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_12_LC_8_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_12_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__15495),
            .in2(_gnd_net_),
            .in3(N__13599),
            .lcout(\COUNTER.counterZ0Z_12 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_11 ),
            .carryout(\COUNTER.counter_1_cry_12 ),
            .clk(N__19115),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_13_LC_8_6_4 .C_ON=1'b1;
    defparam \COUNTER.counter_13_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_13_LC_8_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_13_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__15522),
            .in2(_gnd_net_),
            .in3(N__13674),
            .lcout(\COUNTER.counterZ0Z_13 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_12 ),
            .carryout(\COUNTER.counter_1_cry_13 ),
            .clk(N__19115),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_14_LC_8_6_5 .C_ON=1'b1;
    defparam \COUNTER.counter_14_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_14_LC_8_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_14_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(N__15534),
            .in2(_gnd_net_),
            .in3(N__13671),
            .lcout(\COUNTER.counterZ0Z_14 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_13 ),
            .carryout(\COUNTER.counter_1_cry_14 ),
            .clk(N__19115),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_15_LC_8_6_6 .C_ON=1'b1;
    defparam \COUNTER.counter_15_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_15_LC_8_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_15_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(N__15509),
            .in2(_gnd_net_),
            .in3(N__13668),
            .lcout(\COUNTER.counterZ0Z_15 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_14 ),
            .carryout(\COUNTER.counter_1_cry_15 ),
            .clk(N__19115),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_16_LC_8_6_7 .C_ON=1'b1;
    defparam \COUNTER.counter_16_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_16_LC_8_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_16_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(N__15615),
            .in2(_gnd_net_),
            .in3(N__13665),
            .lcout(\COUNTER.counterZ0Z_16 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_15 ),
            .carryout(\COUNTER.counter_1_cry_16 ),
            .clk(N__19115),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_17_LC_8_7_0 .C_ON=1'b1;
    defparam \COUNTER.counter_17_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_17_LC_8_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_17_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__15642),
            .in2(_gnd_net_),
            .in3(N__13662),
            .lcout(\COUNTER.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\COUNTER.counter_1_cry_17 ),
            .clk(N__19093),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_18_LC_8_7_1 .C_ON=1'b1;
    defparam \COUNTER.counter_18_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_18_LC_8_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_18_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__15654),
            .in2(_gnd_net_),
            .in3(N__13659),
            .lcout(\COUNTER.counterZ0Z_18 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_17 ),
            .carryout(\COUNTER.counter_1_cry_18 ),
            .clk(N__19093),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_19_LC_8_7_2 .C_ON=1'b1;
    defparam \COUNTER.counter_19_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_19_LC_8_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_19_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__15629),
            .in2(_gnd_net_),
            .in3(N__13656),
            .lcout(\COUNTER.counterZ0Z_19 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_18 ),
            .carryout(\COUNTER.counter_1_cry_19 ),
            .clk(N__19093),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_20_LC_8_7_3 .C_ON=1'b1;
    defparam \COUNTER.counter_20_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_20_LC_8_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_20_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__15885),
            .in2(_gnd_net_),
            .in3(N__13653),
            .lcout(\COUNTER.counterZ0Z_20 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_19 ),
            .carryout(\COUNTER.counter_1_cry_20 ),
            .clk(N__19093),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_21_LC_8_7_4 .C_ON=1'b1;
    defparam \COUNTER.counter_21_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_21_LC_8_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_21_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__15912),
            .in2(_gnd_net_),
            .in3(N__13650),
            .lcout(\COUNTER.counterZ0Z_21 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_20 ),
            .carryout(\COUNTER.counter_1_cry_21 ),
            .clk(N__19093),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_22_LC_8_7_5 .C_ON=1'b1;
    defparam \COUNTER.counter_22_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_22_LC_8_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_22_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(N__15924),
            .in2(_gnd_net_),
            .in3(N__13701),
            .lcout(\COUNTER.counterZ0Z_22 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_21 ),
            .carryout(\COUNTER.counter_1_cry_22 ),
            .clk(N__19093),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_23_LC_8_7_6 .C_ON=1'b1;
    defparam \COUNTER.counter_23_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_23_LC_8_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_23_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(N__15899),
            .in2(_gnd_net_),
            .in3(N__13698),
            .lcout(\COUNTER.counterZ0Z_23 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_22 ),
            .carryout(\COUNTER.counter_1_cry_23 ),
            .clk(N__19093),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_24_LC_8_7_7 .C_ON=1'b1;
    defparam \COUNTER.counter_24_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_24_LC_8_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_24_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(N__15945),
            .in2(_gnd_net_),
            .in3(N__13695),
            .lcout(\COUNTER.counterZ0Z_24 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_23 ),
            .carryout(\COUNTER.counter_1_cry_24 ),
            .clk(N__19093),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_25_LC_8_8_0 .C_ON=1'b1;
    defparam \COUNTER.counter_25_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_25_LC_8_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_25_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__15972),
            .in2(_gnd_net_),
            .in3(N__13692),
            .lcout(\COUNTER.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\COUNTER.counter_1_cry_25 ),
            .clk(N__19174),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_26_LC_8_8_1 .C_ON=1'b1;
    defparam \COUNTER.counter_26_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_26_LC_8_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_26_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__15984),
            .in2(_gnd_net_),
            .in3(N__13689),
            .lcout(\COUNTER.counterZ0Z_26 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_25 ),
            .carryout(\COUNTER.counter_1_cry_26 ),
            .clk(N__19174),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_27_LC_8_8_2 .C_ON=1'b1;
    defparam \COUNTER.counter_27_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_27_LC_8_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_27_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__15959),
            .in2(_gnd_net_),
            .in3(N__13686),
            .lcout(\COUNTER.counterZ0Z_27 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_26 ),
            .carryout(\COUNTER.counter_1_cry_27 ),
            .clk(N__19174),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_28_LC_8_8_3 .C_ON=1'b1;
    defparam \COUNTER.counter_28_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_28_LC_8_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_28_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__13800),
            .in2(_gnd_net_),
            .in3(N__13683),
            .lcout(\COUNTER.counterZ0Z_28 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_27 ),
            .carryout(\COUNTER.counter_1_cry_28 ),
            .clk(N__19174),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_29_LC_8_8_4 .C_ON=1'b1;
    defparam \COUNTER.counter_29_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_29_LC_8_8_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \COUNTER.counter_29_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13824),
            .in3(N__13680),
            .lcout(\COUNTER.counterZ0Z_29 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_28 ),
            .carryout(\COUNTER.counter_1_cry_29 ),
            .clk(N__19174),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_30_LC_8_8_5 .C_ON=1'b1;
    defparam \COUNTER.counter_30_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_30_LC_8_8_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \COUNTER.counter_30_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13836),
            .in3(N__13677),
            .lcout(\COUNTER.counterZ0Z_30 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_29 ),
            .carryout(\COUNTER.counter_1_cry_30 ),
            .clk(N__19174),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_31_LC_8_8_6 .C_ON=1'b0;
    defparam \COUNTER.counter_31_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_31_LC_8_8_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.counter_31_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__13811),
            .in2(_gnd_net_),
            .in3(N__13839),
            .lcout(\COUNTER.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19174),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_RNO_LC_8_8_7 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_8_8_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_7_c_RNO_LC_8_8_7  (
            .in0(N__13832),
            .in1(N__13820),
            .in2(N__13812),
            .in3(N__13799),
            .lcout(\COUNTER.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5J285_5_LC_8_9_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5J285_5_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5J285_5_LC_8_9_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.dutycycle_RNI5J285_5_LC_8_9_1  (
            .in0(N__16398),
            .in1(N__16228),
            .in2(N__14838),
            .in3(N__13791),
            .lcout(\POWERLED.N_214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI0AN05_0_0_LC_8_9_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI0AN05_0_0_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI0AN05_0_0_LC_8_9_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \POWERLED.func_state_RNI0AN05_0_0_LC_8_9_2  (
            .in0(N__16229),
            .in1(N__16062),
            .in2(_gnd_net_),
            .in3(N__13776),
            .lcout(\POWERLED.N_248 ),
            .ltout(\POWERLED.N_248_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIV4PD6_1_LC_8_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIV4PD6_1_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIV4PD6_1_LC_8_9_3 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \POWERLED.func_state_RNIV4PD6_1_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__16230),
            .in2(N__13779),
            .in3(N__16285),
            .lcout(\POWERLED.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI0AN05_0_LC_8_9_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI0AN05_0_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI0AN05_0_LC_8_9_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.func_state_RNI0AN05_0_LC_8_9_4  (
            .in0(N__16227),
            .in1(N__16061),
            .in2(_gnd_net_),
            .in3(N__13775),
            .lcout(\POWERLED.N_250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI1UHM1_0_LC_8_9_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI1UHM1_0_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI1UHM1_0_LC_8_9_6 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \POWERLED.func_state_RNI1UHM1_0_LC_8_9_6  (
            .in0(N__16864),
            .in1(N__16356),
            .in2(_gnd_net_),
            .in3(N__16063),
            .lcout(\POWERLED.N_213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIFHLJ_0_LC_8_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIFHLJ_0_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIFHLJ_0_LC_8_10_0 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_RNIFHLJ_0_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__14521),
            .in2(N__14633),
            .in3(N__14318),
            .lcout(\POWERLED.dutycycle_RNIFHLJZ0Z_0 ),
            .ltout(\POWERLED.dutycycle_RNIFHLJZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI16B71_5_LC_8_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI16B71_5_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI16B71_5_LC_8_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNI16B71_5_LC_8_10_1  (
            .in0(N__14070),
            .in1(N__13741),
            .in2(N__13716),
            .in3(N__14615),
            .lcout(\POWERLED.dutycycle_RNI16B71Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_LC_8_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_1_LC_8_10_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \POWERLED.dutycycle_1_LC_8_10_2  (
            .in0(N__14475),
            .in1(N__14565),
            .in2(_gnd_net_),
            .in3(N__14658),
            .lcout(\POWERLED.dutycycleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19181),
            .ce(N__18474),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIFHLJ_0_0_LC_8_10_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIFHLJ_0_0_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIFHLJ_0_0_LC_8_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNIFHLJ_0_0_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__14522),
            .in2(N__14634),
            .in3(N__14319),
            .lcout(\POWERLED.un1_dutycycle_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_0_LC_8_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_0_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_0_LC_8_10_5 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \POWERLED.dutycycle_0_LC_8_10_5  (
            .in0(N__14564),
            .in1(N__14474),
            .in2(N__14556),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19181),
            .ce(N__18474),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_5_LC_8_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_5_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_fast_5_LC_8_10_7 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \POWERLED.dutycycle_fast_5_LC_8_10_7  (
            .in0(N__14492),
            .in1(N__14476),
            .in2(N__14375),
            .in3(N__15862),
            .lcout(\POWERLED.dutycycle_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19181),
            .ce(N__18474),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNID2QT_15_LC_8_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNID2QT_15_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNID2QT_15_LC_8_11_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.dutycycle_RNID2QT_15_LC_8_11_0  (
            .in0(N__14324),
            .in1(N__13953),
            .in2(N__14286),
            .in3(N__14211),
            .lcout(\POWERLED.un2_slp_s3n_2_0_o2_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5QPT_2_LC_8_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5QPT_2_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5QPT_2_LC_8_11_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \POWERLED.dutycycle_RNI5QPT_2_LC_8_11_1  (
            .in0(N__14150),
            .in1(N__14083),
            .in2(N__14037),
            .in3(N__13901),
            .lcout(\POWERLED.un2_slp_s3n_2_0_o2_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI1VLG_10_LC_8_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI1VLG_10_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI1VLG_10_LC_8_11_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI1VLG_10_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__13952),
            .in2(_gnd_net_),
            .in3(N__15033),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_1_44_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIF3561_9_LC_8_11_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIF3561_9_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIF3561_9_LC_8_11_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNIF3561_9_LC_8_11_3  (
            .in0(N__14895),
            .in1(N__13902),
            .in2(N__13854),
            .in3(N__14935),
            .lcout(\POWERLED.dutycycle_RNIF3561Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIC1QT_9_LC_8_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIC1QT_9_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIC1QT_9_LC_8_11_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.dutycycle_RNIC1QT_9_LC_8_11_4  (
            .in0(N__15036),
            .in1(N__14986),
            .in2(N__14945),
            .in3(N__14894),
            .lcout(),
            .ltout(\POWERLED.un2_slp_s3n_2_0_o2_3_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIUTDP2_2_LC_8_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIUTDP2_2_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIUTDP2_2_LC_8_11_5 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \POWERLED.dutycycle_RNIUTDP2_2_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__14853),
            .in2(N__14847),
            .in3(N__14844),
            .lcout(\POWERLED.N_112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNINTA34_1_LC_8_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNINTA34_1_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNINTA34_1_LC_8_11_6 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \POWERLED.func_state_RNINTA34_1_LC_8_11_6  (
            .in0(N__17391),
            .in1(_gnd_net_),
            .in2(N__16299),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI099CL_0_LC_8_11_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI099CL_0_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI099CL_0_LC_8_11_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.func_state_RNI099CL_0_LC_8_11_7  (
            .in0(N__15863),
            .in1(N__15990),
            .in2(N__16189),
            .in3(N__16154),
            .lcout(\POWERLED.count_clk_1_sqmuxa_5_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIPG2D1_2_LC_8_12_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIPG2D1_2_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIPG2D1_2_LC_8_12_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \POWERLED.count_clk_RNIPG2D1_2_LC_8_12_0  (
            .in0(N__15098),
            .in1(N__15059),
            .in2(N__15168),
            .in3(N__15080),
            .lcout(\POWERLED.N_177_5 ),
            .ltout(\POWERLED.N_177_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI2M0Q4_6_LC_8_12_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI2M0Q4_6_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI2M0Q4_6_LC_8_12_1 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \POWERLED.count_clk_RNI2M0Q4_6_LC_8_12_1  (
            .in0(N__15190),
            .in1(N__17653),
            .in2(N__14814),
            .in3(N__16581),
            .lcout(\POWERLED.N_251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI1DHM_6_LC_8_12_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI1DHM_6_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI1DHM_6_LC_8_12_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.count_clk_RNI1DHM_6_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__16702),
            .in2(_gnd_net_),
            .in3(N__15191),
            .lcout(),
            .ltout(\POWERLED.N_368_0_i_i_a6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIBR4E9_6_LC_8_12_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIBR4E9_6_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIBR4E9_6_LC_8_12_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.count_clk_RNIBR4E9_6_LC_8_12_3  (
            .in0(N__14811),
            .in1(N__16582),
            .in2(N__14805),
            .in3(N__15825),
            .lcout(\POWERLED.N_177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_ns_0_i_0_0_a2_1_0_LC_8_12_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_ns_0_i_0_0_a2_1_0_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_ns_0_i_0_0_a2_1_0_LC_8_12_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.func_state_ns_0_i_0_0_a2_1_0_LC_8_12_4  (
            .in0(N__16528),
            .in1(N__16464),
            .in2(_gnd_net_),
            .in3(N__14696),
            .lcout(\POWERLED.N_226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIP4HM_2_LC_8_12_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIP4HM_2_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIP4HM_2_LC_8_12_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \POWERLED.count_clk_RNIP4HM_2_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__15079),
            .in2(_gnd_net_),
            .in3(N__15097),
            .lcout(),
            .ltout(\POWERLED.count_clk_0_sqmuxa_5_0_o2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIP6BO1_4_LC_8_12_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIP6BO1_4_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIP6BO1_4_LC_8_12_6 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \POWERLED.count_clk_RNIP6BO1_4_LC_8_12_6  (
            .in0(N__15164),
            .in1(N__15189),
            .in2(N__15126),
            .in3(N__15058),
            .lcout(\POWERLED.N_141 ),
            .ltout(\POWERLED.N_141_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIS9OC3_4_LC_8_12_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIS9OC3_4_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIS9OC3_4_LC_8_12_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \POWERLED.count_clk_RNIS9OC3_4_LC_8_12_7  (
            .in0(N__16397),
            .in1(_gnd_net_),
            .in2(N__15123),
            .in3(N__16343),
            .lcout(\POWERLED.N_203_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_0_LC_8_13_0 .C_ON=1'b1;
    defparam \POWERLED.count_clk_0_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_0_LC_8_13_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_0_LC_8_13_0  (
            .in0(N__18821),
            .in1(N__17094),
            .in2(N__15120),
            .in3(N__15119),
            .lcout(\POWERLED.count_clkZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\POWERLED.un1_count_clk_1_cry_0 ),
            .clk(N__19223),
            .ce(),
            .sr(N__17021));
    defparam \POWERLED.count_clk_1_LC_8_13_1 .C_ON=1'b1;
    defparam \POWERLED.count_clk_1_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_1_LC_8_13_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_1_LC_8_13_1  (
            .in0(N__18806),
            .in1(N__16607),
            .in2(_gnd_net_),
            .in3(N__15102),
            .lcout(\POWERLED.count_clkZ0Z_1 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_0 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_1 ),
            .clk(N__19223),
            .ce(),
            .sr(N__17021));
    defparam \POWERLED.count_clk_2_LC_8_13_2 .C_ON=1'b1;
    defparam \POWERLED.count_clk_2_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_2_LC_8_13_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_2_LC_8_13_2  (
            .in0(N__18822),
            .in1(N__15099),
            .in2(_gnd_net_),
            .in3(N__15084),
            .lcout(\POWERLED.count_clkZ0Z_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_1 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_2 ),
            .clk(N__19223),
            .ce(),
            .sr(N__17021));
    defparam \POWERLED.count_clk_3_LC_8_13_3 .C_ON=1'b1;
    defparam \POWERLED.count_clk_3_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_3_LC_8_13_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_3_LC_8_13_3  (
            .in0(N__18807),
            .in1(N__15081),
            .in2(_gnd_net_),
            .in3(N__15063),
            .lcout(\POWERLED.count_clkZ0Z_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_2 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_3 ),
            .clk(N__19223),
            .ce(),
            .sr(N__17021));
    defparam \POWERLED.count_clk_4_LC_8_13_4 .C_ON=1'b1;
    defparam \POWERLED.count_clk_4_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_4_LC_8_13_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_4_LC_8_13_4  (
            .in0(N__18823),
            .in1(N__15060),
            .in2(_gnd_net_),
            .in3(N__15045),
            .lcout(\POWERLED.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_3 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_4 ),
            .clk(N__19223),
            .ce(),
            .sr(N__17021));
    defparam \POWERLED.count_clk_5_LC_8_13_5 .C_ON=1'b1;
    defparam \POWERLED.count_clk_5_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_5_LC_8_13_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_5_LC_8_13_5  (
            .in0(N__18808),
            .in1(N__16647),
            .in2(_gnd_net_),
            .in3(N__15042),
            .lcout(\POWERLED.count_clkZ0Z_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_4 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_5 ),
            .clk(N__19223),
            .ce(),
            .sr(N__17021));
    defparam \POWERLED.count_clk_6_LC_8_13_6 .C_ON=1'b1;
    defparam \POWERLED.count_clk_6_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_6_LC_8_13_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_6_LC_8_13_6  (
            .in0(N__18824),
            .in1(N__15192),
            .in2(_gnd_net_),
            .in3(N__15174),
            .lcout(\POWERLED.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_5 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_6 ),
            .clk(N__19223),
            .ce(),
            .sr(N__17021));
    defparam \POWERLED.count_clk_7_LC_8_13_7 .C_ON=1'b1;
    defparam \POWERLED.count_clk_7_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_7_LC_8_13_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_7_LC_8_13_7  (
            .in0(N__18809),
            .in1(N__16703),
            .in2(_gnd_net_),
            .in3(N__15171),
            .lcout(\POWERLED.count_clkZ0Z_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_6 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_7 ),
            .clk(N__19223),
            .ce(),
            .sr(N__17021));
    defparam \POWERLED.count_clk_8_LC_8_14_0 .C_ON=1'b1;
    defparam \POWERLED.count_clk_8_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_8_LC_8_14_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_8_LC_8_14_0  (
            .in0(N__18828),
            .in1(N__15163),
            .in2(_gnd_net_),
            .in3(N__15147),
            .lcout(\POWERLED.count_clkZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\POWERLED.un1_count_clk_1_cry_8 ),
            .clk(N__19222),
            .ce(),
            .sr(N__17014));
    defparam \POWERLED.count_clk_9_LC_8_14_1 .C_ON=1'b1;
    defparam \POWERLED.count_clk_9_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_9_LC_8_14_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_9_LC_8_14_1  (
            .in0(N__18812),
            .in1(N__16628),
            .in2(_gnd_net_),
            .in3(N__15144),
            .lcout(\POWERLED.count_clkZ0Z_9 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_8 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_9 ),
            .clk(N__19222),
            .ce(),
            .sr(N__17014));
    defparam \POWERLED.count_clk_10_LC_8_14_2 .C_ON=1'b1;
    defparam \POWERLED.count_clk_10_LC_8_14_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_10_LC_8_14_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_10_LC_8_14_2  (
            .in0(N__18825),
            .in1(N__17121),
            .in2(_gnd_net_),
            .in3(N__15141),
            .lcout(\POWERLED.count_clkZ0Z_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_9 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_10 ),
            .clk(N__19222),
            .ce(),
            .sr(N__17014));
    defparam \POWERLED.count_clk_11_LC_8_14_3 .C_ON=1'b1;
    defparam \POWERLED.count_clk_11_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_11_LC_8_14_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_11_LC_8_14_3  (
            .in0(N__18810),
            .in1(N__17133),
            .in2(_gnd_net_),
            .in3(N__15138),
            .lcout(\POWERLED.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_10 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_11 ),
            .clk(N__19222),
            .ce(),
            .sr(N__17014));
    defparam \POWERLED.count_clk_12_LC_8_14_4 .C_ON=1'b1;
    defparam \POWERLED.count_clk_12_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_12_LC_8_14_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_12_LC_8_14_4  (
            .in0(N__18826),
            .in1(N__17108),
            .in2(_gnd_net_),
            .in3(N__15135),
            .lcout(\POWERLED.count_clkZ0Z_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_11 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_12 ),
            .clk(N__19222),
            .ce(),
            .sr(N__17014));
    defparam \POWERLED.count_clk_13_LC_8_14_5 .C_ON=1'b1;
    defparam \POWERLED.count_clk_13_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_13_LC_8_14_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_13_LC_8_14_5  (
            .in0(N__18811),
            .in1(N__17052),
            .in2(_gnd_net_),
            .in3(N__15132),
            .lcout(\POWERLED.count_clkZ0Z_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_12 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_13 ),
            .clk(N__19222),
            .ce(),
            .sr(N__17014));
    defparam \POWERLED.count_clk_14_LC_8_14_6 .C_ON=1'b1;
    defparam \POWERLED.count_clk_14_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_14_LC_8_14_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_14_LC_8_14_6  (
            .in0(N__18827),
            .in1(N__17067),
            .in2(_gnd_net_),
            .in3(N__15129),
            .lcout(\POWERLED.count_clkZ0Z_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_13 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_14 ),
            .clk(N__19222),
            .ce(),
            .sr(N__17014));
    defparam \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_8_14_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_8_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_8_14_7  (
            .in0(_gnd_net_),
            .in1(N__17278),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_14 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_esr_15_LC_8_15_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_esr_15_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_esr_15_LC_8_15_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.count_clk_esr_15_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__17081),
            .in2(_gnd_net_),
            .in3(N__15456),
            .lcout(\POWERLED.count_clkZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19242),
            .ce(N__16986),
            .sr(N__17022));
    defparam \PCH_PWRGD.count_RNIESHJ_1_LC_9_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIESHJ_1_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIESHJ_1_LC_9_1_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \PCH_PWRGD.count_RNIESHJ_1_LC_9_1_0  (
            .in0(N__15452),
            .in1(N__15440),
            .in2(N__15429),
            .in3(N__15413),
            .lcout(),
            .ltout(\PCH_PWRGD.un4_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_9_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_9_1_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_9_1_1  (
            .in0(N__15318),
            .in1(N__15261),
            .in2(N__15402),
            .in3(N__15204),
            .lcout(\PCH_PWRGD.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI7J2B_3_LC_9_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI7J2B_3_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI7J2B_3_LC_9_1_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNI7J2B_3_LC_9_1_3  (
            .in0(N__15368),
            .in1(N__15356),
            .in2(N__15345),
            .in3(N__15329),
            .lcout(\PCH_PWRGD.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIN5IJ_0_LC_9_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIN5IJ_0_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIN5IJ_0_LC_9_2_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \PCH_PWRGD.count_RNIN5IJ_0_LC_9_2_0  (
            .in0(N__15311),
            .in1(N__15299),
            .in2(N__15288),
            .in3(N__15272),
            .lcout(\PCH_PWRGD.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_esr_RNIFR521_15_LC_9_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_esr_RNIFR521_15_LC_9_2_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_esr_RNIFR521_15_LC_9_2_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \PCH_PWRGD.count_esr_RNIFR521_15_LC_9_2_7  (
            .in0(N__15254),
            .in1(N__15242),
            .in2(N__15231),
            .in3(N__15215),
            .lcout(\PCH_PWRGD.un4_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_LC_9_4_0 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_0_c_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_LC_9_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(N__15198),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_4_0_),
            .carryout(\COUNTER.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_LC_9_4_1 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_1_c_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_LC_9_4_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_1_c_LC_9_4_1  (
            .in0(_gnd_net_),
            .in1(N__15660),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_0 ),
            .carryout(\COUNTER.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_LC_9_4_2 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_2_c_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_LC_9_4_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_2_c_LC_9_4_2  (
            .in0(_gnd_net_),
            .in1(N__15543),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_1 ),
            .carryout(\COUNTER.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_LC_9_4_3 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_3_c_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_LC_9_4_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_3_c_LC_9_4_3  (
            .in0(_gnd_net_),
            .in1(N__15483),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_2 ),
            .carryout(\COUNTER.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_LC_9_4_4 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_4_c_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_LC_9_4_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_4_c_LC_9_4_4  (
            .in0(_gnd_net_),
            .in1(N__15603),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_3 ),
            .carryout(\COUNTER.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_LC_9_4_5 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_5_c_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_LC_9_4_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_5_c_LC_9_4_5  (
            .in0(_gnd_net_),
            .in1(N__15873),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_4 ),
            .carryout(\COUNTER.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_LC_9_4_6 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_6_c_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_LC_9_4_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_6_c_LC_9_4_6  (
            .in0(_gnd_net_),
            .in1(N__15933),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_5 ),
            .carryout(\COUNTER.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_LC_9_4_7 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_7_c_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_LC_9_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_7_c_LC_9_4_7  (
            .in0(_gnd_net_),
            .in1(N__15474),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_6 ),
            .carryout(\COUNTER.un4_counter_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_THRU_LUT4_0_LC_9_5_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_THRU_LUT4_0_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_THRU_LUT4_0_LC_9_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.un4_counter_7_THRU_LUT4_0_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15462),
            .lcout(\COUNTER.un4_counter_7_THRU_CO ),
            .ltout(\COUNTER.un4_counter_7_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_6_LC_9_5_1 .C_ON=1'b0;
    defparam \COUNTER.counter_6_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_6_LC_9_5_1 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \COUNTER.counter_6_LC_9_5_1  (
            .in0(N__15719),
            .in1(_gnd_net_),
            .in2(N__15459),
            .in3(N__15792),
            .lcout(\COUNTER.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19130),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_LC_9_5_3 .C_ON=1'b0;
    defparam \COUNTER.counter_1_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_1_LC_9_5_3 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_1_LC_9_5_3  (
            .in0(N__15742),
            .in1(N__15674),
            .in2(_gnd_net_),
            .in3(N__15775),
            .lcout(\COUNTER.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19130),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_5_LC_9_5_5 .C_ON=1'b0;
    defparam \COUNTER.counter_5_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_5_LC_9_5_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_5_LC_9_5_5  (
            .in0(N__15786),
            .in1(N__15704),
            .in2(_gnd_net_),
            .in3(N__15773),
            .lcout(\COUNTER.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19130),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_0_LC_9_5_6 .C_ON=1'b0;
    defparam \COUNTER.counter_0_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_0_LC_9_5_6 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \COUNTER.counter_0_LC_9_5_6  (
            .in0(N__15774),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15743),
            .lcout(\COUNTER.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19130),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_RNO_LC_9_5_7 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_9_5_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \COUNTER.un4_counter_1_c_RNO_LC_9_5_7  (
            .in0(N__15718),
            .in1(N__15703),
            .in2(N__15690),
            .in3(N__15673),
            .lcout(\COUNTER.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_RNO_LC_9_6_1 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_9_6_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_4_c_RNO_LC_9_6_1  (
            .in0(N__15653),
            .in1(N__15641),
            .in2(N__15630),
            .in3(N__15614),
            .lcout(\COUNTER.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_RNO_LC_9_6_3 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_9_6_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_2_c_RNO_LC_9_6_3  (
            .in0(N__15593),
            .in1(N__15581),
            .in2(N__15570),
            .in3(N__15554),
            .lcout(\COUNTER.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_RNO_LC_9_6_6 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_9_6_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_3_c_RNO_LC_9_6_6  (
            .in0(N__15533),
            .in1(N__15521),
            .in2(N__15510),
            .in3(N__15494),
            .lcout(\COUNTER.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_RNO_LC_9_7_5 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_9_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_6_c_RNO_LC_9_7_5  (
            .in0(N__15983),
            .in1(N__15971),
            .in2(N__15960),
            .in3(N__15944),
            .lcout(\COUNTER.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_RNO_LC_9_7_6 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_9_7_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_5_c_RNO_LC_9_7_6  (
            .in0(N__15923),
            .in1(N__15911),
            .in2(N__15900),
            .in3(N__15884),
            .lcout(\COUNTER.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_9_8_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_9_8_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_9_8_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_9_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_LC_9_9_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_1_LC_9_9_0 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \POWERLED.func_state_1_LC_9_9_0  (
            .in0(N__16131),
            .in1(N__15798),
            .in2(N__16167),
            .in3(N__16153),
            .lcout(\POWERLED.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19185),
            .ce(N__18473),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_LC_9_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_0_LC_9_9_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.func_state_0_LC_9_9_3  (
            .in0(N__16101),
            .in1(N__15810),
            .in2(N__15864),
            .in3(N__15824),
            .lcout(\POWERLED.func_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19185),
            .ce(N__18473),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_0_0_LC_9_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_0_0_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_0_0_LC_9_10_2 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \POWERLED.func_state_RNO_0_0_LC_9_10_2  (
            .in0(N__16905),
            .in1(N__16123),
            .in2(_gnd_net_),
            .in3(N__16355),
            .lcout(\POWERLED.N_178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_4_1_LC_9_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_4_1_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_4_1_LC_9_10_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.func_state_RNO_4_1_LC_9_10_3  (
            .in0(N__16284),
            .in1(N__16057),
            .in2(_gnd_net_),
            .in3(N__17390),
            .lcout(),
            .ltout(\POWERLED.N_148_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_3_1_LC_9_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_3_1_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_3_1_LC_9_10_4 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \POWERLED.func_state_RNO_3_1_LC_9_10_4  (
            .in0(N__16907),
            .in1(_gnd_net_),
            .in2(N__15804),
            .in3(N__16354),
            .lcout(),
            .ltout(\POWERLED.N_208_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_1_1_LC_9_10_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_1_1_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_1_1_LC_9_10_5 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \POWERLED.func_state_RNO_1_1_LC_9_10_5  (
            .in0(N__16191),
            .in1(N__16906),
            .in2(N__15801),
            .in3(N__16124),
            .lcout(\POWERLED.func_state_ns_i_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_0_1_LC_9_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_0_1_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_0_1_LC_9_10_6 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \POWERLED.func_state_RNO_0_1_LC_9_10_6  (
            .in0(N__16092),
            .in1(N__16190),
            .in2(_gnd_net_),
            .in3(N__16808),
            .lcout(\POWERLED.func_state_ns_i_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI9HME_0_1_LC_9_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI9HME_0_1_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI9HME_0_1_LC_9_10_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.func_state_RNI9HME_0_1_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__16283),
            .in2(_gnd_net_),
            .in3(N__16056),
            .lcout(\POWERLED.N_243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIHPO9A_0_LC_9_11_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIHPO9A_0_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIHPO9A_0_LC_9_11_0 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \POWERLED.func_state_RNIHPO9A_0_LC_9_11_0  (
            .in0(N__16158),
            .in1(N__16122),
            .in2(_gnd_net_),
            .in3(N__16232),
            .lcout(\POWERLED.count_off_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_1_0_LC_9_11_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_1_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_1_0_LC_9_11_1 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \POWERLED.func_state_RNO_1_0_LC_9_11_1  (
            .in0(N__17389),
            .in1(N__16781),
            .in2(N__16085),
            .in3(N__16458),
            .lcout(\POWERLED.N_179 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_2_1_LC_9_11_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_2_1_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_2_1_LC_9_11_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \POWERLED.func_state_RNO_2_1_LC_9_11_2  (
            .in0(N__16287),
            .in1(N__16231),
            .in2(N__16083),
            .in3(N__17388),
            .lcout(\POWERLED.N_211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI9HME_1_LC_9_11_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI9HME_1_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI9HME_1_LC_9_11_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.func_state_RNI9HME_1_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__16286),
            .in2(_gnd_net_),
            .in3(N__16070),
            .lcout(\POWERLED.N_88 ),
            .ltout(\POWERLED.N_88_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIH2SJ1_1_LC_9_11_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIH2SJ1_1_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIH2SJ1_1_LC_9_11_4 .LUT_INIT=16'b1001000110011001;
    LogicCell40 \POWERLED.func_state_RNIH2SJ1_1_LC_9_11_4  (
            .in0(N__16457),
            .in1(N__16526),
            .in2(N__16014),
            .in3(N__16894),
            .lcout(),
            .ltout(\POWERLED.dutycycle_3_sqmuxa_1_i_0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI6KL57_0_LC_9_11_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI6KL57_0_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI6KL57_0_LC_9_11_5 .LUT_INIT=16'b1111010111110100;
    LogicCell40 \POWERLED.func_state_RNI6KL57_0_LC_9_11_5  (
            .in0(N__16525),
            .in1(N__16807),
            .in2(N__16011),
            .in3(N__16322),
            .lcout(\POWERLED.N_366_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI1QOT9_1_LC_9_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI1QOT9_1_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI1QOT9_1_LC_9_11_6 .LUT_INIT=16'b1111101010111010;
    LogicCell40 \POWERLED.func_state_RNI1QOT9_1_LC_9_11_6  (
            .in0(N__16305),
            .in1(N__16396),
            .in2(N__16787),
            .in3(N__17387),
            .lcout(\POWERLED.count_clk_1_sqmuxa_5_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_0_2_LC_9_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_0_2_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_0_2_LC_9_11_7 .LUT_INIT=16'b0111111110101010;
    LogicCell40 \POWERLED.dutycycle_RNO_0_2_LC_9_11_7  (
            .in0(N__16524),
            .in1(N__16288),
            .in2(N__16908),
            .in3(N__16456),
            .lcout(\POWERLED.dutycycle_lm_0_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIORSP5_1_LC_9_12_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIORSP5_1_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIORSP5_1_LC_9_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.func_state_RNIORSP5_1_LC_9_12_0  (
            .in0(N__16344),
            .in1(N__16395),
            .in2(N__16909),
            .in3(N__17372),
            .lcout(\POWERLED.N_205 ),
            .ltout(\POWERLED.N_205_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI5LMRL_1_LC_9_12_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI5LMRL_1_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI5LMRL_1_LC_9_12_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \POWERLED.count_clk_RNI5LMRL_1_LC_9_12_1  (
            .in0(N__16367),
            .in1(N__16920),
            .in2(N__16371),
            .in3(N__16926),
            .lcout(\POWERLED.N_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI4V1H6_1_LC_9_12_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI4V1H6_1_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI4V1H6_1_LC_9_12_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \POWERLED.count_clk_RNI4V1H6_1_LC_9_12_2  (
            .in0(N__16653),
            .in1(N__17373),
            .in2(_gnd_net_),
            .in3(N__17040),
            .lcout(),
            .ltout(\POWERLED.count_clk_0_sqmuxa_5_0_a6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNITU0DB_1_LC_9_12_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNITU0DB_1_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNITU0DB_1_LC_9_12_3 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \POWERLED.count_clk_RNITU0DB_1_LC_9_12_3  (
            .in0(N__16368),
            .in1(N__16895),
            .in2(N__16359),
            .in3(N__16345),
            .lcout(\POWERLED.count_clk_137_tz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIJ13KB_7_LC_9_12_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIJ13KB_7_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIJ13KB_7_LC_9_12_4 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \POWERLED.count_clk_RNIJ13KB_7_LC_9_12_4  (
            .in0(N__16323),
            .in1(N__16701),
            .in2(N__17666),
            .in3(N__16239),
            .lcout(\POWERLED.un2_slp_s3n_2_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIFP6R4_1_LC_9_12_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIFP6R4_1_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIFP6R4_1_LC_9_12_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.func_state_RNIFP6R4_1_LC_9_12_5  (
            .in0(N__17371),
            .in1(N__17649),
            .in2(_gnd_net_),
            .in3(N__16297),
            .lcout(\POWERLED.N_217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIG4MR5_1_LC_9_12_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIG4MR5_1_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIG4MR5_1_LC_9_12_6 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \POWERLED.func_state_RNIG4MR5_1_LC_9_12_6  (
            .in0(N__16298),
            .in1(N__16245),
            .in2(_gnd_net_),
            .in3(N__17370),
            .lcout(\POWERLED.N_149 ),
            .ltout(\POWERLED.N_149_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIS0FM9_7_LC_9_12_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIS0FM9_7_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIS0FM9_7_LC_9_12_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \POWERLED.count_clk_RNIS0FM9_7_LC_9_12_7  (
            .in0(N__16700),
            .in1(N__16233),
            .in2(N__16194),
            .in3(N__16583),
            .lcout(\POWERLED.N_207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNILEIU2_1_LC_9_13_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNILEIU2_1_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNILEIU2_1_LC_9_13_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.count_clk_RNILEIU2_1_LC_9_13_0  (
            .in0(N__17036),
            .in1(N__16605),
            .in2(N__16629),
            .in3(N__16818),
            .lcout(\POWERLED.count_off_1_sqmuxa_i_a6_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI3G101_5_LC_9_13_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI3G101_5_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI3G101_5_LC_9_13_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \POWERLED.count_clk_RNI3G101_5_LC_9_13_1  (
            .in0(N__16645),
            .in1(_gnd_net_),
            .in2(N__16704),
            .in3(N__16910),
            .lcout(\POWERLED.count_off_1_sqmuxa_i_a6_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIA8VP_7_LC_9_13_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIA8VP_7_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIA8VP_7_LC_9_13_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_clk_RNIA8VP_7_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__16693),
            .in2(_gnd_net_),
            .in3(N__16809),
            .lcout(),
            .ltout(\POWERLED.un2_slp_s3n_2_0_a6_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIAIGJ4_7_LC_9_13_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIAIGJ4_7_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIAIGJ4_7_LC_9_13_3 .LUT_INIT=16'b1011101110111010;
    LogicCell40 \POWERLED.count_clk_RNIAIGJ4_7_LC_9_13_3  (
            .in0(N__16788),
            .in1(N__17676),
            .in2(N__16737),
            .in3(N__16584),
            .lcout(),
            .ltout(\POWERLED.un2_slp_s3n_2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI01TCL_7_LC_9_13_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI01TCL_7_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI01TCL_7_LC_9_13_4 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \POWERLED.count_clk_RNI01TCL_7_LC_9_13_4  (
            .in0(N__16707),
            .in1(N__16734),
            .in2(N__16728),
            .in3(N__16721),
            .lcout(\POWERLED.un2_slp_s3n_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIUL2D1_1_LC_9_13_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIUL2D1_1_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIUL2D1_1_LC_9_13_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.count_clk_RNIUL2D1_1_LC_9_13_5  (
            .in0(N__16646),
            .in1(N__16627),
            .in2(N__16705),
            .in3(N__16606),
            .lcout(\POWERLED.count_clk_0_sqmuxa_5_0_a6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIHJP92_1_LC_9_13_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIHJP92_1_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIHJP92_1_LC_9_13_7 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \POWERLED.count_clk_RNIHJP92_1_LC_9_13_7  (
            .in0(N__16644),
            .in1(N__16623),
            .in2(N__16608),
            .in3(N__17035),
            .lcout(\POWERLED.N_146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_LC_9_14_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_LC_9_14_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__18110),
            .in2(_gnd_net_),
            .in3(N__17670),
            .lcout(\VPP_VDDQ.N_238 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIOH1J11_7_LC_9_14_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIOH1J11_7_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIOH1J11_7_LC_9_14_2 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \POWERLED.count_clk_RNIOH1J11_7_LC_9_14_2  (
            .in0(N__17148),
            .in1(N__17139),
            .in2(_gnd_net_),
            .in3(N__18746),
            .lcout(\POWERLED.count_clk_RNIOH1J11Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIUJGM_10_LC_9_14_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIUJGM_10_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIUJGM_10_LC_9_14_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNIUJGM_10_LC_9_14_4  (
            .in0(N__17132),
            .in1(N__17120),
            .in2(N__17109),
            .in3(N__17093),
            .lcout(),
            .ltout(\POWERLED.count_clk_0_sqmuxa_5_0_o2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_esr_RNIKKV71_15_LC_9_14_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_esr_RNIKKV71_15_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_esr_RNIKKV71_15_LC_9_14_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_esr_RNIKKV71_15_LC_9_14_5  (
            .in0(N__17082),
            .in1(N__17066),
            .in2(N__17055),
            .in3(N__17051),
            .lcout(\POWERLED.N_136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_esr_RNO_0_15_LC_9_15_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_esr_RNO_0_15_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_esr_RNO_0_15_LC_9_15_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.count_clk_esr_RNO_0_15_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__18778),
            .in2(_gnd_net_),
            .in3(N__17004),
            .lcout(\POWERLED.N_49_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_11_5_1 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_11_5_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_11_5_1  (
            .in0(N__18027),
            .in1(N__17594),
            .in2(_gnd_net_),
            .in3(N__17561),
            .lcout(vccst_pwrgd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19086),
            .ce(N__18472),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_0_LC_11_5_4 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_0_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.curr_state_0_LC_11_5_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_0_LC_11_5_4  (
            .in0(_gnd_net_),
            .in1(N__17601),
            .in2(_gnd_net_),
            .in3(N__16932),
            .lcout(\ALL_SYS_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19086),
            .ce(N__18472),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_1_LC_11_5_6 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_1_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.curr_state_1_LC_11_5_6 .LUT_INIT=16'b0100010001001110;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_1_LC_11_5_6  (
            .in0(N__17595),
            .in1(N__17184),
            .in2(N__17562),
            .in3(N__18246),
            .lcout(\ALL_SYS_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19086),
            .ce(N__18472),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_RNIHDE82_0_LC_11_6_4 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_RNIHDE82_0_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_RNIHDE82_0_LC_11_6_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_RNIHDE82_0_LC_11_6_4  (
            .in0(N__18019),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17554),
            .lcout(\ALL_SYS_PWRGD.N_247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_RNIK8164_0_LC_11_6_6 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_RNIK8164_0_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_RNIK8164_0_LC_11_6_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_RNIK8164_0_LC_11_6_6  (
            .in0(N__17590),
            .in1(N__17555),
            .in2(_gnd_net_),
            .in3(N__18242),
            .lcout(\ALL_SYS_PWRGD.N_186 ),
            .ltout(\ALL_SYS_PWRGD.N_186_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_RNIDP9H7_1_LC_11_6_7 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_RNIDP9H7_1_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_RNIDP9H7_1_LC_11_6_7 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_RNIDP9H7_1_LC_11_6_7  (
            .in0(N__17592),
            .in1(N__17183),
            .in2(N__17172),
            .in3(N__18737),
            .lcout(\ALL_SYS_PWRGD.curr_state_RNIDP9H7Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_0_LC_11_7_0 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_0_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_0_LC_11_7_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_0_LC_11_7_0  (
            .in0(N__18785),
            .in1(N__17475),
            .in2(N__17529),
            .in3(N__17528),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_0 ),
            .clk(N__19166),
            .ce(),
            .sr(N__17926));
    defparam \ALL_SYS_PWRGD.count_1_LC_11_7_1 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_1_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_1_LC_11_7_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_1_LC_11_7_1  (
            .in0(N__18781),
            .in1(N__17502),
            .in2(_gnd_net_),
            .in3(N__17169),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_0 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_1 ),
            .clk(N__19166),
            .ce(),
            .sr(N__17926));
    defparam \ALL_SYS_PWRGD.count_2_LC_11_7_2 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_2_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_2_LC_11_7_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_2_LC_11_7_2  (
            .in0(N__18786),
            .in1(N__18135),
            .in2(_gnd_net_),
            .in3(N__17166),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_1 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_2 ),
            .clk(N__19166),
            .ce(),
            .sr(N__17926));
    defparam \ALL_SYS_PWRGD.count_3_LC_11_7_3 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_3_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_3_LC_11_7_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_3_LC_11_7_3  (
            .in0(N__18782),
            .in1(N__18174),
            .in2(_gnd_net_),
            .in3(N__17163),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_2 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_3 ),
            .clk(N__19166),
            .ce(),
            .sr(N__17926));
    defparam \ALL_SYS_PWRGD.count_4_LC_11_7_4 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_4_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_4_LC_11_7_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_4_LC_11_7_4  (
            .in0(N__18787),
            .in1(N__18192),
            .in2(_gnd_net_),
            .in3(N__17160),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_3 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_4 ),
            .clk(N__19166),
            .ce(),
            .sr(N__17926));
    defparam \ALL_SYS_PWRGD.count_5_LC_11_7_5 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_5_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_5_LC_11_7_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_5_LC_11_7_5  (
            .in0(N__18783),
            .in1(N__18149),
            .in2(_gnd_net_),
            .in3(N__17157),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_4 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_5 ),
            .clk(N__19166),
            .ce(),
            .sr(N__17926));
    defparam \ALL_SYS_PWRGD.count_6_LC_11_7_6 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_6_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_6_LC_11_7_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_6_LC_11_7_6  (
            .in0(N__18788),
            .in1(N__18219),
            .in2(_gnd_net_),
            .in3(N__17154),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_5 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_6 ),
            .clk(N__19166),
            .ce(),
            .sr(N__17926));
    defparam \ALL_SYS_PWRGD.count_7_LC_11_7_7 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_7_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_7_LC_11_7_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_7_LC_11_7_7  (
            .in0(N__18784),
            .in1(N__18231),
            .in2(_gnd_net_),
            .in3(N__17151),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_6 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_7 ),
            .clk(N__19166),
            .ce(),
            .sr(N__17926));
    defparam \ALL_SYS_PWRGD.count_8_LC_11_8_0 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_8_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_8_LC_11_8_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_8_LC_11_8_0  (
            .in0(N__18795),
            .in1(N__18206),
            .in2(_gnd_net_),
            .in3(N__17322),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_8 ),
            .clk(N__19154),
            .ce(),
            .sr(N__17933));
    defparam \ALL_SYS_PWRGD.count_9_LC_11_8_1 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_9_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_9_LC_11_8_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_9_LC_11_8_1  (
            .in0(N__18791),
            .in1(N__17514),
            .in2(_gnd_net_),
            .in3(N__17319),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_8 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_9 ),
            .clk(N__19154),
            .ce(),
            .sr(N__17933));
    defparam \ALL_SYS_PWRGD.count_10_LC_11_8_2 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_10_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_10_LC_11_8_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_10_LC_11_8_2  (
            .in0(N__18792),
            .in1(N__17489),
            .in2(_gnd_net_),
            .in3(N__17316),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_9 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_10 ),
            .clk(N__19154),
            .ce(),
            .sr(N__17933));
    defparam \ALL_SYS_PWRGD.count_11_LC_11_8_3 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_11_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_11_LC_11_8_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_11_LC_11_8_3  (
            .in0(N__18789),
            .in1(N__18162),
            .in2(_gnd_net_),
            .in3(N__17313),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_10 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_11 ),
            .clk(N__19154),
            .ce(),
            .sr(N__17933));
    defparam \ALL_SYS_PWRGD.count_12_LC_11_8_4 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_12_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_12_LC_11_8_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_12_LC_11_8_4  (
            .in0(N__18793),
            .in1(N__17955),
            .in2(_gnd_net_),
            .in3(N__17310),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_11 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_12 ),
            .clk(N__19154),
            .ce(),
            .sr(N__17933));
    defparam \ALL_SYS_PWRGD.count_13_LC_11_8_5 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_13_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_13_LC_11_8_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_13_LC_11_8_5  (
            .in0(N__18790),
            .in1(N__17982),
            .in2(_gnd_net_),
            .in3(N__17307),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_12 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_13 ),
            .clk(N__19154),
            .ce(),
            .sr(N__17933));
    defparam \ALL_SYS_PWRGD.count_14_LC_11_8_6 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_14_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_14_LC_11_8_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_14_LC_11_8_6  (
            .in0(N__18794),
            .in1(N__17994),
            .in2(_gnd_net_),
            .in3(N__17304),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_13 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_14 ),
            .clk(N__19154),
            .ce(),
            .sr(N__17933));
    defparam \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_8_7 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__17232),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_14 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_esr_15_LC_11_9_0 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_esr_15_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_esr_15_LC_11_9_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALL_SYS_PWRGD.count_esr_15_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__17969),
            .in2(_gnd_net_),
            .in3(N__17187),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19012),
            .ce(N__17895),
            .sr(N__17934));
    defparam \POWERLED.un1_count_off_1_cry_0_c_LC_11_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_off_1_cry_0_c_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_off_1_cry_0_c_LC_11_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_off_1_cry_0_c_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__17879),
            .in2(N__17861),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\POWERLED.un1_count_off_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_1_LC_11_10_1 .C_ON=1'b1;
    defparam \POWERLED.count_off_1_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_1_LC_11_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_1_LC_11_10_1  (
            .in0(N__19361),
            .in1(N__17714),
            .in2(_gnd_net_),
            .in3(N__17346),
            .lcout(\POWERLED.count_offZ0Z_1 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_0 ),
            .carryout(\POWERLED.un1_count_off_1_cry_1 ),
            .clk(N__19155),
            .ce(N__18477),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_off_1_cry_1_THRU_LUT4_0_LC_11_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_off_1_cry_1_THRU_LUT4_0_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_off_1_cry_1_THRU_LUT4_0_LC_11_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.un1_count_off_1_cry_1_THRU_LUT4_0_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__19423),
            .in2(_gnd_net_),
            .in3(N__17343),
            .lcout(\POWERLED.un1_count_off_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_1 ),
            .carryout(\POWERLED.un1_count_off_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_3_LC_11_10_3 .C_ON=1'b1;
    defparam \POWERLED.count_off_3_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_3_LC_11_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_3_LC_11_10_3  (
            .in0(N__19362),
            .in1(N__17408),
            .in2(_gnd_net_),
            .in3(N__17340),
            .lcout(\POWERLED.count_offZ0Z_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_2 ),
            .carryout(\POWERLED.un1_count_off_1_cry_3 ),
            .clk(N__19155),
            .ce(N__18477),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_4_LC_11_10_4 .C_ON=1'b1;
    defparam \POWERLED.count_off_4_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_4_LC_11_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_4_LC_11_10_4  (
            .in0(N__19374),
            .in1(N__17441),
            .in2(_gnd_net_),
            .in3(N__17337),
            .lcout(\POWERLED.count_offZ0Z_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_3 ),
            .carryout(\POWERLED.un1_count_off_1_cry_4 ),
            .clk(N__19155),
            .ce(N__18477),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_off_1_cry_4_THRU_LUT4_0_LC_11_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_off_1_cry_4_THRU_LUT4_0_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_off_1_cry_4_THRU_LUT4_0_LC_11_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.un1_count_off_1_cry_4_THRU_LUT4_0_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__19393),
            .in2(_gnd_net_),
            .in3(N__17334),
            .lcout(\POWERLED.un1_count_off_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_4 ),
            .carryout(\POWERLED.un1_count_off_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_off_1_cry_5_THRU_LUT4_0_LC_11_10_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_off_1_cry_5_THRU_LUT4_0_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_off_1_cry_5_THRU_LUT4_0_LC_11_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.un1_count_off_1_cry_5_THRU_LUT4_0_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__19267),
            .in2(_gnd_net_),
            .in3(N__17331),
            .lcout(\POWERLED.un1_count_off_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_5 ),
            .carryout(\POWERLED.un1_count_off_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_7_LC_11_10_7 .C_ON=1'b1;
    defparam \POWERLED.count_off_7_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_7_LC_11_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_7_LC_11_10_7  (
            .in0(N__19363),
            .in1(N__17423),
            .in2(_gnd_net_),
            .in3(N__17328),
            .lcout(\POWERLED.count_offZ0Z_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_6 ),
            .carryout(\POWERLED.un1_count_off_1_cry_7 ),
            .clk(N__19155),
            .ce(N__18477),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_8_LC_11_11_0 .C_ON=1'b1;
    defparam \POWERLED.count_off_8_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_8_LC_11_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_8_LC_11_11_0  (
            .in0(N__19359),
            .in1(N__17822),
            .in2(_gnd_net_),
            .in3(N__17325),
            .lcout(\POWERLED.count_offZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\POWERLED.un1_count_off_1_cry_8 ),
            .clk(N__19212),
            .ce(N__18481),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_9_LC_11_11_1 .C_ON=1'b1;
    defparam \POWERLED.count_off_9_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_9_LC_11_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_9_LC_11_11_1  (
            .in0(N__19366),
            .in1(N__17835),
            .in2(_gnd_net_),
            .in3(N__17463),
            .lcout(\POWERLED.count_offZ0Z_9 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_8 ),
            .carryout(\POWERLED.un1_count_off_1_cry_9 ),
            .clk(N__19212),
            .ce(N__18481),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_10_LC_11_11_2 .C_ON=1'b1;
    defparam \POWERLED.count_off_10_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_10_LC_11_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_10_LC_11_11_2  (
            .in0(N__19356),
            .in1(N__17802),
            .in2(_gnd_net_),
            .in3(N__17460),
            .lcout(\POWERLED.count_offZ0Z_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_9 ),
            .carryout(\POWERLED.un1_count_off_1_cry_10 ),
            .clk(N__19212),
            .ce(N__18481),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_11_LC_11_11_3 .C_ON=1'b1;
    defparam \POWERLED.count_off_11_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_11_LC_11_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_11_LC_11_11_3  (
            .in0(N__19364),
            .in1(N__17774),
            .in2(_gnd_net_),
            .in3(N__17457),
            .lcout(\POWERLED.count_offZ0Z_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_10 ),
            .carryout(\POWERLED.un1_count_off_1_cry_11 ),
            .clk(N__19212),
            .ce(N__18481),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_12_LC_11_11_4 .C_ON=1'b1;
    defparam \POWERLED.count_off_12_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_12_LC_11_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_12_LC_11_11_4  (
            .in0(N__19357),
            .in1(N__17742),
            .in2(_gnd_net_),
            .in3(N__17454),
            .lcout(\POWERLED.count_offZ0Z_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_11 ),
            .carryout(\POWERLED.un1_count_off_1_cry_12 ),
            .clk(N__19212),
            .ce(N__18481),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_13_LC_11_11_5 .C_ON=1'b1;
    defparam \POWERLED.count_off_13_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_13_LC_11_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_13_LC_11_11_5  (
            .in0(N__19365),
            .in1(N__17754),
            .in2(_gnd_net_),
            .in3(N__17451),
            .lcout(\POWERLED.count_offZ0Z_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_12 ),
            .carryout(\POWERLED.un1_count_off_1_cry_13 ),
            .clk(N__19212),
            .ce(N__18481),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_14_LC_11_11_6 .C_ON=1'b1;
    defparam \POWERLED.count_off_14_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_14_LC_11_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_14_LC_11_11_6  (
            .in0(N__19358),
            .in1(N__17789),
            .in2(_gnd_net_),
            .in3(N__17448),
            .lcout(\POWERLED.count_offZ0Z_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_13 ),
            .carryout(\POWERLED.un1_count_off_1_cry_14 ),
            .clk(N__19212),
            .ce(N__18481),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_15_LC_11_11_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_15_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_15_LC_11_11_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \POWERLED.count_off_15_LC_11_11_7  (
            .in0(N__17729),
            .in1(N__19360),
            .in2(_gnd_net_),
            .in3(N__17445),
            .lcout(\POWERLED.count_offZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19212),
            .ce(N__18481),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIS3P11_2_LC_11_12_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIS3P11_2_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIS3P11_2_LC_11_12_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \POWERLED.count_off_RNIS3P11_2_LC_11_12_0  (
            .in0(N__19427),
            .in1(N__17442),
            .in2(N__17427),
            .in3(N__17409),
            .lcout(),
            .ltout(\POWERLED.func_state_ns_0_a2_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIIKVR3_10_LC_11_12_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIIKVR3_10_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIIKVR3_10_LC_11_12_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.count_off_RNIIKVR3_10_LC_11_12_1  (
            .in0(N__17700),
            .in1(N__17760),
            .in2(N__17394),
            .in3(N__17808),
            .lcout(\POWERLED.count_off_RNIIKVR3Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI8GP11_5_LC_11_12_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI8GP11_5_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI8GP11_5_LC_11_12_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \POWERLED.count_off_RNI8GP11_5_LC_11_12_2  (
            .in0(N__19397),
            .in1(N__17834),
            .in2(N__17823),
            .in3(N__19271),
            .lcout(\POWERLED.func_state_ns_0_a2_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI4D6S_10_LC_11_12_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI4D6S_10_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI4D6S_10_LC_11_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI4D6S_10_LC_11_12_3  (
            .in0(N__17801),
            .in1(N__17790),
            .in2(N__17775),
            .in3(N__17860),
            .lcout(\POWERLED.func_state_ns_0_a2_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIAJ6S_15_LC_11_12_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIAJ6S_15_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIAJ6S_15_LC_11_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNIAJ6S_15_LC_11_12_6  (
            .in0(N__17753),
            .in1(N__17741),
            .in2(N__17730),
            .in3(N__17715),
            .lcout(\POWERLED.func_state_ns_0_a2_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIJKKQ_LC_11_13_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIJKKQ_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIJKKQ_LC_11_13_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNIJKKQ_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__17694),
            .in2(_gnd_net_),
            .in3(N__17675),
            .lcout(vpp_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_LC_12_5_5 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_LC_12_5_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_LC_12_5_5  (
            .in0(N__18023),
            .in1(N__17593),
            .in2(_gnd_net_),
            .in3(N__17557),
            .lcout(\ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_RNIUU4I2_0_LC_12_6_0 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_RNIUU4I2_0_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_RNIUU4I2_0_LC_12_6_0 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_RNIUU4I2_0_LC_12_6_0  (
            .in0(N__18015),
            .in1(N__17591),
            .in2(_gnd_net_),
            .in3(N__17556),
            .lcout(\ALL_SYS_PWRGD.un1_curr_state10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_RNIV07U_10_LC_12_7_0 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_RNIV07U_10_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_RNIV07U_10_LC_12_7_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \ALL_SYS_PWRGD.count_RNIV07U_10_LC_12_7_0  (
            .in0(N__17513),
            .in1(N__17501),
            .in2(N__17490),
            .in3(N__17474),
            .lcout(),
            .ltout(\ALL_SYS_PWRGD.un4_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_12_7_1 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_12_7_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_12_7_1  (
            .in0(N__17943),
            .in1(N__18123),
            .in2(N__18249),
            .in3(N__18180),
            .lcout(\ALL_SYS_PWRGD.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_12_7_3 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_12_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_12_7_3  (
            .in0(N__18230),
            .in1(N__18218),
            .in2(N__18207),
            .in3(N__18191),
            .lcout(\ALL_SYS_PWRGD.un4_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_RNI027U_11_LC_12_7_5 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_RNI027U_11_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_RNI027U_11_LC_12_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ALL_SYS_PWRGD.count_RNI027U_11_LC_12_7_5  (
            .in0(N__18173),
            .in1(N__18161),
            .in2(N__18150),
            .in3(N__18134),
            .lcout(\ALL_SYS_PWRGD.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_1_LC_12_7_6 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_1_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_1_LC_12_7_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_1_LC_12_7_6  (
            .in0(N__18117),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18093),
            .lcout(),
            .ltout(\ALL_SYS_PWRGD.m4_0_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_LC_12_7_7 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_LC_12_7_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_LC_12_7_7  (
            .in0(N__18087),
            .in1(N__18075),
            .in2(N__18042),
            .in3(N__18039),
            .lcout(\ALL_SYS_PWRGD.N_245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_12_8_3 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_12_8_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_12_8_3  (
            .in0(N__17993),
            .in1(N__17981),
            .in2(N__17970),
            .in3(N__17954),
            .lcout(\ALL_SYS_PWRGD.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_12_8_4 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_12_8_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_12_8_4  (
            .in0(N__17925),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18740),
            .lcout(\ALL_SYS_PWRGD.N_49_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_0_LC_12_10_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_0_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_0_LC_12_10_0 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \POWERLED.count_off_0_LC_12_10_0  (
            .in0(N__19367),
            .in1(N__19296),
            .in2(N__17862),
            .in3(N__17880),
            .lcout(\POWERLED.count_offZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19232),
            .ce(N__18490),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_2_LC_12_10_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_2_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_2_LC_12_10_1 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \POWERLED.count_off_2_LC_12_10_1  (
            .in0(N__19297),
            .in1(N__19434),
            .in2(N__19428),
            .in3(N__19369),
            .lcout(\POWERLED.count_offZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19232),
            .ce(N__18490),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_5_LC_12_10_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_5_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_5_LC_12_10_3 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \POWERLED.count_off_5_LC_12_10_3  (
            .in0(N__19298),
            .in1(N__19404),
            .in2(N__19398),
            .in3(N__19370),
            .lcout(\POWERLED.count_offZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19232),
            .ce(N__18490),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_6_LC_12_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_6_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_6_LC_12_10_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \POWERLED.count_off_6_LC_12_10_4  (
            .in0(N__19368),
            .in1(N__19299),
            .in2(N__19272),
            .in3(N__19278),
            .lcout(\POWERLED.count_offZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19232),
            .ce(N__18490),
            .sr(_gnd_net_));
endmodule // TOP
