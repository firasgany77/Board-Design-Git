-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 11 2022 18:28:00

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VCCST_ENn : out std_logic;
    GPIO_FPGA_PM_3 : in std_logic;
    GPIO_FPGA_PCH_2 : in std_logic;
    VR_READY_VCCINAUX : in std_logic;
    VCCST_OK : in std_logic;
    VCCIO_EN : out std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    GPIO_FPGA_SV_4 : in std_logic;
    GPIO_FPGA_PM_4 : in std_logic;
    VDDQ_EN : out std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    GPIO_FPGA_PCH_4 : in std_logic;
    VCCIO_OK : in std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    SLP_SUSn : in std_logic;
    MAIN_12V_MON : in std_logic;
    GPIO_FPGA_SV_3 : in std_logic;
    GPIO_FPGA_HDR_3 : in std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    PLTRSTn : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    GPIO_FPGA_SV_1 : in std_logic;
    GPIO_FPGA_HDR_1 : in std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    V105A_EN : out std_logic;
    SYS_PWROK : out std_logic;
    GPIO_FPGA_PM_2 : in std_logic;
    GPIO_FPGA_PCH_1 : in std_logic;
    HDA_SDO_FPGA : out std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SLP_S4n : in std_logic;
    GPIO_FPGA_PCH_3 : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    V1P8_OK : in std_logic;
    DSW_PWROK : out std_logic;
    PM_PWROK : in std_logic;
    GPIO_FPGA_SV_2 : in std_logic;
    GPIO_FPGA_PCH_5 : in std_logic;
    V5A_EN : out std_logic;
    FPGA_GPIO_WD : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_EN : out std_logic;
    V105A_OK : in std_logic;
    SLP_S5n : in std_logic;
    GPIO_FPGA_HDR_2 : in std_logic;
    FP_RSTn : in std_logic;
    GPIO_FPGA_PM_1 : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__35653\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35623\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35615\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35532\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35515\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35453\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35399\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35033\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34951\ : std_logic;
signal \N__34948\ : std_logic;
signal \N__34945\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34891\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34396\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34230\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34145\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34055\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34036\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33952\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33863\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33813\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33004\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32809\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32803\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32791\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32707\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32608\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32441\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32066\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32038\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31974\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31943\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31901\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31318\ : std_logic;
signal \N__31315\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31141\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30934\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30805\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30301\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30085\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29801\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29197\ : std_logic;
signal \N__29194\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28888\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28739\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28697\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28581\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28301\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28277\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27383\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27314\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26374\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26112\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25620\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25604\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24334\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \b2v_inst16.count_4_3\ : std_logic;
signal \b2v_inst16.count_4_5\ : std_logic;
signal \bfn_1_2_0_\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_1\ : std_logic;
signal \b2v_inst16.countZ0Z_3\ : std_logic;
signal \b2v_inst16.count_rst_8\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_2_cZ0\ : std_logic;
signal \b2v_inst16.countZ0Z_4\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_3\ : std_logic;
signal \b2v_inst16.countZ0Z_5\ : std_logic;
signal \b2v_inst16.count_rst_10\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_4\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_5\ : std_logic;
signal \b2v_inst16.countZ0Z_7\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_6\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_7\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_8\ : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_9\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_10_cZ0\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_11\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_12\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_13\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_14\ : std_logic;
signal \b2v_inst16.count_rst_7\ : std_logic;
signal \b2v_inst16.count_4_2\ : std_logic;
signal \b2v_inst16.count_rst_1\ : std_logic;
signal \b2v_inst16.count_4_12\ : std_logic;
signal \b2v_inst16.count_rst_0\ : std_logic;
signal \b2v_inst16.count_4_11\ : std_logic;
signal \b2v_inst16.count_rst_11\ : std_logic;
signal \b2v_inst16.count_4_6\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_12_cascade_\ : std_logic;
signal \b2v_inst200.count_RNIC03N_3Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst200.count_RNI_0_0_cascade_\ : std_logic;
signal \b2v_inst200.count_2_11\ : std_logic;
signal \b2v_inst200.count_2_10\ : std_logic;
signal \b2v_inst200.count_2_8\ : std_logic;
signal \b2v_inst200.count_2_0\ : std_logic;
signal \b2v_inst200.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_13\ : std_logic;
signal \b2v_inst200.count_2_6\ : std_logic;
signal \b2v_inst200.count_2_14\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_10\ : std_logic;
signal \b2v_inst200.count_2_3\ : std_logic;
signal \b2v_inst200.count_2_4\ : std_logic;
signal \b2v_inst200.count_2_5\ : std_logic;
signal \b2v_inst200.count_2_9\ : std_logic;
signal \b2v_inst200.countZ0Z_9_cascade_\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_9\ : std_logic;
signal \b2v_inst200.count_2_12\ : std_logic;
signal \b2v_inst200.count_2_13\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_1\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_2\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_3\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_4\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_6\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_7_cZ0\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_8_cZ0\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_9_cZ0\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_10_cZ0\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_11\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_12\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_13\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_14\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0\ : std_logic;
signal \b2v_inst11.count_clk_0_15\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_6\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_8\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_7\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_9\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_4\ : std_logic;
signal \b2v_inst11.count_off_1_2\ : std_logic;
signal \b2v_inst11.count_offZ0Z_2\ : std_logic;
signal \b2v_inst11.count_off_1_2_cascade_\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_1_cascade_\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_0\ : std_logic;
signal \b2v_inst11.count_off_0_5\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_axb_2\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_1\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_2_cZ0\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_3_cZ0\ : std_logic;
signal \b2v_inst11.count_offZ0Z_5\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_4_cZ0\ : std_logic;
signal \b2v_inst11.un3_count_off_1_axb_6\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_5\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_6\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_7\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_8\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_9\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_10\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_11\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_12\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_13\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_14\ : std_logic;
signal \b2v_inst11.count_off_1_3_cascade_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_axb_3\ : std_logic;
signal \b2v_inst11.count_offZ0Z_4\ : std_logic;
signal \b2v_inst11.count_off_1_3\ : std_logic;
signal \b2v_inst11.count_offZ0Z_4_cascade_\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_2\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362\ : std_logic;
signal \b2v_inst11.count_offZ0Z_3\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672\ : std_logic;
signal \b2v_inst11.count_off_0_4\ : std_logic;
signal \b2v_inst11.count_off_0_14\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5\ : std_logic;
signal \b2v_inst16.count_rst_12\ : std_logic;
signal \b2v_inst16.count_4_7\ : std_logic;
signal \b2v_inst16.count_rst_9\ : std_logic;
signal \b2v_inst16.count_4_4\ : std_logic;
signal \b2v_inst16.count_rst_6_cascade_\ : std_logic;
signal \b2v_inst16.count_rst_6\ : std_logic;
signal \b2v_inst16.countZ0Z_11\ : std_logic;
signal \b2v_inst16.countZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst16.un4_count_1_axb_1\ : std_logic;
signal \b2v_inst16.count_4_1\ : std_logic;
signal \b2v_inst16.countZ0Z_2\ : std_logic;
signal \b2v_inst16.countZ0Z_6\ : std_logic;
signal \b2v_inst16.countZ0Z_12\ : std_logic;
signal \b2v_inst16.un13_clk_100khz_9\ : std_logic;
signal \b2v_inst16.un13_clk_100khz_8\ : std_logic;
signal \b2v_inst16.un13_clk_100khz_10_cascade_\ : std_logic;
signal \b2v_inst16.un13_clk_100khz_i_cascade_\ : std_logic;
signal \b2v_inst16.count_4_0\ : std_logic;
signal \b2v_inst16.count_rst_5_cascade_\ : std_logic;
signal \b2v_inst16.count_4_13\ : std_logic;
signal \b2v_inst16.count_rst_2\ : std_logic;
signal \b2v_inst16.countZ0Z_13\ : std_logic;
signal \b2v_inst16.countZ0Z_0\ : std_logic;
signal \b2v_inst16.countZ0Z_13_cascade_\ : std_logic;
signal \b2v_inst16.un13_clk_100khz_11\ : std_logic;
signal \b2v_inst16.countZ0Z_15\ : std_logic;
signal \b2v_inst16.count_rst_4\ : std_logic;
signal \b2v_inst16.count_4_15\ : std_logic;
signal \b2v_inst16.count_4_14\ : std_logic;
signal \b2v_inst16.count_rst_3\ : std_logic;
signal \b2v_inst16.countZ0Z_14\ : std_logic;
signal \b2v_inst200.count_2_15\ : std_logic;
signal \b2v_inst200.count_2_7\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_11\ : std_logic;
signal \b2v_inst200.count_0_16\ : std_logic;
signal \b2v_inst200.count_0_17\ : std_logic;
signal \b2v_inst200.count_2_1\ : std_logic;
signal \b2v_inst200.count_2_2\ : std_logic;
signal \b2v_inst200.count_en_g\ : std_logic;
signal \b2v_inst200.countZ0Z_0\ : std_logic;
signal \b2v_inst200.count_1_0\ : std_logic;
signal \bfn_2_6_0_\ : std_logic;
signal \b2v_inst200.countZ0Z_1\ : std_logic;
signal \b2v_inst200.count_RNIC03N_5Z0Z_0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_1_cy\ : std_logic;
signal \b2v_inst200.countZ0Z_2\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst200.countZ0Z_3\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst200.countZ0Z_4\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst200.countZ0Z_5\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst200.countZ0Z_6\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_5\ : std_logic;
signal \b2v_inst200.countZ0Z_7\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_7\ : std_logic;
signal \b2v_inst200.countZ0Z_8\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_7_c_RNIP33EZ0\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal \b2v_inst200.countZ0Z_9\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_8\ : std_logic;
signal \b2v_inst200.countZ0Z_10\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_9_c_RNIR75EZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst200.countZ0Z_11\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_10_c_RNI3AZ0Z29\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst200.countZ0Z_12\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst200.countZ0Z_13\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst200.countZ0Z_14\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst200.countZ0Z_15\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_15\ : std_logic;
signal \b2v_inst200.countZ0Z_16\ : std_logic;
signal \b2v_inst200.count_1_16\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \b2v_inst200.countZ0Z_17\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_16\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AAZ0\ : std_logic;
signal \b2v_inst11.count_clk_0_11\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_0_0\ : std_logic;
signal \b2v_inst11.count_clk_0_10\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_10\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_11\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_10_cascade_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_15\ : std_logic;
signal \b2v_inst11.un2_count_clk_17_0_o2_1_4_cascade_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_14\ : std_logic;
signal \b2v_inst11.count_clk_0_13\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CAZ0\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_13\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DAZ0\ : std_logic;
signal \b2v_inst11.count_clk_0_14\ : std_logic;
signal \b2v_inst11.count_clk_en_cascade_\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_2\ : std_logic;
signal \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_\ : std_logic;
signal \b2v_inst11.N_373\ : std_logic;
signal \b2v_inst11.N_373_cascade_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_8\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_6\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_4\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_2\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_3\ : std_logic;
signal \b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_7\ : std_logic;
signal \b2v_inst11.count_clk_RNIZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_en_0\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_12\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BAZ0\ : std_logic;
signal \b2v_inst11.count_clk_0_12\ : std_logic;
signal \b2v_inst11.count_clk_RNI_0Z0Z_0\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_0\ : std_logic;
signal \b2v_inst11.count_clk_0_1\ : std_logic;
signal \b2v_inst11.count_clk_RNIZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_5\ : std_logic;
signal \b2v_inst11.N_187\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_9\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_1\ : std_logic;
signal \b2v_inst11.count_clk_RNIZ0Z_5\ : std_logic;
signal \b2v_inst11.N_172\ : std_logic;
signal \b2v_inst11.N_421\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_i_1\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_0_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNICC5V2_0_1\ : std_logic;
signal \b2v_inst11.count_off_1_11_cascade_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_axb_11\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_12\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_4_cascade_\ : std_logic;
signal \b2v_inst11.count_off_0_12\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5\ : std_logic;
signal \b2v_inst11.count_offZ0Z_12\ : std_logic;
signal \b2v_inst11.count_off_1_11\ : std_logic;
signal \b2v_inst11.count_offZ0Z_11\ : std_logic;
signal \b2v_inst11.count_offZ0Z_12_cascade_\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_5\ : std_logic;
signal \b2v_inst11.count_offZ0Z_6\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2\ : std_logic;
signal \b2v_inst11.count_off_1_9\ : std_logic;
signal \b2v_inst11.count_off_1_9_cascade_\ : std_logic;
signal \b2v_inst11.count_offZ0Z_9\ : std_logic;
signal \b2v_inst11.un3_count_off_1_axb_9\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92\ : std_logic;
signal \b2v_inst11.count_off_1_6\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2\ : std_logic;
signal \b2v_inst11.count_off_0_15\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5\ : std_logic;
signal \b2v_inst11.count_offZ0Z_15\ : std_logic;
signal \b2v_inst11.count_offZ0Z_13\ : std_logic;
signal \b2v_inst11.count_offZ0Z_14\ : std_logic;
signal \b2v_inst11.count_offZ0Z_15_cascade_\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_11\ : std_logic;
signal \b2v_inst11.count_off_0_8\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2\ : std_logic;
signal \b2v_inst11.count_offZ0Z_8\ : std_logic;
signal \b2v_inst11.count_offZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_3\ : std_logic;
signal \b2v_inst11.count_offZ0Z_7\ : std_logic;
signal \b2v_inst11.count_off_1_7\ : std_logic;
signal \b2v_inst11.un3_count_off_1_axb_7\ : std_logic;
signal \bfn_4_1_0_\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_s_8_cascade_\ : std_logic;
signal \bfn_4_2_0_\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_i_0_8\ : std_logic;
signal \bfn_4_3_0_\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_7\ : std_logic;
signal \bfn_4_4_0_\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un40_sum_i_5_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_10\ : std_logic;
signal \b2v_inst16.count_rst\ : std_logic;
signal \b2v_inst16.count_4_10\ : std_logic;
signal \bfn_4_6_0_\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_5\ : std_logic;
signal \b2v_inst200.count_enZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_i_29\ : std_logic;
signal \b2v_inst11.mult1_un40_sum_i_l_ofx_4\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_s_4_sf\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_3\ : std_logic;
signal \b2v_inst11.count_clk_en\ : std_logic;
signal \b2v_inst11.N_150_N\ : std_logic;
signal \b2v_inst11.N_152_N_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_12_cascade_\ : std_logic;
signal \b2v_inst11.N_155_N_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_en_12\ : std_logic;
signal \b2v_inst11.dutycycle_en_12_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_15\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_12_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_10Z0Z_9_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_en_10\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_13\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_9_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_13_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_10_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIJU083Z0Z_8_cascade_\ : std_logic;
signal \b2v_inst11.N_108_f0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIHTFQZ0Z_8\ : std_logic;
signal \b2v_inst11.dutycycle_RNI2NK31Z0Z_8_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_e_1_8\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_8\ : std_logic;
signal \b2v_inst11.N_108_f0\ : std_logic;
signal \b2v_inst11.dutycycle_e_1_8_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIJU083_0Z0Z_8\ : std_logic;
signal \delayed_vccin_vccinaux_ok_RNIM6F44_0\ : std_logic;
signal \b2v_inst11.N_289_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_i_0_2_cascade_\ : std_logic;
signal \b2v_inst11.N_302_cascade_\ : std_logic;
signal \b2v_inst11.N_301_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIGKEF3Z0Z_12\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_12\ : std_logic;
signal \b2v_inst11.dutycycle_RNIGKEF3Z0Z_12_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_10_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_56_a0_3_0_cascade_\ : std_logic;
signal \b2v_inst11.N_232_N\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_325_N_cascade_\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_323_N\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_324_N\ : std_logic;
signal \b2v_inst11.N_322\ : std_logic;
signal \b2v_inst11.count_offZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_offZ0Z_1\ : std_logic;
signal \b2v_inst11.count_off_RNIZ0Z_1\ : std_logic;
signal \b2v_inst11.count_off_RNIZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.count_off_0_1\ : std_logic;
signal \b2v_inst11.count_offZ0Z_0\ : std_logic;
signal \b2v_inst11.count_off_0_0\ : std_logic;
signal \b2v_inst11.count_off_0_10\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2\ : std_logic;
signal \b2v_inst11.count_offZ0Z_10\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5\ : std_logic;
signal \b2v_inst11.count_off_0_13\ : std_logic;
signal \b2v_inst11.count_off_enZ0\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2\ : std_logic;
signal \bfn_5_1_0_\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_i_0_8\ : std_logic;
signal \bfn_5_2_0_\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_s_8\ : std_logic;
signal \bfn_5_4_0_\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_2_c\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_3_c\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_4_c\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_5_c\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_6_c\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_i_0_8\ : std_logic;
signal \bfn_5_5_0_\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_7\ : std_logic;
signal \bfn_5_6_0_\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_l_fx_3\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_l_fx_6\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_s_6\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un40_sum_i_5\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_i_8\ : std_logic;
signal \b2v_inst11.m15_e_2\ : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_0_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_1_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_2_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_3_cZ0\ : std_logic;
signal \b2v_inst11.mult1_un110_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_4_cZ0\ : std_logic;
signal \b2v_inst11.mult1_un103_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_5_cZ0\ : std_logic;
signal \b2v_inst11.mult1_un96_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_6_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_7_cZ0\ : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal \b2v_inst11.mult1_un82_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_8_cZ0\ : std_logic;
signal \b2v_inst11.mult1_un75_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_9_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_10\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_11\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_12\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_13\ : std_logic;
signal \b2v_inst11.mult1_un47_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_15\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \b2v_inst11.CO2\ : std_logic;
signal \b2v_inst11.CO2_THRU_CO\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_10\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_15\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_44_0_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_6Z0Z_9_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_11\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_15\ : std_logic;
signal \b2v_inst11.un1_m7_1_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_i3_mux\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_11\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_44_0_2_tz\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_39_0_0_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_39_0_0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_39_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_41_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_13\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_5Z0Z_9_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_10_1_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_12\ : std_logic;
signal \b2v_inst11.m18_i_1_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_11Z0Z_9\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_5Z0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_5Z0Z_9\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_8Z0Z_9\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_11\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_13_1\ : std_logic;
signal \b2v_inst11.G_6_i_0_cascade_\ : std_logic;
signal \b2v_inst11.G_6_i_a4_1_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_7_1\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_11\ : std_logic;
signal \b2v_inst11.dutycycle_RNIGKEF3Z0Z_11\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_8_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_11\ : std_logic;
signal \b2v_inst11.N_354\ : std_logic;
signal \b2v_inst11.N_354_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_11\ : std_logic;
signal \b2v_inst11.g2_1_1\ : std_logic;
signal \b2v_inst11.g3_0_1_cascade_\ : std_logic;
signal \b2v_inst11.N_14_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_6Z0Z_5\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_6Z0Z_5_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_RNI_0Z0Z_1\ : std_logic;
signal \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_0_0\ : std_logic;
signal \b2v_inst11.N_122\ : std_logic;
signal \b2v_inst11.N_357\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_a2_0\ : std_logic;
signal \b2v_inst11.N_327\ : std_logic;
signal \b2v_inst11.N_328\ : std_logic;
signal \b2v_inst11.func_state_1_m0_0_0_0_cascade_\ : std_logic;
signal \bfn_6_1_0_\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_s_8_cascade_\ : std_logic;
signal \bfn_6_2_0_\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_i_0_8\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_axb_4_l_fx\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_axb_7_l_fx\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un68_sum\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un117_sum\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un124_sum\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un89_sum\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_s_8\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un54_sum\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un61_sum\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_s_8\ : std_logic;
signal \b2v_inst16.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst16.curr_state_7_0_cascade_\ : std_logic;
signal \b2v_inst16.un13_clk_100khz_i\ : std_logic;
signal \b2v_inst16.curr_state_0_1\ : std_logic;
signal \b2v_inst16.delayed_vddq_pwrgdZ0\ : std_logic;
signal b2v_inst16_un2_vpp_en_0_i : std_logic;
signal \b2v_inst16.curr_state_1_0\ : std_logic;
signal \b2v_inst16.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst16.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_0\ : std_logic;
signal \b2v_inst200.count_RNIC03N_3Z0Z_0\ : std_logic;
signal \V105A_EN_c\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_5\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_10\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_5\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_14\ : std_logic;
signal \b2v_inst11.dutycycle_en_11\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_13_cascade_\ : std_logic;
signal \b2v_inst11.un2_count_clk_17_0_a2_1_4\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_4\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_50_a4_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_10\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_7\ : std_logic;
signal \VCCST_OK_c\ : std_logic;
signal \VDDQ_OK_c\ : std_logic;
signal \VCCIO_EN_c\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_3\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_7_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_9\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIAI7C4Z0Z_4_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_eena_2_0_1\ : std_logic;
signal \b2v_inst11.func_state_RNI3JFN6Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI3JFN6Z0Z_4\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_4\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_9\ : std_logic;
signal \b2v_inst11.func_state_RNI3JFN6Z0Z_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI0KJ31Z0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI74A23Z0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_e_1_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNI74A23Z0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_e_1_7_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI01TT1Z0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNI25OT3Z0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNIGALV4Z0Z_0\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNIGSFQZ0Z_7\ : std_logic;
signal \bfn_6_13_0_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_0_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDUZ0Z8\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_2\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_3\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_4\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_5_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_6_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_7_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHPZ0Z49\ : std_logic;
signal \bfn_6_14_0_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_2\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_8_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_9_cZ0\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_7\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNPZ0Z5\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_10\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_10\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQZ0Z5\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_11\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_9\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_12\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_13\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_12\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_5Z0Z_5_cascade_\ : std_logic;
signal \b2v_inst11.N_156\ : std_logic;
signal \b2v_inst11.N_156_cascade_\ : std_logic;
signal \b2v_inst11.N_331\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_307_N\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_5Z0Z_5\ : std_logic;
signal \b2v_inst11.N_4_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNI_0Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNINJ641_0Z0Z_0\ : std_logic;
signal \b2v_inst11.func_state_RNINJ641_0Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_off_RNIQCBN4Z0Z_9_cascade_\ : std_logic;
signal \b2v_inst11.N_333\ : std_logic;
signal \b2v_inst11.func_state_RNI_1Z0Z_1\ : std_logic;
signal \b2v_inst11.func_state_1_m2s2_i_1\ : std_logic;
signal \b2v_inst11.N_73\ : std_logic;
signal \b2v_inst11.func_state_1_m0_0\ : std_logic;
signal \b2v_inst11.N_73_cascade_\ : std_logic;
signal \b2v_inst11.count_off_RNIQCBN4Z0Z_9\ : std_logic;
signal \b2v_inst11.func_state_1_m0_1\ : std_logic;
signal \bfn_7_2_0_\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_i_0_8\ : std_logic;
signal \bfn_7_3_0_\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un138_sum\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un131_sum\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_i\ : std_logic;
signal \b2v_inst11.un1_count_cry_0_i\ : std_logic;
signal \bfn_7_5_0_\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1\ : std_logic;
signal \b2v_inst11.N_5647_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_0\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_2\ : std_logic;
signal \b2v_inst11.N_5648_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_1\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_3\ : std_logic;
signal \b2v_inst11.N_5649_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_2\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_4\ : std_logic;
signal \b2v_inst11.N_5650_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_3\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_5\ : std_logic;
signal \b2v_inst11.N_5651_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_4\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_6\ : std_logic;
signal \b2v_inst11.N_5652_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_5\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_7\ : std_logic;
signal \b2v_inst11.N_5653_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_6\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_7\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_8\ : std_logic;
signal \b2v_inst11.N_5654_i\ : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_9\ : std_logic;
signal \b2v_inst11.N_5655_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_8\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_10\ : std_logic;
signal \b2v_inst11.N_5656_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_9\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_11\ : std_logic;
signal \b2v_inst11.N_5657_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_10\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_12\ : std_logic;
signal \b2v_inst11.N_5658_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_11\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_13\ : std_logic;
signal \b2v_inst11.N_5659_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_12\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_14\ : std_logic;
signal \b2v_inst11.N_5660_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_13\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_i_8\ : std_logic;
signal \b2v_inst11.N_5661_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_14\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_15_cZ0\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \b2v_inst36.curr_state_RNI8TT2Z0Z_0\ : std_logic;
signal \b2v_inst11.pwm_out_en_cascade_\ : std_logic;
signal \PWRBTN_LED_c\ : std_logic;
signal \b2v_inst11.pwm_out_1_sqmuxa_0\ : std_logic;
signal \b2v_inst11.curr_state_0_0\ : std_logic;
signal \b2v_inst11.curr_state_3_0\ : std_logic;
signal \b2v_inst11.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_0_sqmuxa_i_cascade_\ : std_logic;
signal \b2v_inst11.N_349\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_32_and_i_o2_0_0_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNIAI7C4Z0Z_10_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_5\ : std_logic;
signal \b2v_inst11.N_418\ : std_logic;
signal \b2v_inst11.func_state_RNIJU083Z0Z_0\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_43_and_i_o2_0_0_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJTZ0Z69\ : std_logic;
signal \b2v_inst11.dutycycle_RNI4I3C2Z0Z_10\ : std_logic;
signal \b2v_inst11.dutycycle_RNI4I3C2Z0Z_10_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIAI7C4Z0Z_10\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_10\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_5\ : std_logic;
signal \b2v_inst11.d_i3_mux_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_5\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_3\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_3\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8\ : std_logic;
signal \b2v_inst11.dutycycle_e_1_3\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_3\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_6_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_5Z0Z_3\ : std_logic;
signal \b2v_inst11.func_state_RNINJ641_0Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.g0_2_3\ : std_logic;
signal \b2v_inst11.g0_2_2\ : std_logic;
signal \b2v_inst11.g0_1_1_0\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_2_i_o3_out\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_1\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_1_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNI_1Z0Z_0\ : std_logic;
signal \b2v_inst11.func_state_RNI_0Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_func_state25_4_i_a2_1_cascade_\ : std_logic;
signal \b2v_inst11.N_321\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIZ0\ : std_logic;
signal \b2v_inst11.g1\ : std_logic;
signal \b2v_inst11.dutycycle_0_6\ : std_logic;
signal \b2v_inst11.g1_cascade_\ : std_logic;
signal \b2v_inst11.g1_0\ : std_logic;
signal \b2v_inst11.dutycycle_eena\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_0\ : std_logic;
signal \b2v_inst11.dutycycle_eena_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_0\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_sx\ : std_logic;
signal \b2v_inst11.func_state_RNI_0Z0Z_1\ : std_logic;
signal \b2v_inst11.func_state_1_m0_0_0_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_0\ : std_logic;
signal \b2v_inst11.N_360\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.func_stateZ0Z_0\ : std_logic;
signal \b2v_inst11.func_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.N_3013_i_cascade_\ : std_logic;
signal \b2v_inst11.N_330\ : std_logic;
signal \b2v_inst11.func_state_RNI_0Z0Z_0\ : std_logic;
signal \b2v_inst11.g1_1\ : std_logic;
signal \b2v_inst11.func_state_RNI673P9Z0Z_0\ : std_logic;
signal \b2v_inst11.func_stateZ1Z_0\ : std_logic;
signal \b2v_inst11.count_off_RNIZ0Z_9\ : std_logic;
signal \b2v_inst11.N_335_cascade_\ : std_logic;
signal \b2v_inst11.count_off_RNIQ1RAS1Z0Z_9\ : std_logic;
signal \b2v_inst11.func_state_1_ss0_i_0_o2_0\ : std_logic;
signal \b2v_inst36.count_rst_11_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst36.count_1_7\ : std_logic;
signal \b2v_inst36.count_rst_9_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_5_cascade_\ : std_logic;
signal \b2v_inst36.count_1_5\ : std_logic;
signal \b2v_inst36.count_rst_7\ : std_logic;
signal \b2v_inst36.count_rst_6_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst36.count_1_8\ : std_logic;
signal \b2v_inst36.count_rst_4_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_10_cascade_\ : std_logic;
signal \b2v_inst36.count_1_10\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_i_0_8\ : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_1\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_axb_7\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_i_0_8\ : std_logic;
signal \b2v_inst11.count_0_14\ : std_logic;
signal \b2v_inst11.count_0_6\ : std_logic;
signal \b2v_inst11.count_0_15\ : std_logic;
signal \b2v_inst11.count_0_7\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \b2v_inst11.un1_count_cry_1\ : std_logic;
signal \b2v_inst11.un1_count_cry_2\ : std_logic;
signal \b2v_inst11.un1_count_cry_3\ : std_logic;
signal \b2v_inst11.un1_count_cry_4\ : std_logic;
signal \b2v_inst11.un1_count_cry_5_c_RNIMQUDZ0\ : std_logic;
signal \b2v_inst11.un1_count_cry_5\ : std_logic;
signal \b2v_inst11.un1_count_cry_6_c_RNINSVDZ0\ : std_logic;
signal \b2v_inst11.un1_count_cry_6\ : std_logic;
signal \b2v_inst11.un1_count_cry_7\ : std_logic;
signal \b2v_inst11.un1_count_cry_8\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \b2v_inst11.un1_count_cry_9\ : std_logic;
signal \b2v_inst11.un1_count_cry_10\ : std_logic;
signal \b2v_inst11.un1_count_cry_11\ : std_logic;
signal \b2v_inst11.un1_count_cry_12\ : std_logic;
signal \b2v_inst11.un1_count_cry_13_c_RNI5AUZ0Z6\ : std_logic;
signal \b2v_inst11.un1_count_cry_13\ : std_logic;
signal \b2v_inst11.un1_count_cry_14\ : std_logic;
signal \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6\ : std_logic;
signal \b2v_inst11.un1_count_cry_9_c_RNIQ23EZ0\ : std_logic;
signal \b2v_inst11.count_0_10\ : std_logic;
signal \b2v_inst11.un1_count_cry_10_c_RNI24RZ0Z6\ : std_logic;
signal \b2v_inst11.count_0_11\ : std_logic;
signal \b2v_inst11.un1_count_cry_1_c_RNIIIQDZ0\ : std_logic;
signal \b2v_inst11.count_0_2\ : std_logic;
signal \b2v_inst11.un1_count_cry_11_c_RNI36SZ0Z6\ : std_logic;
signal \b2v_inst11.count_0_12\ : std_logic;
signal \G_2727_cascade_\ : std_logic;
signal \b2v_inst5.curr_state_2_1\ : std_logic;
signal \N_229_cascade_\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \curr_state_RNI5VS71_0_1_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un145_sum\ : std_logic;
signal \RSMRSTn_RNI8DFE_cascade_\ : std_logic;
signal \b2v_inst11.g0_1_1\ : std_logic;
signal \b2v_inst11.N_182\ : std_logic;
signal \b2v_inst11.func_state_RNIT4D71_0Z0Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_0_5\ : std_logic;
signal \b2v_inst11.g1_4_0\ : std_logic;
signal \b2v_inst11.func_state_RNIT4D71_0Z0Z_1_cascade_\ : std_logic;
signal \dutycycle_RNIIOE3D_0_5_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_5_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_3_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_2\ : std_logic;
signal \b2v_inst11.un1_i3_mux_1\ : std_logic;
signal \b2v_inst11.g0_6_2\ : std_logic;
signal \b2v_inst11.m15_e_3\ : std_logic;
signal \b2v_inst11.un1_dutycycle_inv_4_0\ : std_logic;
signal \b2v_inst11.g0_9_1\ : std_logic;
signal \b2v_inst11.g1_0_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_164_0\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_5\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_i\ : std_logic;
signal \b2v_inst11.N_3013_i\ : std_logic;
signal \b2v_inst11.N_221_iZ0\ : std_logic;
signal \b2v_inst11.func_state_cascade_\ : std_logic;
signal \b2v_inst11.N_303_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_eena_1\ : std_logic;
signal \b2v_inst11.N_70\ : std_logic;
signal \b2v_inst11.dutycycle_eena_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_2\ : std_logic;
signal \b2v_inst11.dutycycle_eena_0\ : std_logic;
signal \b2v_inst11.N_169\ : std_logic;
signal \b2v_inst11.N_375\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_sxZ0_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_47keep_fast\ : std_logic;
signal \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_1\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_26_and_i_o2_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNINJ641_0Z0Z_5\ : std_logic;
signal \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_cascade_\ : std_logic;
signal \b2v_inst11.N_183\ : std_logic;
signal \b2v_inst11.func_state_RNI_3Z0Z_1\ : std_logic;
signal \b2v_inst11.N_183_cascade_\ : std_logic;
signal \b2v_inst11.N_114_f0_1\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_6\ : std_logic;
signal \b2v_inst11.N_379\ : std_logic;
signal \b2v_inst6.curr_state_RNI8OKQ2Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_52_and_i_a2Z0Z_1\ : std_logic;
signal \b2v_inst11.func_state_RNIDINH9Z0Z_0\ : std_logic;
signal \b2v_inst11.func_stateZ0Z_1\ : std_logic;
signal \b2v_inst6.curr_state_RNI8OKQ2Z0Z_0\ : std_logic;
signal \b2v_inst6.delayed_vccin_vccinaux_ok_0\ : std_logic;
signal \SYNTHESIZED_WIRE_49_i_0_o3_0\ : std_logic;
signal \VPP_OK_c\ : std_logic;
signal \VDDQ_EN_c\ : std_logic;
signal \VCCIO_OK_c\ : std_logic;
signal \V5S_OK_c\ : std_logic;
signal \b2v_inst31.un8_outputZ0Z_0\ : std_logic;
signal \V33S_OK_c\ : std_logic;
signal \VCCIN_EN_c\ : std_logic;
signal \bfn_9_1_0_\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst36.countZ0Z_5\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_5\ : std_logic;
signal \b2v_inst36.countZ0Z_7\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_7\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_8\ : std_logic;
signal \bfn_9_2_0_\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_9_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst36.count_1_12\ : std_logic;
signal \b2v_inst36.count_en_cascade_\ : std_logic;
signal \b2v_inst36.count_rst_2\ : std_logic;
signal \b2v_inst36.count_rst_0\ : std_logic;
signal \b2v_inst36.count_1_14\ : std_logic;
signal \b2v_inst36.count_rst\ : std_logic;
signal \b2v_inst36.count_1_15\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_0\ : std_logic;
signal \bfn_9_4_0_\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_0\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_2_s\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_1\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_s_7\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_3\ : std_logic;
signal \G_2890\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_axb_6\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_5\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0\ : std_logic;
signal \b2v_inst11.dutycycle\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_i\ : std_logic;
signal \b2v_inst11.countZ0Z_2\ : std_logic;
signal \b2v_inst11.countZ0Z_7\ : std_logic;
signal \b2v_inst11.countZ0Z_15\ : std_logic;
signal \b2v_inst11.countZ0Z_11\ : std_logic;
signal \b2v_inst11.countZ0Z_10\ : std_logic;
signal \b2v_inst11.countZ0Z_12\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlt6\ : std_logic;
signal \b2v_inst11.countZ0Z_6\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlto15_5_cascade_\ : std_logic;
signal \b2v_inst11.countZ0Z_14\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlto15_7_cascade_\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlto15_4\ : std_logic;
signal \b2v_inst11.count_RNIZ0Z_13\ : std_logic;
signal \b2v_inst11.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst11.count_RNIZ0Z_13_cascade_\ : std_logic;
signal \b2v_inst11.countZ0Z_3\ : std_logic;
signal \b2v_inst11.un1_count_cry_2_c_RNIJKRDZ0\ : std_logic;
signal \b2v_inst11.count_0_3\ : std_logic;
signal \b2v_inst11.countZ0Z_13\ : std_logic;
signal \b2v_inst11.un1_count_cry_12_c_RNI48TZ0Z6\ : std_logic;
signal \b2v_inst11.count_0_13\ : std_logic;
signal \b2v_inst11.countZ0Z_4\ : std_logic;
signal \b2v_inst11.un1_count_cry_3_c_RNIKMSDZ0\ : std_logic;
signal \b2v_inst11.count_0_4\ : std_logic;
signal \b2v_inst11.countZ0Z_5\ : std_logic;
signal \b2v_inst11.un1_count_cry_4_c_RNILOTDZ0\ : std_logic;
signal \b2v_inst11.count_0_5\ : std_logic;
signal \b2v_inst11.count_0_0\ : std_logic;
signal \b2v_inst11.count_RNI_2_0\ : std_logic;
signal \b2v_inst11.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_RNIZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.countZ0Z_1\ : std_logic;
signal \b2v_inst11.countZ0Z_0\ : std_logic;
signal \b2v_inst11.countZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.count_0_sqmuxa_i\ : std_logic;
signal \b2v_inst11.count_0_1\ : std_logic;
signal \b2v_inst11.countZ0Z_8\ : std_logic;
signal \b2v_inst11.un1_count_cry_7_c_RNIOU0EZ0\ : std_logic;
signal \b2v_inst11.count_0_8\ : std_logic;
signal \b2v_inst11.countZ0Z_9\ : std_logic;
signal \b2v_inst11.un1_count_cry_8_c_RNIP02EZ0\ : std_logic;
signal \b2v_inst11.count_0_9\ : std_logic;
signal \b2v_inst5.curr_state_3_0\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_0\ : std_logic;
signal \G_2727\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst5.m4_0\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_4\ : std_logic;
signal \b2v_inst11.dutycycle_RNITBKN1Z0Z_7\ : std_logic;
signal \N_229\ : std_logic;
signal \b2v_inst5.count_enZ0_cascade_\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO\ : std_logic;
signal \b2v_inst11.g0_2_1\ : std_logic;
signal \b2v_inst11.pwm_outZ0\ : std_logic;
signal \b2v_inst11.pwm_out_1_sqmuxa\ : std_logic;
signal \b2v_inst20.un4_counter_0_and\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \b2v_inst20.un4_counter_0\ : std_logic;
signal \b2v_inst20.un4_counter_1\ : std_logic;
signal \b2v_inst20.un4_counter_2\ : std_logic;
signal \b2v_inst20.un4_counter_3\ : std_logic;
signal \b2v_inst20.un4_counter_4\ : std_logic;
signal \b2v_inst20.un4_counter_5\ : std_logic;
signal \b2v_inst20.un4_counter_6\ : std_logic;
signal b2v_inst20_un4_counter_7 : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \b2v_inst20.un4_counter_1_and\ : std_logic;
signal \curr_state_RNI5VS71_0_1\ : std_logic;
signal \RSMRSTn_0\ : std_logic;
signal \b2v_inst11.N_234_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_52_and_i_0_0_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_47keep_rep1\ : std_logic;
signal \b2v_inst20_un4_counter_7_THRU_CO\ : std_logic;
signal \dutycycle_RNIIOE3D_0_5\ : std_logic;
signal b2v_inst11_count_off_1_sqmuxa_0_0_0 : std_logic;
signal \G_26_0_a5_1_0\ : std_logic;
signal \G_26_0_a5_2_1_cascade_\ : std_logic;
signal \G_26_0_0\ : std_logic;
signal \b2v_inst11.g2_0_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_172_m4\ : std_logic;
signal \b2v_inst11_un1_dutycycle_172_m3_0_0_0_cascade_\ : std_logic;
signal \b2v_inst11.g2_1\ : std_logic;
signal \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z2\ : std_logic;
signal \b2v_inst11.g4_cascade_\ : std_logic;
signal b2v_inst16_delayed_vddq_pwrgd_en : std_logic;
signal \b2v_inst11.N_5\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_xZ0\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_3\ : std_logic;
signal \b2v_inst11.N_12\ : std_logic;
signal \b2v_inst11.func_state_RNINJ641_0Z0Z_1\ : std_logic;
signal \N_4\ : std_logic;
signal \G_26_0_a5_2\ : std_logic;
signal \b2v_inst11.N_158\ : std_logic;
signal \b2v_inst11.N_3046_i\ : std_logic;
signal \b2v_inst11.g3_0\ : std_logic;
signal \b2v_inst11.g2_0_cascade_\ : std_logic;
signal \RSMRSTn_RNI8DFE\ : std_logic;
signal \b2v_inst11.N_228_N_0\ : std_logic;
signal \b2v_inst6.delayed_vccin_vccinaux_okZ0\ : std_logic;
signal \b2v_inst11.g1_4_2_0\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_8\ : std_logic;
signal \N_19_i\ : std_logic;
signal \b2v_inst11.g0_8_0_0\ : std_logic;
signal \SLP_S4n_c\ : std_logic;
signal \GPIO_FPGA_PCH_5_c\ : std_logic;
signal \b2v_inst11.func_state\ : std_logic;
signal \SLP_S3n_c\ : std_logic;
signal \b2v_inst11.count_clk_RNIZ0Z_3\ : std_logic;
signal \b2v_inst11.g1_2_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_6\ : std_logic;
signal \b2v_inst11.g1_2\ : std_logic;
signal \b2v_inst6.countZ0Z_11_cascade_\ : std_logic;
signal \b2v_inst6.count_3_11\ : std_logic;
signal \b2v_inst6.curr_state_RNIDMSJ1Z0Z_1\ : std_logic;
signal \b2v_inst6.count_rst_10\ : std_logic;
signal \b2v_inst6.count_rst_3_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_4_cascade_\ : std_logic;
signal \b2v_inst6.count_3_4\ : std_logic;
signal \G_2746_cascade_\ : std_logic;
signal \b2v_inst6.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst6.curr_state_2_0\ : std_logic;
signal \VR_READY_VCCIN_c\ : std_logic;
signal \VR_READY_VCCINAUX_c\ : std_logic;
signal \SYNTHESIZED_WIRE_48_i_0_o3_2\ : std_logic;
signal \b2v_inst6.N_413_cascade_\ : std_logic;
signal \b2v_inst6.curr_state_7_1_cascade_\ : std_logic;
signal \b2v_inst6.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst6.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst6.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst6.N_413\ : std_logic;
signal \b2v_inst6.curr_state_1_1\ : std_logic;
signal \b2v_inst36.countZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst36.count_rst_13\ : std_logic;
signal \b2v_inst36.countZ0Z_14\ : std_logic;
signal \b2v_inst36.countZ0Z_15\ : std_logic;
signal \b2v_inst36.count_1_1\ : std_logic;
signal \b2v_inst36.count_rst_12_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_2\ : std_logic;
signal \b2v_inst36.countZ0Z_2_cascade_\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_1_THRU_CO\ : std_logic;
signal \b2v_inst36.count_1_2\ : std_logic;
signal \b2v_inst36.countZ0Z_3\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst36.count_1_3\ : std_logic;
signal \b2v_inst36.countZ0Z_8\ : std_logic;
signal \b2v_inst36.countZ0Z_10\ : std_logic;
signal \b2v_inst36.countZ0Z_1\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_11\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_10_cascade_\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_8\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_6\ : std_logic;
signal \b2v_inst36.count_rst_3\ : std_logic;
signal \b2v_inst36.countZ0Z_11\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \b2v_inst36.countZ0Z_11_cascade_\ : std_logic;
signal \b2v_inst36.count_1_11\ : std_logic;
signal \b2v_inst36.count_rst_8\ : std_logic;
signal \b2v_inst36.count_1_6\ : std_logic;
signal \b2v_inst36.countZ0Z_12\ : std_logic;
signal \b2v_inst36.countZ0Z_6_cascade_\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_9\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst36.curr_state_7_0_cascade_\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst36.DSW_PWROK_0\ : std_logic;
signal \b2v_inst36.curr_state_3_1\ : std_logic;
signal \b2v_inst36.curr_state_7_1\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst36.curr_state_4_0\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_1\ : std_logic;
signal \V33DSW_OK_c\ : std_logic;
signal \b2v_inst36.N_2925_i\ : std_logic;
signal \b2v_inst5.count_0_14\ : std_logic;
signal \b2v_inst5.count_0_7\ : std_logic;
signal \b2v_inst16.countZ0Z_8\ : std_logic;
signal \b2v_inst16.count_rst_13\ : std_logic;
signal \b2v_inst16.count_4_8\ : std_logic;
signal \b2v_inst16.countZ0Z_9\ : std_logic;
signal \b2v_inst16.count_rst_14\ : std_logic;
signal \b2v_inst16.count_4_9\ : std_logic;
signal \b2v_inst16.count_en\ : std_logic;
signal \b2v_inst36.count_1_4\ : std_logic;
signal \b2v_inst36.count_rst_10\ : std_logic;
signal \b2v_inst36.countZ0Z_4\ : std_logic;
signal \b2v_inst5.N_2906_i_cascade_\ : std_logic;
signal \b2v_inst5.count_1_i_a2_1_0_cascade_\ : std_logic;
signal \b2v_inst5.count_0_12\ : std_logic;
signal \b2v_inst5.count_1_i_a2_0_0\ : std_logic;
signal \b2v_inst5.count_0_5\ : std_logic;
signal \b2v_inst5.count_0_6\ : std_logic;
signal \b2v_inst5.count_1_i_a2_2_0\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_5\ : std_logic;
signal \b2v_inst5.count_rst_9\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_6\ : std_logic;
signal \b2v_inst5.count_rst_8\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_5\ : std_logic;
signal \b2v_inst5.countZ0Z_7\ : std_logic;
signal \b2v_inst5.count_rst_7\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_7\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_8\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_12\ : std_logic;
signal \b2v_inst5.count_rst_2\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst5.countZ0Z_14\ : std_logic;
signal \b2v_inst5.count_rst_0\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst5.countZ0Z_15\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst5.count_rst\ : std_logic;
signal \b2v_inst5.count_0_15\ : std_logic;
signal \b2v_inst20.counterZ0Z_1\ : std_logic;
signal \b2v_inst20.counterZ0Z_0\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \b2v_inst20.counterZ0Z_2\ : std_logic;
signal \b2v_inst20.counter_1_cry_1_THRU_CO\ : std_logic;
signal \b2v_inst20.counter_1_cry_1\ : std_logic;
signal \b2v_inst20.counterZ0Z_3\ : std_logic;
signal \b2v_inst20.counter_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst20.counter_1_cry_2\ : std_logic;
signal \b2v_inst20.counterZ0Z_4\ : std_logic;
signal \b2v_inst20.counter_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst20.counter_1_cry_3\ : std_logic;
signal \b2v_inst20.counterZ0Z_5\ : std_logic;
signal \b2v_inst20.counter_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst20.counter_1_cry_4\ : std_logic;
signal \b2v_inst20.counterZ0Z_6\ : std_logic;
signal \b2v_inst20.counter_1_cry_5_THRU_CO\ : std_logic;
signal \b2v_inst20.counter_1_cry_5\ : std_logic;
signal \b2v_inst20.counterZ0Z_7\ : std_logic;
signal \b2v_inst20.counter_1_cry_6\ : std_logic;
signal \b2v_inst20.counter_1_cry_7\ : std_logic;
signal \b2v_inst20.counter_1_cry_8\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \b2v_inst20.counter_1_cry_9\ : std_logic;
signal \b2v_inst20.counter_1_cry_10\ : std_logic;
signal \b2v_inst20.counter_1_cry_11\ : std_logic;
signal \b2v_inst20.counter_1_cry_12\ : std_logic;
signal \b2v_inst20.counter_1_cry_13\ : std_logic;
signal \b2v_inst20.counter_1_cry_14\ : std_logic;
signal \b2v_inst20.counter_1_cry_15\ : std_logic;
signal \b2v_inst20.counter_1_cry_16\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \b2v_inst20.counter_1_cry_17\ : std_logic;
signal \b2v_inst20.counter_1_cry_18\ : std_logic;
signal \b2v_inst20.counter_1_cry_19\ : std_logic;
signal \b2v_inst20.counter_1_cry_20\ : std_logic;
signal \b2v_inst20.counter_1_cry_21\ : std_logic;
signal \b2v_inst20.counter_1_cry_22\ : std_logic;
signal \b2v_inst20.counter_1_cry_23\ : std_logic;
signal \b2v_inst20.counter_1_cry_24\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \b2v_inst20.counter_1_cry_25\ : std_logic;
signal \b2v_inst20.counter_1_cry_26\ : std_logic;
signal \b2v_inst20.counter_1_cry_27\ : std_logic;
signal \b2v_inst20.counter_1_cry_28\ : std_logic;
signal \b2v_inst20.counter_1_cry_29\ : std_logic;
signal \b2v_inst20.counter_1_cry_30\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_5\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_7\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_8\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst6.count_rst_4_cascade_\ : std_logic;
signal \b2v_inst6.count_3_5\ : std_logic;
signal \b2v_inst6.count_rst_2_cascade_\ : std_logic;
signal \b2v_inst6.count_rst_8_cascade_\ : std_logic;
signal \b2v_inst6.count_rst_9\ : std_logic;
signal \b2v_inst6.count_3_10\ : std_logic;
signal \b2v_inst6.countZ0Z_11\ : std_logic;
signal \b2v_inst6.count_rst_6_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_7\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \b2v_inst6.countZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst6.count_3_7\ : std_logic;
signal \b2v_inst6.count_rst_7_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_8\ : std_logic;
signal \b2v_inst6.countZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst6.count_3_8\ : std_logic;
signal \b2v_inst6.countZ0Z_9\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \b2v_inst6.count_3_9\ : std_logic;
signal \b2v_inst36.N_2928_i_cascade_\ : std_logic;
signal \b2v_inst36.count_1_13\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_12_c_RNIS7LZ0Z1\ : std_logic;
signal \b2v_inst36.countZ0Z_13\ : std_logic;
signal \b2v_inst36.countZ0Z_9\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_8_c_RNIH8IZ0Z8\ : std_logic;
signal \b2v_inst36.count_1_9\ : std_logic;
signal \b2v_inst36.count_rst_14\ : std_logic;
signal \b2v_inst36.countZ0Z_0\ : std_logic;
signal \b2v_inst36.N_2928_i\ : std_logic;
signal \b2v_inst36.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst36.N_1_i\ : std_logic;
signal \b2v_inst36.count_1_0\ : std_logic;
signal \b2v_inst36.count_en\ : std_logic;
signal \b2v_inst36.count_0_sqmuxa\ : std_logic;
signal \b2v_inst5.count_rst_5\ : std_logic;
signal \b2v_inst5.count_rst_5_cascade_\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_9\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_9_cascade_\ : std_logic;
signal \b2v_inst5.count_0_9\ : std_logic;
signal \b2v_inst5.count_rst_4_cascade_\ : std_logic;
signal \b2v_inst5.countZ0Z_10\ : std_logic;
signal \b2v_inst5.countZ0Z_10_cascade_\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_9_THRU_CO\ : std_logic;
signal \b2v_inst5.count_0_10\ : std_logic;
signal \b2v_inst5.count_RNIRHC7IZ0Z_2_cascade_\ : std_logic;
signal \b2v_inst5.countZ0Z_0\ : std_logic;
signal \b2v_inst5.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst5.count_RNIZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst5.count_RNIZ0Z_0\ : std_logic;
signal \b2v_inst5.count_0_1\ : std_logic;
signal \b2v_inst5.count_1_i_a2_11_0\ : std_logic;
signal \b2v_inst5.N_2906_i\ : std_logic;
signal \b2v_inst5.count_0_0\ : std_logic;
signal \b2v_inst5.count_0_3\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9\ : std_logic;
signal \b2v_inst5.countZ0Z_3\ : std_logic;
signal \b2v_inst5.count_1_i_a2_6_0\ : std_logic;
signal \b2v_inst5.count_1_i_a2_4_0_cascade_\ : std_logic;
signal \b2v_inst5.count_1_i_a2_12_0\ : std_logic;
signal \b2v_inst5.count_0_2\ : std_logic;
signal \b2v_inst5.count_rst_12\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_2\ : std_logic;
signal \b2v_inst5.countZ0Z_1\ : std_logic;
signal \b2v_inst5.count_1_i_a2_3_0\ : std_logic;
signal \b2v_inst5.count_0_11\ : std_logic;
signal \b2v_inst5.count_rst_3\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_11\ : std_logic;
signal \b2v_inst5.count_1_i_a2_5_0\ : std_logic;
signal \b2v_inst5.count_rst_6_cascade_\ : std_logic;
signal \b2v_inst5.countZ0Z_8\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst5.countZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst5.count_0_8\ : std_logic;
signal \b2v_inst5.count_rst_10\ : std_logic;
signal \b2v_inst5.count_rst_10_cascade_\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_4\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_4_cascade_\ : std_logic;
signal \b2v_inst5.count_0_4\ : std_logic;
signal \b2v_inst5.N_390\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_12_THRU_CO\ : std_logic;
signal \b2v_inst5.count_0_sqmuxa\ : std_logic;
signal \b2v_inst5.count_enZ0\ : std_logic;
signal \b2v_inst5.count_rst_1_cascade_\ : std_logic;
signal \b2v_inst5.count_0_13\ : std_logic;
signal \b2v_inst5.countZ0Z_13\ : std_logic;
signal \b2v_inst20.counterZ0Z_11\ : std_logic;
signal \b2v_inst20.counterZ0Z_8\ : std_logic;
signal \b2v_inst20.counterZ0Z_10\ : std_logic;
signal \b2v_inst20.counterZ0Z_9\ : std_logic;
signal \b2v_inst20.un4_counter_2_and\ : std_logic;
signal \b2v_inst20.counterZ0Z_12\ : std_logic;
signal \b2v_inst20.counterZ0Z_14\ : std_logic;
signal \b2v_inst20.counterZ0Z_15\ : std_logic;
signal \b2v_inst20.counterZ0Z_13\ : std_logic;
signal \b2v_inst20.un4_counter_3_and\ : std_logic;
signal \b2v_inst20.counterZ0Z_19\ : std_logic;
signal \b2v_inst20.counterZ0Z_16\ : std_logic;
signal \b2v_inst20.counterZ0Z_17\ : std_logic;
signal \b2v_inst20.counterZ0Z_18\ : std_logic;
signal \b2v_inst20.un4_counter_4_and\ : std_logic;
signal \b2v_inst20.counterZ0Z_23\ : std_logic;
signal \b2v_inst20.counterZ0Z_22\ : std_logic;
signal \b2v_inst20.counterZ0Z_21\ : std_logic;
signal \b2v_inst20.counterZ0Z_20\ : std_logic;
signal \b2v_inst20.un4_counter_5_and\ : std_logic;
signal \b2v_inst20.counterZ0Z_24\ : std_logic;
signal \b2v_inst20.counterZ0Z_27\ : std_logic;
signal \b2v_inst20.counterZ0Z_25\ : std_logic;
signal \b2v_inst20.counterZ0Z_26\ : std_logic;
signal \b2v_inst20.un4_counter_6_and\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \N_405\ : std_logic;
signal \GPIO_FPGA_PCH_1_c\ : std_logic;
signal \b2v_inst200.count_RNI_0_0\ : std_logic;
signal \N_405_cascade_\ : std_logic;
signal \b2v_inst200.m6_i_0_cascade_\ : std_logic;
signal \b2v_inst200.N_57_cascade_\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \N_406_cascade_\ : std_logic;
signal \b2v_inst200.N_55\ : std_logic;
signal \N_406\ : std_logic;
signal \b2v_inst200.curr_state_0_1\ : std_logic;
signal \b2v_inst200.N_202_cascade_\ : std_logic;
signal \HDA_SDO_FPGA_c\ : std_logic;
signal \b2v_inst20.counterZ0Z_29\ : std_logic;
signal \b2v_inst20.counterZ0Z_28\ : std_logic;
signal \b2v_inst20.counterZ0Z_31\ : std_logic;
signal \b2v_inst20.counterZ0Z_30\ : std_logic;
signal \b2v_inst20.un4_counter_7_and\ : std_logic;
signal \b2v_inst200.m11_0_a3_0\ : std_logic;
signal \b2v_inst200.N_202\ : std_logic;
signal \G_2788\ : std_logic;
signal \b2v_inst200.curr_state_0_2\ : std_logic;
signal \G_2788_cascade_\ : std_logic;
signal \SYNTHESIZED_WIRE_47keep\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_2\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_2_cascade_\ : std_logic;
signal \b2v_inst200.HDA_SDO_FPGA_0\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_1\ : std_logic;
signal \N_219\ : std_logic;
signal \b2v_inst200.m6_i_0\ : std_logic;
signal \b2v_inst200.curr_state_0_0\ : std_logic;
signal b2v_inst16_delayed_vddq_pwrgd_en_g : std_logic;
signal \b2v_inst6.count_rst_0_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst6.count_3_1\ : std_logic;
signal \b2v_inst6.count_rst_1\ : std_logic;
signal \b2v_inst6.count_3_2\ : std_logic;
signal \b2v_inst6.count_3_6\ : std_logic;
signal \b2v_inst6.count_rst_5\ : std_logic;
signal \b2v_inst6.countZ0Z_6\ : std_logic;
signal \b2v_inst6.countZ0Z_10\ : std_logic;
signal \b2v_inst6.countZ0Z_2\ : std_logic;
signal \b2v_inst6.countZ0Z_6_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_1\ : std_logic;
signal \b2v_inst6.countZ0Z_12\ : std_logic;
signal \b2v_inst6.count_rst_11\ : std_logic;
signal \b2v_inst6.count_3_12\ : std_logic;
signal \b2v_inst6.countZ0Z_13\ : std_logic;
signal \b2v_inst6.count_rst_12\ : std_logic;
signal \b2v_inst6.count_3_13\ : std_logic;
signal \b2v_inst6.countZ0Z_14\ : std_logic;
signal \b2v_inst6.count_rst_13\ : std_logic;
signal \b2v_inst6.count_3_14\ : std_logic;
signal \b2v_inst6.count_3_15\ : std_logic;
signal \b2v_inst6.count_rst_14\ : std_logic;
signal \b2v_inst6.countZ0Z_15\ : std_logic;
signal \V5A_OK_c\ : std_logic;
signal \V33A_OK_c\ : std_logic;
signal \V1P8A_OK_c\ : std_logic;
signal \V105A_OK_c\ : std_logic;
signal \SYNTHESIZED_WIRE_26\ : std_logic;
signal \b2v_inst6.count_rst_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst6.count_3_0\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst6.count_3_3\ : std_logic;
signal \FPGA_OSC_0_c_g\ : std_logic;
signal \b2v_inst6.count_en\ : std_logic;
signal \b2v_inst6.count_0_sqmuxa\ : std_logic;
signal \b2v_inst6.countZ0Z_5\ : std_logic;
signal \b2v_inst6.countZ0Z_3\ : std_logic;
signal \b2v_inst6.countZ0Z_4\ : std_logic;
signal \b2v_inst6.countZ0Z_0\ : std_logic;
signal \b2v_inst6.un12_clk_100khz_10\ : std_logic;
signal \b2v_inst6.un12_clk_100khz_9\ : std_logic;
signal \b2v_inst6.un12_clk_100khz_11_cascade_\ : std_logic;
signal \b2v_inst6.un12_clk_100khz_8\ : std_logic;
signal \b2v_inst6.N_1_i\ : std_logic;
signal \b2v_inst6.N_1_i_cascade_\ : std_logic;
signal \b2v_inst6.N_1_i_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \FPGA_OSC_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \HDA_SDO_FPGA_wire\ : std_logic;
signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \VCCIO_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \V105A_EN_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \VCCST_ENn_wire\ : std_logic;
signal \VCCST_OK_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \GPIO_FPGA_PCH_5_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \V105A_OK_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \GPIO_FPGA_PCH_1_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \VCCIO_EN_wire\ : std_logic;

begin
    \FPGA_OSC_wire\ <= FPGA_OSC;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \V5A_OK_wire\ <= V5A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V5S_ENn <= \V5S_ENn_wire\;
    \SLP_S4n_wire\ <= SLP_S4n;
    HDA_SDO_FPGA <= \HDA_SDO_FPGA_wire\;
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    \SLP_S3n_wire\ <= SLP_S3n;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    \VPP_OK_wire\ <= VPP_OK;
    V33A_ENn <= \V33A_ENn_wire\;
    \V5S_OK_wire\ <= V5S_OK;
    \V33A_OK_wire\ <= V33A_OK;
    VPP_EN <= \VPP_EN_wire\;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \VCCIO_OK_wire\ <= VCCIO_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    RSMRSTn <= \RSMRSTn_wire\;
    V105A_EN <= \V105A_EN_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    VCCST_ENn <= \VCCST_ENn_wire\;
    \VCCST_OK_wire\ <= VCCST_OK;
    DSW_PWROK <= \DSW_PWROK_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \GPIO_FPGA_PCH_5_wire\ <= GPIO_FPGA_PCH_5;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \V105A_OK_wire\ <= V105A_OK;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \GPIO_FPGA_PCH_1_wire\ <= GPIO_FPGA_PCH_1;
    V5A_EN <= \V5A_EN_wire\;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    VCCIO_EN <= \VCCIO_EN_wire\;

    \FPGA_OSC_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__35651\,
            GLOBALBUFFEROUTPUT => \FPGA_OSC_0_c_g\
        );

    \FPGA_OSC_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35653\,
            DIN => \N__35652\,
            DOUT => \N__35651\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \FPGA_OSC_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35653\,
            PADOUT => \N__35652\,
            PADIN => \N__35651\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V1P8A_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35642\,
            DIN => \N__35641\,
            DOUT => \N__35640\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \V1P8A_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35642\,
            PADOUT => \N__35641\,
            PADIN => \N__35640\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V1P8A_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V5A_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35633\,
            DIN => \N__35632\,
            DOUT => \N__35631\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \V5A_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35633\,
            PADOUT => \N__35632\,
            PADIN => \N__35631\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V5A_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PCH_PWROK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35624\,
            DIN => \N__35623\,
            DOUT => \N__35622\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \PCH_PWROK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35624\,
            PADOUT => \N__35623\,
            PADIN => \N__35622\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17640\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCIN_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35615\,
            DIN => \N__35614\,
            DOUT => \N__35613\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \VCCIN_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35615\,
            PADOUT => \N__35614\,
            PADIN => \N__35613\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24954\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33S_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35606\,
            DIN => \N__35605\,
            DOUT => \N__35604\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \V33S_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35606\,
            PADOUT => \N__35605\,
            PADIN => \N__35604\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V33S_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V5S_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35597\,
            DIN => \N__35596\,
            DOUT => \N__35595\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \V5S_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35597\,
            PADOUT => \N__35596\,
            PADIN => \N__35595\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29685\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SLP_S4n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35588\,
            DIN => \N__35587\,
            DOUT => \N__35586\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \SLP_S4n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35588\,
            PADOUT => \N__35587\,
            PADIN => \N__35586\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SLP_S4n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HDA_SDO_FPGA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35579\,
            DIN => \N__35578\,
            DOUT => \N__35577\,
            PACKAGEPIN => \HDA_SDO_FPGA_wire\
        );

    \HDA_SDO_FPGA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35579\,
            PADOUT => \N__35578\,
            PADIN => \N__35577\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33505\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VR_READY_VCCINAUX_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35570\,
            DIN => \N__35569\,
            DOUT => \N__35568\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \VR_READY_VCCINAUX_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35570\,
            PADOUT => \N__35569\,
            PADIN => \N__35568\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VR_READY_VCCINAUX_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SLP_S3n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35561\,
            DIN => \N__35560\,
            DOUT => \N__35559\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \SLP_S3n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35561\,
            PADOUT => \N__35560\,
            PADIN => \N__35559\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SLP_S3n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCST_PWRGD_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35552\,
            DIN => \N__35551\,
            DOUT => \N__35550\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \VCCST_PWRGD_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35552\,
            PADOUT => \N__35551\,
            PADIN => \N__35550\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17625\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VPP_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35543\,
            DIN => \N__35542\,
            DOUT => \N__35541\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \VPP_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35543\,
            PADOUT => \N__35542\,
            PADIN => \N__35541\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VPP_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33A_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35534\,
            DIN => \N__35533\,
            DOUT => \N__35532\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \V33A_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35534\,
            PADOUT => \N__35533\,
            PADIN => \N__35532\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V5S_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35525\,
            DIN => \N__35524\,
            DOUT => \N__35523\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \V5S_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35525\,
            PADOUT => \N__35524\,
            PADIN => \N__35523\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V5S_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33A_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35516\,
            DIN => \N__35515\,
            DOUT => \N__35514\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \V33A_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35516\,
            PADOUT => \N__35515\,
            PADIN => \N__35514\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V33A_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VPP_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35507\,
            DIN => \N__35506\,
            DOUT => \N__35505\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \VPP_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35507\,
            PADOUT => \N__35506\,
            PADIN => \N__35505\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20290\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PWRBTN_LED_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35498\,
            DIN => \N__35497\,
            DOUT => \N__35496\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \PWRBTN_LED_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35498\,
            PADOUT => \N__35497\,
            PADIN => \N__35496\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22144\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCIO_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35489\,
            DIN => \N__35488\,
            DOUT => \N__35487\,
            PACKAGEPIN => \VCCIO_OK_wire\
        );

    \VCCIO_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35489\,
            PADOUT => \N__35488\,
            PADIN => \N__35487\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VCCIO_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33S_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35480\,
            DIN => \N__35479\,
            DOUT => \N__35478\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \V33S_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35480\,
            PADOUT => \N__35479\,
            PADIN => \N__35478\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29686\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RSMRSTn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35471\,
            DIN => \N__35470\,
            DOUT => \N__35469\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \RSMRSTn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35471\,
            PADOUT => \N__35470\,
            PADIN => \N__35469\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29119\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V105A_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35462\,
            DIN => \N__35461\,
            DOUT => \N__35460\,
            PACKAGEPIN => \V105A_EN_wire\
        );

    \V105A_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35462\,
            PADOUT => \N__35461\,
            PADIN => \N__35460\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20494\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V1P8A_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35453\,
            DIN => \N__35452\,
            DOUT => \N__35451\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \V1P8A_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35453\,
            PADOUT => \N__35452\,
            PADIN => \N__35451\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VDDQ_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35444\,
            DIN => \N__35443\,
            DOUT => \N__35442\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \VDDQ_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35444\,
            PADOUT => \N__35443\,
            PADIN => \N__35442\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VDDQ_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCST_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35435\,
            DIN => \N__35434\,
            DOUT => \N__35433\,
            PACKAGEPIN => \VCCST_ENn_wire\
        );

    \VCCST_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35435\,
            PADOUT => \N__35434\,
            PADIN => \N__35433\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25096\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCST_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35426\,
            DIN => \N__35425\,
            DOUT => \N__35424\,
            PACKAGEPIN => \VCCST_OK_wire\
        );

    \VCCST_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35426\,
            PADOUT => \N__35425\,
            PADIN => \N__35424\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VCCST_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DSW_PWROK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35417\,
            DIN => \N__35416\,
            DOUT => \N__35415\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \DSW_PWROK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35417\,
            PADOUT => \N__35416\,
            PADIN => \N__35415\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20493\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SYS_PWROK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35408\,
            DIN => \N__35407\,
            DOUT => \N__35406\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \SYS_PWROK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35408\,
            PADOUT => \N__35407\,
            PADIN => \N__35406\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17641\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO_FPGA_PCH_5_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35399\,
            DIN => \N__35398\,
            DOUT => \N__35397\,
            PACKAGEPIN => \GPIO_FPGA_PCH_5_wire\
        );

    \GPIO_FPGA_PCH_5_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35399\,
            PADOUT => \N__35398\,
            PADIN => \N__35397\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \GPIO_FPGA_PCH_5_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33DSW_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35390\,
            DIN => \N__35389\,
            DOUT => \N__35388\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \V33DSW_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35390\,
            PADOUT => \N__35389\,
            PADIN => \N__35388\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V33DSW_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V105A_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35381\,
            DIN => \N__35380\,
            DOUT => \N__35379\,
            PACKAGEPIN => \V105A_OK_wire\
        );

    \V105A_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35381\,
            PADOUT => \N__35380\,
            PADIN => \N__35379\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V105A_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VR_READY_VCCIN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35372\,
            DIN => \N__35371\,
            DOUT => \N__35370\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \VR_READY_VCCIN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35372\,
            PADOUT => \N__35371\,
            PADIN => \N__35370\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VR_READY_VCCIN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VDDQ_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35363\,
            DIN => \N__35362\,
            DOUT => \N__35361\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \VDDQ_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35363\,
            PADOUT => \N__35362\,
            PADIN => \N__35361\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24994\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO_FPGA_PCH_1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35354\,
            DIN => \N__35353\,
            DOUT => \N__35352\,
            PACKAGEPIN => \GPIO_FPGA_PCH_1_wire\
        );

    \GPIO_FPGA_PCH_1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__35354\,
            PADOUT => \N__35353\,
            PADIN => \N__35352\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \GPIO_FPGA_PCH_1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V5A_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35345\,
            DIN => \N__35344\,
            DOUT => \N__35343\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \V5A_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35345\,
            PADOUT => \N__35344\,
            PADIN => \N__35343\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20125\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCINAUX_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35336\,
            DIN => \N__35335\,
            DOUT => \N__35334\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \VCCINAUX_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35336\,
            PADOUT => \N__35335\,
            PADIN => \N__35334\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24955\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCIO_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35327\,
            DIN => \N__35326\,
            DOUT => \N__35325\,
            PACKAGEPIN => \VCCIO_EN_wire\
        );

    \VCCIO_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__35327\,
            PADOUT => \N__35326\,
            PADIN => \N__35325\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20605\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__8172\ : SRMux
    port map (
            O => \N__35308\,
            I => \N__35304\
        );

    \I__8171\ : SRMux
    port map (
            O => \N__35307\,
            I => \N__35301\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__35304\,
            I => \N__35298\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__35301\,
            I => \N__35285\
        );

    \I__8168\ : IoSpan4Mux
    port map (
            O => \N__35298\,
            I => \N__35285\
        );

    \I__8167\ : SRMux
    port map (
            O => \N__35297\,
            I => \N__35280\
        );

    \I__8166\ : InMux
    port map (
            O => \N__35296\,
            I => \N__35280\
        );

    \I__8165\ : SRMux
    port map (
            O => \N__35295\,
            I => \N__35267\
        );

    \I__8164\ : SRMux
    port map (
            O => \N__35294\,
            I => \N__35264\
        );

    \I__8163\ : InMux
    port map (
            O => \N__35293\,
            I => \N__35255\
        );

    \I__8162\ : InMux
    port map (
            O => \N__35292\,
            I => \N__35255\
        );

    \I__8161\ : InMux
    port map (
            O => \N__35291\,
            I => \N__35255\
        );

    \I__8160\ : InMux
    port map (
            O => \N__35290\,
            I => \N__35255\
        );

    \I__8159\ : Span4Mux_s1_v
    port map (
            O => \N__35285\,
            I => \N__35250\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__35280\,
            I => \N__35250\
        );

    \I__8157\ : InMux
    port map (
            O => \N__35279\,
            I => \N__35239\
        );

    \I__8156\ : InMux
    port map (
            O => \N__35278\,
            I => \N__35239\
        );

    \I__8155\ : InMux
    port map (
            O => \N__35277\,
            I => \N__35239\
        );

    \I__8154\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35239\
        );

    \I__8153\ : InMux
    port map (
            O => \N__35275\,
            I => \N__35239\
        );

    \I__8152\ : InMux
    port map (
            O => \N__35274\,
            I => \N__35234\
        );

    \I__8151\ : InMux
    port map (
            O => \N__35273\,
            I => \N__35234\
        );

    \I__8150\ : InMux
    port map (
            O => \N__35272\,
            I => \N__35229\
        );

    \I__8149\ : InMux
    port map (
            O => \N__35271\,
            I => \N__35229\
        );

    \I__8148\ : SRMux
    port map (
            O => \N__35270\,
            I => \N__35219\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__35267\,
            I => \N__35214\
        );

    \I__8146\ : LocalMux
    port map (
            O => \N__35264\,
            I => \N__35214\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__35255\,
            I => \N__35211\
        );

    \I__8144\ : Span4Mux_v
    port map (
            O => \N__35250\,
            I => \N__35206\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__35239\,
            I => \N__35206\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__35234\,
            I => \N__35196\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__35229\,
            I => \N__35196\
        );

    \I__8140\ : SRMux
    port map (
            O => \N__35228\,
            I => \N__35193\
        );

    \I__8139\ : InMux
    port map (
            O => \N__35227\,
            I => \N__35186\
        );

    \I__8138\ : InMux
    port map (
            O => \N__35226\,
            I => \N__35186\
        );

    \I__8137\ : InMux
    port map (
            O => \N__35225\,
            I => \N__35186\
        );

    \I__8136\ : InMux
    port map (
            O => \N__35224\,
            I => \N__35179\
        );

    \I__8135\ : InMux
    port map (
            O => \N__35223\,
            I => \N__35179\
        );

    \I__8134\ : InMux
    port map (
            O => \N__35222\,
            I => \N__35179\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__35219\,
            I => \N__35175\
        );

    \I__8132\ : Span4Mux_v
    port map (
            O => \N__35214\,
            I => \N__35168\
        );

    \I__8131\ : Span4Mux_v
    port map (
            O => \N__35211\,
            I => \N__35168\
        );

    \I__8130\ : Span4Mux_s1_v
    port map (
            O => \N__35206\,
            I => \N__35168\
        );

    \I__8129\ : InMux
    port map (
            O => \N__35205\,
            I => \N__35157\
        );

    \I__8128\ : InMux
    port map (
            O => \N__35204\,
            I => \N__35157\
        );

    \I__8127\ : InMux
    port map (
            O => \N__35203\,
            I => \N__35157\
        );

    \I__8126\ : InMux
    port map (
            O => \N__35202\,
            I => \N__35157\
        );

    \I__8125\ : InMux
    port map (
            O => \N__35201\,
            I => \N__35157\
        );

    \I__8124\ : Span4Mux_s2_h
    port map (
            O => \N__35196\,
            I => \N__35154\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__35193\,
            I => \N__35147\
        );

    \I__8122\ : LocalMux
    port map (
            O => \N__35186\,
            I => \N__35147\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__35179\,
            I => \N__35147\
        );

    \I__8120\ : InMux
    port map (
            O => \N__35178\,
            I => \N__35144\
        );

    \I__8119\ : Odrv4
    port map (
            O => \N__35175\,
            I => \b2v_inst6.count_0_sqmuxa\
        );

    \I__8118\ : Odrv4
    port map (
            O => \N__35168\,
            I => \b2v_inst6.count_0_sqmuxa\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__35157\,
            I => \b2v_inst6.count_0_sqmuxa\
        );

    \I__8116\ : Odrv4
    port map (
            O => \N__35154\,
            I => \b2v_inst6.count_0_sqmuxa\
        );

    \I__8115\ : Odrv4
    port map (
            O => \N__35147\,
            I => \b2v_inst6.count_0_sqmuxa\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__35144\,
            I => \b2v_inst6.count_0_sqmuxa\
        );

    \I__8113\ : InMux
    port map (
            O => \N__35131\,
            I => \N__35127\
        );

    \I__8112\ : CascadeMux
    port map (
            O => \N__35130\,
            I => \N__35122\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__35127\,
            I => \N__35119\
        );

    \I__8110\ : InMux
    port map (
            O => \N__35126\,
            I => \N__35116\
        );

    \I__8109\ : InMux
    port map (
            O => \N__35125\,
            I => \N__35113\
        );

    \I__8108\ : InMux
    port map (
            O => \N__35122\,
            I => \N__35110\
        );

    \I__8107\ : Span4Mux_v
    port map (
            O => \N__35119\,
            I => \N__35107\
        );

    \I__8106\ : LocalMux
    port map (
            O => \N__35116\,
            I => \N__35104\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__35113\,
            I => \b2v_inst6.countZ0Z_5\
        );

    \I__8104\ : LocalMux
    port map (
            O => \N__35110\,
            I => \b2v_inst6.countZ0Z_5\
        );

    \I__8103\ : Odrv4
    port map (
            O => \N__35107\,
            I => \b2v_inst6.countZ0Z_5\
        );

    \I__8102\ : Odrv4
    port map (
            O => \N__35104\,
            I => \b2v_inst6.countZ0Z_5\
        );

    \I__8101\ : CascadeMux
    port map (
            O => \N__35095\,
            I => \N__35089\
        );

    \I__8100\ : CascadeMux
    port map (
            O => \N__35094\,
            I => \N__35086\
        );

    \I__8099\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35083\
        );

    \I__8098\ : InMux
    port map (
            O => \N__35092\,
            I => \N__35080\
        );

    \I__8097\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35077\
        );

    \I__8096\ : InMux
    port map (
            O => \N__35086\,
            I => \N__35074\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__35083\,
            I => \N__35071\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__35080\,
            I => \b2v_inst6.countZ0Z_3\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__35077\,
            I => \b2v_inst6.countZ0Z_3\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__35074\,
            I => \b2v_inst6.countZ0Z_3\
        );

    \I__8091\ : Odrv4
    port map (
            O => \N__35071\,
            I => \b2v_inst6.countZ0Z_3\
        );

    \I__8090\ : CascadeMux
    port map (
            O => \N__35062\,
            I => \N__35059\
        );

    \I__8089\ : InMux
    port map (
            O => \N__35059\,
            I => \N__35055\
        );

    \I__8088\ : InMux
    port map (
            O => \N__35058\,
            I => \N__35051\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__35055\,
            I => \N__35048\
        );

    \I__8086\ : CascadeMux
    port map (
            O => \N__35054\,
            I => \N__35045\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__35051\,
            I => \N__35042\
        );

    \I__8084\ : Span4Mux_s3_h
    port map (
            O => \N__35048\,
            I => \N__35039\
        );

    \I__8083\ : InMux
    port map (
            O => \N__35045\,
            I => \N__35036\
        );

    \I__8082\ : Span4Mux_s2_h
    port map (
            O => \N__35042\,
            I => \N__35033\
        );

    \I__8081\ : Odrv4
    port map (
            O => \N__35039\,
            I => \b2v_inst6.countZ0Z_4\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__35036\,
            I => \b2v_inst6.countZ0Z_4\
        );

    \I__8079\ : Odrv4
    port map (
            O => \N__35033\,
            I => \b2v_inst6.countZ0Z_4\
        );

    \I__8078\ : CascadeMux
    port map (
            O => \N__35026\,
            I => \N__35022\
        );

    \I__8077\ : InMux
    port map (
            O => \N__35025\,
            I => \N__35017\
        );

    \I__8076\ : InMux
    port map (
            O => \N__35022\,
            I => \N__35013\
        );

    \I__8075\ : InMux
    port map (
            O => \N__35021\,
            I => \N__35008\
        );

    \I__8074\ : InMux
    port map (
            O => \N__35020\,
            I => \N__35008\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__35017\,
            I => \N__35005\
        );

    \I__8072\ : InMux
    port map (
            O => \N__35016\,
            I => \N__35002\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__35013\,
            I => \N__34999\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__35008\,
            I => \N__34996\
        );

    \I__8069\ : Odrv4
    port map (
            O => \N__35005\,
            I => \b2v_inst6.countZ0Z_0\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__35002\,
            I => \b2v_inst6.countZ0Z_0\
        );

    \I__8067\ : Odrv4
    port map (
            O => \N__34999\,
            I => \b2v_inst6.countZ0Z_0\
        );

    \I__8066\ : Odrv12
    port map (
            O => \N__34996\,
            I => \b2v_inst6.countZ0Z_0\
        );

    \I__8065\ : InMux
    port map (
            O => \N__34987\,
            I => \N__34984\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__34984\,
            I => \b2v_inst6.un12_clk_100khz_10\
        );

    \I__8063\ : InMux
    port map (
            O => \N__34981\,
            I => \N__34978\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__34978\,
            I => \N__34975\
        );

    \I__8061\ : Odrv4
    port map (
            O => \N__34975\,
            I => \b2v_inst6.un12_clk_100khz_9\
        );

    \I__8060\ : CascadeMux
    port map (
            O => \N__34972\,
            I => \b2v_inst6.un12_clk_100khz_11_cascade_\
        );

    \I__8059\ : InMux
    port map (
            O => \N__34969\,
            I => \N__34966\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__34966\,
            I => \N__34963\
        );

    \I__8057\ : Odrv4
    port map (
            O => \N__34963\,
            I => \b2v_inst6.un12_clk_100khz_8\
        );

    \I__8056\ : InMux
    port map (
            O => \N__34960\,
            I => \N__34954\
        );

    \I__8055\ : InMux
    port map (
            O => \N__34959\,
            I => \N__34954\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__34954\,
            I => \N__34951\
        );

    \I__8053\ : Span4Mux_h
    port map (
            O => \N__34951\,
            I => \N__34948\
        );

    \I__8052\ : Odrv4
    port map (
            O => \N__34948\,
            I => \b2v_inst6.N_1_i\
        );

    \I__8051\ : CascadeMux
    port map (
            O => \N__34945\,
            I => \b2v_inst6.N_1_i_cascade_\
        );

    \I__8050\ : InMux
    port map (
            O => \N__34942\,
            I => \N__34930\
        );

    \I__8049\ : InMux
    port map (
            O => \N__34941\,
            I => \N__34930\
        );

    \I__8048\ : InMux
    port map (
            O => \N__34940\,
            I => \N__34917\
        );

    \I__8047\ : InMux
    port map (
            O => \N__34939\,
            I => \N__34917\
        );

    \I__8046\ : InMux
    port map (
            O => \N__34938\,
            I => \N__34917\
        );

    \I__8045\ : InMux
    port map (
            O => \N__34937\,
            I => \N__34917\
        );

    \I__8044\ : InMux
    port map (
            O => \N__34936\,
            I => \N__34917\
        );

    \I__8043\ : InMux
    port map (
            O => \N__34935\,
            I => \N__34911\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__34930\,
            I => \N__34908\
        );

    \I__8041\ : CascadeMux
    port map (
            O => \N__34929\,
            I => \N__34905\
        );

    \I__8040\ : CascadeMux
    port map (
            O => \N__34928\,
            I => \N__34900\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__34917\,
            I => \N__34897\
        );

    \I__8038\ : InMux
    port map (
            O => \N__34916\,
            I => \N__34891\
        );

    \I__8037\ : InMux
    port map (
            O => \N__34915\,
            I => \N__34886\
        );

    \I__8036\ : InMux
    port map (
            O => \N__34914\,
            I => \N__34886\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__34911\,
            I => \N__34881\
        );

    \I__8034\ : Span4Mux_v
    port map (
            O => \N__34908\,
            I => \N__34881\
        );

    \I__8033\ : InMux
    port map (
            O => \N__34905\,
            I => \N__34872\
        );

    \I__8032\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34872\
        );

    \I__8031\ : InMux
    port map (
            O => \N__34903\,
            I => \N__34872\
        );

    \I__8030\ : InMux
    port map (
            O => \N__34900\,
            I => \N__34872\
        );

    \I__8029\ : Span4Mux_h
    port map (
            O => \N__34897\,
            I => \N__34869\
        );

    \I__8028\ : InMux
    port map (
            O => \N__34896\,
            I => \N__34862\
        );

    \I__8027\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34862\
        );

    \I__8026\ : InMux
    port map (
            O => \N__34894\,
            I => \N__34862\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__34891\,
            I => \b2v_inst6.N_1_i_i\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__34886\,
            I => \b2v_inst6.N_1_i_i\
        );

    \I__8023\ : Odrv4
    port map (
            O => \N__34881\,
            I => \b2v_inst6.N_1_i_i\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__34872\,
            I => \b2v_inst6.N_1_i_i\
        );

    \I__8021\ : Odrv4
    port map (
            O => \N__34869\,
            I => \b2v_inst6.N_1_i_i\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__34862\,
            I => \b2v_inst6.N_1_i_i\
        );

    \I__8019\ : InMux
    port map (
            O => \N__34849\,
            I => \N__34845\
        );

    \I__8018\ : InMux
    port map (
            O => \N__34848\,
            I => \N__34842\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__34845\,
            I => \b2v_inst6.countZ0Z_14\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__34842\,
            I => \b2v_inst6.countZ0Z_14\
        );

    \I__8015\ : InMux
    port map (
            O => \N__34837\,
            I => \N__34831\
        );

    \I__8014\ : InMux
    port map (
            O => \N__34836\,
            I => \N__34831\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__34831\,
            I => \b2v_inst6.count_rst_13\
        );

    \I__8012\ : InMux
    port map (
            O => \N__34828\,
            I => \N__34825\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__34825\,
            I => \b2v_inst6.count_3_14\
        );

    \I__8010\ : InMux
    port map (
            O => \N__34822\,
            I => \N__34819\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__34819\,
            I => \b2v_inst6.count_3_15\
        );

    \I__8008\ : InMux
    port map (
            O => \N__34816\,
            I => \N__34812\
        );

    \I__8007\ : InMux
    port map (
            O => \N__34815\,
            I => \N__34809\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__34812\,
            I => \b2v_inst6.count_rst_14\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__34809\,
            I => \b2v_inst6.count_rst_14\
        );

    \I__8004\ : CascadeMux
    port map (
            O => \N__34804\,
            I => \N__34800\
        );

    \I__8003\ : InMux
    port map (
            O => \N__34803\,
            I => \N__34797\
        );

    \I__8002\ : InMux
    port map (
            O => \N__34800\,
            I => \N__34794\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__34797\,
            I => \b2v_inst6.countZ0Z_15\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__34794\,
            I => \b2v_inst6.countZ0Z_15\
        );

    \I__7999\ : InMux
    port map (
            O => \N__34789\,
            I => \N__34786\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__34786\,
            I => \V5A_OK_c\
        );

    \I__7997\ : InMux
    port map (
            O => \N__34783\,
            I => \N__34780\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__34780\,
            I => \V33A_OK_c\
        );

    \I__7995\ : CascadeMux
    port map (
            O => \N__34777\,
            I => \N__34774\
        );

    \I__7994\ : InMux
    port map (
            O => \N__34774\,
            I => \N__34771\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__34771\,
            I => \V1P8A_OK_c\
        );

    \I__7992\ : InMux
    port map (
            O => \N__34768\,
            I => \N__34765\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__34765\,
            I => \N__34762\
        );

    \I__7990\ : IoSpan4Mux
    port map (
            O => \N__34762\,
            I => \N__34759\
        );

    \I__7989\ : Odrv4
    port map (
            O => \N__34759\,
            I => \V105A_OK_c\
        );

    \I__7988\ : InMux
    port map (
            O => \N__34756\,
            I => \N__34744\
        );

    \I__7987\ : InMux
    port map (
            O => \N__34755\,
            I => \N__34744\
        );

    \I__7986\ : InMux
    port map (
            O => \N__34754\,
            I => \N__34744\
        );

    \I__7985\ : InMux
    port map (
            O => \N__34753\,
            I => \N__34744\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__34744\,
            I => \N__34740\
        );

    \I__7983\ : InMux
    port map (
            O => \N__34743\,
            I => \N__34737\
        );

    \I__7982\ : Span12Mux_v
    port map (
            O => \N__34740\,
            I => \N__34732\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__34737\,
            I => \N__34732\
        );

    \I__7980\ : Odrv12
    port map (
            O => \N__34732\,
            I => \SYNTHESIZED_WIRE_26\
        );

    \I__7979\ : CascadeMux
    port map (
            O => \N__34729\,
            I => \b2v_inst6.count_rst_cascade_\
        );

    \I__7978\ : CascadeMux
    port map (
            O => \N__34726\,
            I => \b2v_inst6.countZ0Z_0_cascade_\
        );

    \I__7977\ : InMux
    port map (
            O => \N__34723\,
            I => \N__34720\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__34720\,
            I => \b2v_inst6.count_3_0\
        );

    \I__7975\ : InMux
    port map (
            O => \N__34717\,
            I => \N__34713\
        );

    \I__7974\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34710\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__34713\,
            I => \N__34707\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__34710\,
            I => \N__34704\
        );

    \I__7971\ : Odrv4
    port map (
            O => \N__34707\,
            I => \b2v_inst6.un2_count_1_cry_2_THRU_CO\
        );

    \I__7970\ : Odrv4
    port map (
            O => \N__34704\,
            I => \b2v_inst6.un2_count_1_cry_2_THRU_CO\
        );

    \I__7969\ : InMux
    port map (
            O => \N__34699\,
            I => \N__34696\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__34696\,
            I => \N__34693\
        );

    \I__7967\ : Odrv4
    port map (
            O => \N__34693\,
            I => \b2v_inst6.count_3_3\
        );

    \I__7966\ : ClkMux
    port map (
            O => \N__34690\,
            I => \N__34441\
        );

    \I__7965\ : ClkMux
    port map (
            O => \N__34689\,
            I => \N__34441\
        );

    \I__7964\ : ClkMux
    port map (
            O => \N__34688\,
            I => \N__34441\
        );

    \I__7963\ : ClkMux
    port map (
            O => \N__34687\,
            I => \N__34441\
        );

    \I__7962\ : ClkMux
    port map (
            O => \N__34686\,
            I => \N__34441\
        );

    \I__7961\ : ClkMux
    port map (
            O => \N__34685\,
            I => \N__34441\
        );

    \I__7960\ : ClkMux
    port map (
            O => \N__34684\,
            I => \N__34441\
        );

    \I__7959\ : ClkMux
    port map (
            O => \N__34683\,
            I => \N__34441\
        );

    \I__7958\ : ClkMux
    port map (
            O => \N__34682\,
            I => \N__34441\
        );

    \I__7957\ : ClkMux
    port map (
            O => \N__34681\,
            I => \N__34441\
        );

    \I__7956\ : ClkMux
    port map (
            O => \N__34680\,
            I => \N__34441\
        );

    \I__7955\ : ClkMux
    port map (
            O => \N__34679\,
            I => \N__34441\
        );

    \I__7954\ : ClkMux
    port map (
            O => \N__34678\,
            I => \N__34441\
        );

    \I__7953\ : ClkMux
    port map (
            O => \N__34677\,
            I => \N__34441\
        );

    \I__7952\ : ClkMux
    port map (
            O => \N__34676\,
            I => \N__34441\
        );

    \I__7951\ : ClkMux
    port map (
            O => \N__34675\,
            I => \N__34441\
        );

    \I__7950\ : ClkMux
    port map (
            O => \N__34674\,
            I => \N__34441\
        );

    \I__7949\ : ClkMux
    port map (
            O => \N__34673\,
            I => \N__34441\
        );

    \I__7948\ : ClkMux
    port map (
            O => \N__34672\,
            I => \N__34441\
        );

    \I__7947\ : ClkMux
    port map (
            O => \N__34671\,
            I => \N__34441\
        );

    \I__7946\ : ClkMux
    port map (
            O => \N__34670\,
            I => \N__34441\
        );

    \I__7945\ : ClkMux
    port map (
            O => \N__34669\,
            I => \N__34441\
        );

    \I__7944\ : ClkMux
    port map (
            O => \N__34668\,
            I => \N__34441\
        );

    \I__7943\ : ClkMux
    port map (
            O => \N__34667\,
            I => \N__34441\
        );

    \I__7942\ : ClkMux
    port map (
            O => \N__34666\,
            I => \N__34441\
        );

    \I__7941\ : ClkMux
    port map (
            O => \N__34665\,
            I => \N__34441\
        );

    \I__7940\ : ClkMux
    port map (
            O => \N__34664\,
            I => \N__34441\
        );

    \I__7939\ : ClkMux
    port map (
            O => \N__34663\,
            I => \N__34441\
        );

    \I__7938\ : ClkMux
    port map (
            O => \N__34662\,
            I => \N__34441\
        );

    \I__7937\ : ClkMux
    port map (
            O => \N__34661\,
            I => \N__34441\
        );

    \I__7936\ : ClkMux
    port map (
            O => \N__34660\,
            I => \N__34441\
        );

    \I__7935\ : ClkMux
    port map (
            O => \N__34659\,
            I => \N__34441\
        );

    \I__7934\ : ClkMux
    port map (
            O => \N__34658\,
            I => \N__34441\
        );

    \I__7933\ : ClkMux
    port map (
            O => \N__34657\,
            I => \N__34441\
        );

    \I__7932\ : ClkMux
    port map (
            O => \N__34656\,
            I => \N__34441\
        );

    \I__7931\ : ClkMux
    port map (
            O => \N__34655\,
            I => \N__34441\
        );

    \I__7930\ : ClkMux
    port map (
            O => \N__34654\,
            I => \N__34441\
        );

    \I__7929\ : ClkMux
    port map (
            O => \N__34653\,
            I => \N__34441\
        );

    \I__7928\ : ClkMux
    port map (
            O => \N__34652\,
            I => \N__34441\
        );

    \I__7927\ : ClkMux
    port map (
            O => \N__34651\,
            I => \N__34441\
        );

    \I__7926\ : ClkMux
    port map (
            O => \N__34650\,
            I => \N__34441\
        );

    \I__7925\ : ClkMux
    port map (
            O => \N__34649\,
            I => \N__34441\
        );

    \I__7924\ : ClkMux
    port map (
            O => \N__34648\,
            I => \N__34441\
        );

    \I__7923\ : ClkMux
    port map (
            O => \N__34647\,
            I => \N__34441\
        );

    \I__7922\ : ClkMux
    port map (
            O => \N__34646\,
            I => \N__34441\
        );

    \I__7921\ : ClkMux
    port map (
            O => \N__34645\,
            I => \N__34441\
        );

    \I__7920\ : ClkMux
    port map (
            O => \N__34644\,
            I => \N__34441\
        );

    \I__7919\ : ClkMux
    port map (
            O => \N__34643\,
            I => \N__34441\
        );

    \I__7918\ : ClkMux
    port map (
            O => \N__34642\,
            I => \N__34441\
        );

    \I__7917\ : ClkMux
    port map (
            O => \N__34641\,
            I => \N__34441\
        );

    \I__7916\ : ClkMux
    port map (
            O => \N__34640\,
            I => \N__34441\
        );

    \I__7915\ : ClkMux
    port map (
            O => \N__34639\,
            I => \N__34441\
        );

    \I__7914\ : ClkMux
    port map (
            O => \N__34638\,
            I => \N__34441\
        );

    \I__7913\ : ClkMux
    port map (
            O => \N__34637\,
            I => \N__34441\
        );

    \I__7912\ : ClkMux
    port map (
            O => \N__34636\,
            I => \N__34441\
        );

    \I__7911\ : ClkMux
    port map (
            O => \N__34635\,
            I => \N__34441\
        );

    \I__7910\ : ClkMux
    port map (
            O => \N__34634\,
            I => \N__34441\
        );

    \I__7909\ : ClkMux
    port map (
            O => \N__34633\,
            I => \N__34441\
        );

    \I__7908\ : ClkMux
    port map (
            O => \N__34632\,
            I => \N__34441\
        );

    \I__7907\ : ClkMux
    port map (
            O => \N__34631\,
            I => \N__34441\
        );

    \I__7906\ : ClkMux
    port map (
            O => \N__34630\,
            I => \N__34441\
        );

    \I__7905\ : ClkMux
    port map (
            O => \N__34629\,
            I => \N__34441\
        );

    \I__7904\ : ClkMux
    port map (
            O => \N__34628\,
            I => \N__34441\
        );

    \I__7903\ : ClkMux
    port map (
            O => \N__34627\,
            I => \N__34441\
        );

    \I__7902\ : ClkMux
    port map (
            O => \N__34626\,
            I => \N__34441\
        );

    \I__7901\ : ClkMux
    port map (
            O => \N__34625\,
            I => \N__34441\
        );

    \I__7900\ : ClkMux
    port map (
            O => \N__34624\,
            I => \N__34441\
        );

    \I__7899\ : ClkMux
    port map (
            O => \N__34623\,
            I => \N__34441\
        );

    \I__7898\ : ClkMux
    port map (
            O => \N__34622\,
            I => \N__34441\
        );

    \I__7897\ : ClkMux
    port map (
            O => \N__34621\,
            I => \N__34441\
        );

    \I__7896\ : ClkMux
    port map (
            O => \N__34620\,
            I => \N__34441\
        );

    \I__7895\ : ClkMux
    port map (
            O => \N__34619\,
            I => \N__34441\
        );

    \I__7894\ : ClkMux
    port map (
            O => \N__34618\,
            I => \N__34441\
        );

    \I__7893\ : ClkMux
    port map (
            O => \N__34617\,
            I => \N__34441\
        );

    \I__7892\ : ClkMux
    port map (
            O => \N__34616\,
            I => \N__34441\
        );

    \I__7891\ : ClkMux
    port map (
            O => \N__34615\,
            I => \N__34441\
        );

    \I__7890\ : ClkMux
    port map (
            O => \N__34614\,
            I => \N__34441\
        );

    \I__7889\ : ClkMux
    port map (
            O => \N__34613\,
            I => \N__34441\
        );

    \I__7888\ : ClkMux
    port map (
            O => \N__34612\,
            I => \N__34441\
        );

    \I__7887\ : ClkMux
    port map (
            O => \N__34611\,
            I => \N__34441\
        );

    \I__7886\ : ClkMux
    port map (
            O => \N__34610\,
            I => \N__34441\
        );

    \I__7885\ : ClkMux
    port map (
            O => \N__34609\,
            I => \N__34441\
        );

    \I__7884\ : ClkMux
    port map (
            O => \N__34608\,
            I => \N__34441\
        );

    \I__7883\ : GlobalMux
    port map (
            O => \N__34441\,
            I => \N__34438\
        );

    \I__7882\ : gio2CtrlBuf
    port map (
            O => \N__34438\,
            I => \FPGA_OSC_0_c_g\
        );

    \I__7881\ : CEMux
    port map (
            O => \N__34435\,
            I => \N__34431\
        );

    \I__7880\ : CEMux
    port map (
            O => \N__34434\,
            I => \N__34422\
        );

    \I__7879\ : LocalMux
    port map (
            O => \N__34431\,
            I => \N__34411\
        );

    \I__7878\ : CEMux
    port map (
            O => \N__34430\,
            I => \N__34408\
        );

    \I__7877\ : CEMux
    port map (
            O => \N__34429\,
            I => \N__34405\
        );

    \I__7876\ : InMux
    port map (
            O => \N__34428\,
            I => \N__34396\
        );

    \I__7875\ : InMux
    port map (
            O => \N__34427\,
            I => \N__34396\
        );

    \I__7874\ : InMux
    port map (
            O => \N__34426\,
            I => \N__34396\
        );

    \I__7873\ : InMux
    port map (
            O => \N__34425\,
            I => \N__34396\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__34422\,
            I => \N__34393\
        );

    \I__7871\ : CEMux
    port map (
            O => \N__34421\,
            I => \N__34390\
        );

    \I__7870\ : CEMux
    port map (
            O => \N__34420\,
            I => \N__34387\
        );

    \I__7869\ : InMux
    port map (
            O => \N__34419\,
            I => \N__34382\
        );

    \I__7868\ : InMux
    port map (
            O => \N__34418\,
            I => \N__34382\
        );

    \I__7867\ : CEMux
    port map (
            O => \N__34417\,
            I => \N__34373\
        );

    \I__7866\ : InMux
    port map (
            O => \N__34416\,
            I => \N__34373\
        );

    \I__7865\ : InMux
    port map (
            O => \N__34415\,
            I => \N__34373\
        );

    \I__7864\ : InMux
    port map (
            O => \N__34414\,
            I => \N__34373\
        );

    \I__7863\ : Span4Mux_s3_h
    port map (
            O => \N__34411\,
            I => \N__34365\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__34408\,
            I => \N__34358\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__34405\,
            I => \N__34358\
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__34396\,
            I => \N__34358\
        );

    \I__7859\ : Span4Mux_s1_v
    port map (
            O => \N__34393\,
            I => \N__34353\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__34390\,
            I => \N__34353\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__34387\,
            I => \N__34350\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__34382\,
            I => \N__34347\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__34373\,
            I => \N__34342\
        );

    \I__7854\ : InMux
    port map (
            O => \N__34372\,
            I => \N__34333\
        );

    \I__7853\ : InMux
    port map (
            O => \N__34371\,
            I => \N__34333\
        );

    \I__7852\ : InMux
    port map (
            O => \N__34370\,
            I => \N__34333\
        );

    \I__7851\ : InMux
    port map (
            O => \N__34369\,
            I => \N__34333\
        );

    \I__7850\ : InMux
    port map (
            O => \N__34368\,
            I => \N__34330\
        );

    \I__7849\ : Span4Mux_h
    port map (
            O => \N__34365\,
            I => \N__34325\
        );

    \I__7848\ : Span4Mux_s3_h
    port map (
            O => \N__34358\,
            I => \N__34325\
        );

    \I__7847\ : Span4Mux_s1_h
    port map (
            O => \N__34353\,
            I => \N__34318\
        );

    \I__7846\ : Span4Mux_s1_h
    port map (
            O => \N__34350\,
            I => \N__34318\
        );

    \I__7845\ : Span4Mux_s1_v
    port map (
            O => \N__34347\,
            I => \N__34318\
        );

    \I__7844\ : InMux
    port map (
            O => \N__34346\,
            I => \N__34313\
        );

    \I__7843\ : InMux
    port map (
            O => \N__34345\,
            I => \N__34313\
        );

    \I__7842\ : Span4Mux_s3_h
    port map (
            O => \N__34342\,
            I => \N__34310\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__34333\,
            I => \N__34305\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__34330\,
            I => \N__34305\
        );

    \I__7839\ : Odrv4
    port map (
            O => \N__34325\,
            I => \b2v_inst6.count_en\
        );

    \I__7838\ : Odrv4
    port map (
            O => \N__34318\,
            I => \b2v_inst6.count_en\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__34313\,
            I => \b2v_inst6.count_en\
        );

    \I__7836\ : Odrv4
    port map (
            O => \N__34310\,
            I => \b2v_inst6.count_en\
        );

    \I__7835\ : Odrv12
    port map (
            O => \N__34305\,
            I => \b2v_inst6.count_en\
        );

    \I__7834\ : CascadeMux
    port map (
            O => \N__34294\,
            I => \b2v_inst6.countZ0Z_1_cascade_\
        );

    \I__7833\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34288\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__34288\,
            I => \b2v_inst6.count_3_1\
        );

    \I__7831\ : InMux
    port map (
            O => \N__34285\,
            I => \N__34279\
        );

    \I__7830\ : InMux
    port map (
            O => \N__34284\,
            I => \N__34279\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__34279\,
            I => \b2v_inst6.count_rst_1\
        );

    \I__7828\ : InMux
    port map (
            O => \N__34276\,
            I => \N__34273\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__34273\,
            I => \b2v_inst6.count_3_2\
        );

    \I__7826\ : InMux
    port map (
            O => \N__34270\,
            I => \N__34267\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__34267\,
            I => \b2v_inst6.count_3_6\
        );

    \I__7824\ : InMux
    port map (
            O => \N__34264\,
            I => \N__34258\
        );

    \I__7823\ : InMux
    port map (
            O => \N__34263\,
            I => \N__34258\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__34258\,
            I => \b2v_inst6.count_rst_5\
        );

    \I__7821\ : InMux
    port map (
            O => \N__34255\,
            I => \N__34252\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__34252\,
            I => \b2v_inst6.countZ0Z_6\
        );

    \I__7819\ : InMux
    port map (
            O => \N__34249\,
            I => \N__34246\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__34246\,
            I => \N__34243\
        );

    \I__7817\ : Span4Mux_s0_h
    port map (
            O => \N__34243\,
            I => \N__34239\
        );

    \I__7816\ : InMux
    port map (
            O => \N__34242\,
            I => \N__34236\
        );

    \I__7815\ : Odrv4
    port map (
            O => \N__34239\,
            I => \b2v_inst6.countZ0Z_10\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__34236\,
            I => \b2v_inst6.countZ0Z_10\
        );

    \I__7813\ : InMux
    port map (
            O => \N__34231\,
            I => \N__34227\
        );

    \I__7812\ : InMux
    port map (
            O => \N__34230\,
            I => \N__34224\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__34227\,
            I => \b2v_inst6.countZ0Z_2\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__34224\,
            I => \b2v_inst6.countZ0Z_2\
        );

    \I__7809\ : CascadeMux
    port map (
            O => \N__34219\,
            I => \b2v_inst6.countZ0Z_6_cascade_\
        );

    \I__7808\ : InMux
    port map (
            O => \N__34216\,
            I => \N__34209\
        );

    \I__7807\ : InMux
    port map (
            O => \N__34215\,
            I => \N__34209\
        );

    \I__7806\ : InMux
    port map (
            O => \N__34214\,
            I => \N__34206\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__34209\,
            I => \b2v_inst6.countZ0Z_1\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__34206\,
            I => \b2v_inst6.countZ0Z_1\
        );

    \I__7803\ : InMux
    port map (
            O => \N__34201\,
            I => \N__34197\
        );

    \I__7802\ : InMux
    port map (
            O => \N__34200\,
            I => \N__34194\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__34197\,
            I => \b2v_inst6.countZ0Z_12\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__34194\,
            I => \b2v_inst6.countZ0Z_12\
        );

    \I__7799\ : InMux
    port map (
            O => \N__34189\,
            I => \N__34183\
        );

    \I__7798\ : InMux
    port map (
            O => \N__34188\,
            I => \N__34183\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__34183\,
            I => \b2v_inst6.count_rst_11\
        );

    \I__7796\ : InMux
    port map (
            O => \N__34180\,
            I => \N__34177\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__34177\,
            I => \b2v_inst6.count_3_12\
        );

    \I__7794\ : InMux
    port map (
            O => \N__34174\,
            I => \N__34170\
        );

    \I__7793\ : InMux
    port map (
            O => \N__34173\,
            I => \N__34167\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__34170\,
            I => \b2v_inst6.countZ0Z_13\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__34167\,
            I => \b2v_inst6.countZ0Z_13\
        );

    \I__7790\ : InMux
    port map (
            O => \N__34162\,
            I => \N__34156\
        );

    \I__7789\ : InMux
    port map (
            O => \N__34161\,
            I => \N__34156\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__34156\,
            I => \b2v_inst6.count_rst_12\
        );

    \I__7787\ : InMux
    port map (
            O => \N__34153\,
            I => \N__34150\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__34150\,
            I => \b2v_inst6.count_3_13\
        );

    \I__7785\ : InMux
    port map (
            O => \N__34147\,
            I => \N__34142\
        );

    \I__7784\ : InMux
    port map (
            O => \N__34146\,
            I => \N__34139\
        );

    \I__7783\ : InMux
    port map (
            O => \N__34145\,
            I => \N__34136\
        );

    \I__7782\ : LocalMux
    port map (
            O => \N__34142\,
            I => \N__34129\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__34139\,
            I => \N__34129\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__34136\,
            I => \N__34129\
        );

    \I__7779\ : Span12Mux_s9_v
    port map (
            O => \N__34129\,
            I => \N__34126\
        );

    \I__7778\ : Odrv12
    port map (
            O => \N__34126\,
            I => \b2v_inst200.m11_0_a3_0\
        );

    \I__7777\ : CascadeMux
    port map (
            O => \N__34123\,
            I => \N__34120\
        );

    \I__7776\ : InMux
    port map (
            O => \N__34120\,
            I => \N__34117\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__34117\,
            I => \b2v_inst200.N_202\
        );

    \I__7774\ : InMux
    port map (
            O => \N__34114\,
            I => \N__34111\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__34111\,
            I => \N__34108\
        );

    \I__7772\ : Odrv4
    port map (
            O => \N__34108\,
            I => \G_2788\
        );

    \I__7771\ : InMux
    port map (
            O => \N__34105\,
            I => \N__34102\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__34102\,
            I => \N__34099\
        );

    \I__7769\ : Odrv4
    port map (
            O => \N__34099\,
            I => \b2v_inst200.curr_state_0_2\
        );

    \I__7768\ : CascadeMux
    port map (
            O => \N__34096\,
            I => \G_2788_cascade_\
        );

    \I__7767\ : InMux
    port map (
            O => \N__34093\,
            I => \N__34080\
        );

    \I__7766\ : InMux
    port map (
            O => \N__34092\,
            I => \N__34080\
        );

    \I__7765\ : CascadeMux
    port map (
            O => \N__34091\,
            I => \N__34066\
        );

    \I__7764\ : InMux
    port map (
            O => \N__34090\,
            I => \N__34061\
        );

    \I__7763\ : InMux
    port map (
            O => \N__34089\,
            I => \N__34041\
        );

    \I__7762\ : InMux
    port map (
            O => \N__34088\,
            I => \N__34041\
        );

    \I__7761\ : InMux
    port map (
            O => \N__34087\,
            I => \N__34041\
        );

    \I__7760\ : InMux
    port map (
            O => \N__34086\,
            I => \N__34041\
        );

    \I__7759\ : CascadeMux
    port map (
            O => \N__34085\,
            I => \N__34038\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__34080\,
            I => \N__34033\
        );

    \I__7757\ : InMux
    port map (
            O => \N__34079\,
            I => \N__34024\
        );

    \I__7756\ : InMux
    port map (
            O => \N__34078\,
            I => \N__34024\
        );

    \I__7755\ : InMux
    port map (
            O => \N__34077\,
            I => \N__34024\
        );

    \I__7754\ : InMux
    port map (
            O => \N__34076\,
            I => \N__34024\
        );

    \I__7753\ : InMux
    port map (
            O => \N__34075\,
            I => \N__34017\
        );

    \I__7752\ : InMux
    port map (
            O => \N__34074\,
            I => \N__34017\
        );

    \I__7751\ : InMux
    port map (
            O => \N__34073\,
            I => \N__34017\
        );

    \I__7750\ : InMux
    port map (
            O => \N__34072\,
            I => \N__34012\
        );

    \I__7749\ : InMux
    port map (
            O => \N__34071\,
            I => \N__34012\
        );

    \I__7748\ : InMux
    port map (
            O => \N__34070\,
            I => \N__34007\
        );

    \I__7747\ : InMux
    port map (
            O => \N__34069\,
            I => \N__34007\
        );

    \I__7746\ : InMux
    port map (
            O => \N__34066\,
            I => \N__34003\
        );

    \I__7745\ : InMux
    port map (
            O => \N__34065\,
            I => \N__33998\
        );

    \I__7744\ : InMux
    port map (
            O => \N__34064\,
            I => \N__33998\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__34061\,
            I => \N__33995\
        );

    \I__7742\ : InMux
    port map (
            O => \N__34060\,
            I => \N__33991\
        );

    \I__7741\ : InMux
    port map (
            O => \N__34059\,
            I => \N__33986\
        );

    \I__7740\ : InMux
    port map (
            O => \N__34058\,
            I => \N__33986\
        );

    \I__7739\ : InMux
    port map (
            O => \N__34057\,
            I => \N__33983\
        );

    \I__7738\ : InMux
    port map (
            O => \N__34056\,
            I => \N__33974\
        );

    \I__7737\ : InMux
    port map (
            O => \N__34055\,
            I => \N__33974\
        );

    \I__7736\ : InMux
    port map (
            O => \N__34054\,
            I => \N__33974\
        );

    \I__7735\ : InMux
    port map (
            O => \N__34053\,
            I => \N__33974\
        );

    \I__7734\ : InMux
    port map (
            O => \N__34052\,
            I => \N__33967\
        );

    \I__7733\ : InMux
    port map (
            O => \N__34051\,
            I => \N__33967\
        );

    \I__7732\ : InMux
    port map (
            O => \N__34050\,
            I => \N__33967\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__34041\,
            I => \N__33964\
        );

    \I__7730\ : InMux
    port map (
            O => \N__34038\,
            I => \N__33957\
        );

    \I__7729\ : InMux
    port map (
            O => \N__34037\,
            I => \N__33957\
        );

    \I__7728\ : InMux
    port map (
            O => \N__34036\,
            I => \N__33957\
        );

    \I__7727\ : Span4Mux_h
    port map (
            O => \N__34033\,
            I => \N__33952\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__34024\,
            I => \N__33952\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__34017\,
            I => \N__33949\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__34012\,
            I => \N__33946\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__34007\,
            I => \N__33943\
        );

    \I__7722\ : InMux
    port map (
            O => \N__34006\,
            I => \N__33940\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__34003\,
            I => \N__33933\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__33998\,
            I => \N__33933\
        );

    \I__7719\ : Span4Mux_h
    port map (
            O => \N__33995\,
            I => \N__33933\
        );

    \I__7718\ : InMux
    port map (
            O => \N__33994\,
            I => \N__33930\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__33991\,
            I => \N__33924\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__33986\,
            I => \N__33924\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__33983\,
            I => \N__33919\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__33974\,
            I => \N__33919\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__33967\,
            I => \N__33912\
        );

    \I__7712\ : Span4Mux_h
    port map (
            O => \N__33964\,
            I => \N__33912\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__33957\,
            I => \N__33912\
        );

    \I__7710\ : Sp12to4
    port map (
            O => \N__33952\,
            I => \N__33907\
        );

    \I__7709\ : Span12Mux_s2_h
    port map (
            O => \N__33949\,
            I => \N__33907\
        );

    \I__7708\ : Span4Mux_s0_h
    port map (
            O => \N__33946\,
            I => \N__33899\
        );

    \I__7707\ : Span4Mux_v
    port map (
            O => \N__33943\,
            I => \N__33899\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__33940\,
            I => \N__33896\
        );

    \I__7705\ : Span4Mux_v
    port map (
            O => \N__33933\,
            I => \N__33891\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__33930\,
            I => \N__33891\
        );

    \I__7703\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33888\
        );

    \I__7702\ : Span12Mux_v
    port map (
            O => \N__33924\,
            I => \N__33885\
        );

    \I__7701\ : Span12Mux_s8_v
    port map (
            O => \N__33919\,
            I => \N__33880\
        );

    \I__7700\ : Sp12to4
    port map (
            O => \N__33912\,
            I => \N__33880\
        );

    \I__7699\ : Span12Mux_v
    port map (
            O => \N__33907\,
            I => \N__33877\
        );

    \I__7698\ : InMux
    port map (
            O => \N__33906\,
            I => \N__33870\
        );

    \I__7697\ : InMux
    port map (
            O => \N__33905\,
            I => \N__33870\
        );

    \I__7696\ : InMux
    port map (
            O => \N__33904\,
            I => \N__33870\
        );

    \I__7695\ : Span4Mux_h
    port map (
            O => \N__33899\,
            I => \N__33863\
        );

    \I__7694\ : Span4Mux_h
    port map (
            O => \N__33896\,
            I => \N__33863\
        );

    \I__7693\ : Span4Mux_h
    port map (
            O => \N__33891\,
            I => \N__33863\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__33888\,
            I => \SYNTHESIZED_WIRE_47keep\
        );

    \I__7691\ : Odrv12
    port map (
            O => \N__33885\,
            I => \SYNTHESIZED_WIRE_47keep\
        );

    \I__7690\ : Odrv12
    port map (
            O => \N__33880\,
            I => \SYNTHESIZED_WIRE_47keep\
        );

    \I__7689\ : Odrv12
    port map (
            O => \N__33877\,
            I => \SYNTHESIZED_WIRE_47keep\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__33870\,
            I => \SYNTHESIZED_WIRE_47keep\
        );

    \I__7687\ : Odrv4
    port map (
            O => \N__33863\,
            I => \SYNTHESIZED_WIRE_47keep\
        );

    \I__7686\ : InMux
    port map (
            O => \N__33850\,
            I => \N__33844\
        );

    \I__7685\ : InMux
    port map (
            O => \N__33849\,
            I => \N__33844\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__33844\,
            I => \b2v_inst200.curr_stateZ0Z_2\
        );

    \I__7683\ : CascadeMux
    port map (
            O => \N__33841\,
            I => \b2v_inst200.curr_stateZ0Z_2_cascade_\
        );

    \I__7682\ : InMux
    port map (
            O => \N__33838\,
            I => \N__33835\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__33835\,
            I => \b2v_inst200.HDA_SDO_FPGA_0\
        );

    \I__7680\ : InMux
    port map (
            O => \N__33832\,
            I => \N__33823\
        );

    \I__7679\ : InMux
    port map (
            O => \N__33831\,
            I => \N__33823\
        );

    \I__7678\ : InMux
    port map (
            O => \N__33830\,
            I => \N__33823\
        );

    \I__7677\ : LocalMux
    port map (
            O => \N__33823\,
            I => \N__33818\
        );

    \I__7676\ : InMux
    port map (
            O => \N__33822\,
            I => \N__33813\
        );

    \I__7675\ : InMux
    port map (
            O => \N__33821\,
            I => \N__33813\
        );

    \I__7674\ : Odrv4
    port map (
            O => \N__33818\,
            I => \b2v_inst200.curr_stateZ0Z_0\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__33813\,
            I => \b2v_inst200.curr_stateZ0Z_0\
        );

    \I__7672\ : InMux
    port map (
            O => \N__33808\,
            I => \N__33797\
        );

    \I__7671\ : InMux
    port map (
            O => \N__33807\,
            I => \N__33797\
        );

    \I__7670\ : InMux
    port map (
            O => \N__33806\,
            I => \N__33794\
        );

    \I__7669\ : InMux
    port map (
            O => \N__33805\,
            I => \N__33785\
        );

    \I__7668\ : InMux
    port map (
            O => \N__33804\,
            I => \N__33785\
        );

    \I__7667\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33785\
        );

    \I__7666\ : InMux
    port map (
            O => \N__33802\,
            I => \N__33785\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__33797\,
            I => \b2v_inst200.curr_stateZ0Z_1\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__33794\,
            I => \b2v_inst200.curr_stateZ0Z_1\
        );

    \I__7663\ : LocalMux
    port map (
            O => \N__33785\,
            I => \b2v_inst200.curr_stateZ0Z_1\
        );

    \I__7662\ : InMux
    port map (
            O => \N__33778\,
            I => \N__33774\
        );

    \I__7661\ : CascadeMux
    port map (
            O => \N__33777\,
            I => \N__33771\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__33774\,
            I => \N__33764\
        );

    \I__7659\ : InMux
    port map (
            O => \N__33771\,
            I => \N__33759\
        );

    \I__7658\ : InMux
    port map (
            O => \N__33770\,
            I => \N__33759\
        );

    \I__7657\ : InMux
    port map (
            O => \N__33769\,
            I => \N__33752\
        );

    \I__7656\ : InMux
    port map (
            O => \N__33768\,
            I => \N__33752\
        );

    \I__7655\ : InMux
    port map (
            O => \N__33767\,
            I => \N__33752\
        );

    \I__7654\ : Span4Mux_h
    port map (
            O => \N__33764\,
            I => \N__33749\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__33759\,
            I => \N__33746\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__33752\,
            I => \N__33743\
        );

    \I__7651\ : Span4Mux_h
    port map (
            O => \N__33749\,
            I => \N__33738\
        );

    \I__7650\ : Span4Mux_s2_h
    port map (
            O => \N__33746\,
            I => \N__33738\
        );

    \I__7649\ : Span4Mux_s2_h
    port map (
            O => \N__33743\,
            I => \N__33735\
        );

    \I__7648\ : Odrv4
    port map (
            O => \N__33738\,
            I => \N_219\
        );

    \I__7647\ : Odrv4
    port map (
            O => \N__33735\,
            I => \N_219\
        );

    \I__7646\ : InMux
    port map (
            O => \N__33730\,
            I => \N__33727\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__33727\,
            I => \b2v_inst200.m6_i_0\
        );

    \I__7644\ : InMux
    port map (
            O => \N__33724\,
            I => \N__33721\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__33721\,
            I => \b2v_inst200.curr_state_0_0\
        );

    \I__7642\ : InMux
    port map (
            O => \N__33718\,
            I => \N__33709\
        );

    \I__7641\ : InMux
    port map (
            O => \N__33717\,
            I => \N__33706\
        );

    \I__7640\ : InMux
    port map (
            O => \N__33716\,
            I => \N__33703\
        );

    \I__7639\ : InMux
    port map (
            O => \N__33715\,
            I => \N__33698\
        );

    \I__7638\ : InMux
    port map (
            O => \N__33714\,
            I => \N__33698\
        );

    \I__7637\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33693\
        );

    \I__7636\ : InMux
    port map (
            O => \N__33712\,
            I => \N__33693\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__33709\,
            I => \N__33690\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__33706\,
            I => \N__33675\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__33703\,
            I => \N__33672\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__33698\,
            I => \N__33669\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__33693\,
            I => \N__33666\
        );

    \I__7630\ : Glb2LocalMux
    port map (
            O => \N__33690\,
            I => \N__33631\
        );

    \I__7629\ : CEMux
    port map (
            O => \N__33689\,
            I => \N__33631\
        );

    \I__7628\ : CEMux
    port map (
            O => \N__33688\,
            I => \N__33631\
        );

    \I__7627\ : CEMux
    port map (
            O => \N__33687\,
            I => \N__33631\
        );

    \I__7626\ : CEMux
    port map (
            O => \N__33686\,
            I => \N__33631\
        );

    \I__7625\ : CEMux
    port map (
            O => \N__33685\,
            I => \N__33631\
        );

    \I__7624\ : CEMux
    port map (
            O => \N__33684\,
            I => \N__33631\
        );

    \I__7623\ : CEMux
    port map (
            O => \N__33683\,
            I => \N__33631\
        );

    \I__7622\ : CEMux
    port map (
            O => \N__33682\,
            I => \N__33631\
        );

    \I__7621\ : CEMux
    port map (
            O => \N__33681\,
            I => \N__33631\
        );

    \I__7620\ : CEMux
    port map (
            O => \N__33680\,
            I => \N__33631\
        );

    \I__7619\ : CEMux
    port map (
            O => \N__33679\,
            I => \N__33631\
        );

    \I__7618\ : CEMux
    port map (
            O => \N__33678\,
            I => \N__33631\
        );

    \I__7617\ : Glb2LocalMux
    port map (
            O => \N__33675\,
            I => \N__33631\
        );

    \I__7616\ : Glb2LocalMux
    port map (
            O => \N__33672\,
            I => \N__33631\
        );

    \I__7615\ : Glb2LocalMux
    port map (
            O => \N__33669\,
            I => \N__33631\
        );

    \I__7614\ : Glb2LocalMux
    port map (
            O => \N__33666\,
            I => \N__33631\
        );

    \I__7613\ : GlobalMux
    port map (
            O => \N__33631\,
            I => \N__33628\
        );

    \I__7612\ : gio2CtrlBuf
    port map (
            O => \N__33628\,
            I => b2v_inst16_delayed_vddq_pwrgd_en_g
        );

    \I__7611\ : CascadeMux
    port map (
            O => \N__33625\,
            I => \b2v_inst6.count_rst_0_cascade_\
        );

    \I__7610\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33619\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__33619\,
            I => \GPIO_FPGA_PCH_1_c\
        );

    \I__7608\ : InMux
    port map (
            O => \N__33616\,
            I => \N__33613\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__33613\,
            I => \N__33610\
        );

    \I__7606\ : Span4Mux_v
    port map (
            O => \N__33610\,
            I => \N__33605\
        );

    \I__7605\ : InMux
    port map (
            O => \N__33609\,
            I => \N__33599\
        );

    \I__7604\ : InMux
    port map (
            O => \N__33608\,
            I => \N__33599\
        );

    \I__7603\ : Sp12to4
    port map (
            O => \N__33605\,
            I => \N__33596\
        );

    \I__7602\ : CascadeMux
    port map (
            O => \N__33604\,
            I => \N__33587\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__33599\,
            I => \N__33582\
        );

    \I__7600\ : Span12Mux_s11_h
    port map (
            O => \N__33596\,
            I => \N__33579\
        );

    \I__7599\ : InMux
    port map (
            O => \N__33595\,
            I => \N__33570\
        );

    \I__7598\ : InMux
    port map (
            O => \N__33594\,
            I => \N__33570\
        );

    \I__7597\ : InMux
    port map (
            O => \N__33593\,
            I => \N__33570\
        );

    \I__7596\ : InMux
    port map (
            O => \N__33592\,
            I => \N__33570\
        );

    \I__7595\ : InMux
    port map (
            O => \N__33591\,
            I => \N__33561\
        );

    \I__7594\ : InMux
    port map (
            O => \N__33590\,
            I => \N__33561\
        );

    \I__7593\ : InMux
    port map (
            O => \N__33587\,
            I => \N__33561\
        );

    \I__7592\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33561\
        );

    \I__7591\ : InMux
    port map (
            O => \N__33585\,
            I => \N__33558\
        );

    \I__7590\ : Odrv4
    port map (
            O => \N__33582\,
            I => \b2v_inst200.count_RNI_0_0\
        );

    \I__7589\ : Odrv12
    port map (
            O => \N__33579\,
            I => \b2v_inst200.count_RNI_0_0\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__33570\,
            I => \b2v_inst200.count_RNI_0_0\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__33561\,
            I => \b2v_inst200.count_RNI_0_0\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__33558\,
            I => \b2v_inst200.count_RNI_0_0\
        );

    \I__7585\ : CascadeMux
    port map (
            O => \N__33547\,
            I => \N_405_cascade_\
        );

    \I__7584\ : CascadeMux
    port map (
            O => \N__33544\,
            I => \b2v_inst200.m6_i_0_cascade_\
        );

    \I__7583\ : CascadeMux
    port map (
            O => \N__33541\,
            I => \b2v_inst200.N_57_cascade_\
        );

    \I__7582\ : CascadeMux
    port map (
            O => \N__33538\,
            I => \b2v_inst200.curr_stateZ0Z_0_cascade_\
        );

    \I__7581\ : CascadeMux
    port map (
            O => \N__33535\,
            I => \N_406_cascade_\
        );

    \I__7580\ : InMux
    port map (
            O => \N__33532\,
            I => \N__33529\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__33529\,
            I => \b2v_inst200.N_55\
        );

    \I__7578\ : CascadeMux
    port map (
            O => \N__33526\,
            I => \N__33523\
        );

    \I__7577\ : InMux
    port map (
            O => \N__33523\,
            I => \N__33517\
        );

    \I__7576\ : InMux
    port map (
            O => \N__33522\,
            I => \N__33517\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__33517\,
            I => \N_406\
        );

    \I__7574\ : InMux
    port map (
            O => \N__33514\,
            I => \N__33511\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__33511\,
            I => \b2v_inst200.curr_state_0_1\
        );

    \I__7572\ : CascadeMux
    port map (
            O => \N__33508\,
            I => \b2v_inst200.N_202_cascade_\
        );

    \I__7571\ : IoInMux
    port map (
            O => \N__33505\,
            I => \N__33502\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__33502\,
            I => \N__33499\
        );

    \I__7569\ : IoSpan4Mux
    port map (
            O => \N__33499\,
            I => \N__33496\
        );

    \I__7568\ : Span4Mux_s3_h
    port map (
            O => \N__33496\,
            I => \N__33493\
        );

    \I__7567\ : Span4Mux_h
    port map (
            O => \N__33493\,
            I => \N__33490\
        );

    \I__7566\ : Span4Mux_h
    port map (
            O => \N__33490\,
            I => \N__33487\
        );

    \I__7565\ : Odrv4
    port map (
            O => \N__33487\,
            I => \HDA_SDO_FPGA_c\
        );

    \I__7564\ : InMux
    port map (
            O => \N__33484\,
            I => \N__33480\
        );

    \I__7563\ : InMux
    port map (
            O => \N__33483\,
            I => \N__33477\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__33480\,
            I => \b2v_inst20.counterZ0Z_29\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__33477\,
            I => \b2v_inst20.counterZ0Z_29\
        );

    \I__7560\ : InMux
    port map (
            O => \N__33472\,
            I => \N__33468\
        );

    \I__7559\ : InMux
    port map (
            O => \N__33471\,
            I => \N__33465\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__33468\,
            I => \b2v_inst20.counterZ0Z_28\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__33465\,
            I => \b2v_inst20.counterZ0Z_28\
        );

    \I__7556\ : CascadeMux
    port map (
            O => \N__33460\,
            I => \N__33456\
        );

    \I__7555\ : InMux
    port map (
            O => \N__33459\,
            I => \N__33453\
        );

    \I__7554\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33450\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__33453\,
            I => \b2v_inst20.counterZ0Z_31\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__33450\,
            I => \b2v_inst20.counterZ0Z_31\
        );

    \I__7551\ : InMux
    port map (
            O => \N__33445\,
            I => \N__33441\
        );

    \I__7550\ : InMux
    port map (
            O => \N__33444\,
            I => \N__33438\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__33441\,
            I => \b2v_inst20.counterZ0Z_30\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__33438\,
            I => \b2v_inst20.counterZ0Z_30\
        );

    \I__7547\ : InMux
    port map (
            O => \N__33433\,
            I => \N__33430\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__33430\,
            I => \N__33427\
        );

    \I__7545\ : Span4Mux_h
    port map (
            O => \N__33427\,
            I => \N__33424\
        );

    \I__7544\ : Odrv4
    port map (
            O => \N__33424\,
            I => \b2v_inst20.un4_counter_7_and\
        );

    \I__7543\ : InMux
    port map (
            O => \N__33421\,
            I => \N__33417\
        );

    \I__7542\ : InMux
    port map (
            O => \N__33420\,
            I => \N__33414\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__33417\,
            I => \b2v_inst20.counterZ0Z_11\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__33414\,
            I => \b2v_inst20.counterZ0Z_11\
        );

    \I__7539\ : InMux
    port map (
            O => \N__33409\,
            I => \N__33405\
        );

    \I__7538\ : InMux
    port map (
            O => \N__33408\,
            I => \N__33402\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__33405\,
            I => \b2v_inst20.counterZ0Z_8\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__33402\,
            I => \b2v_inst20.counterZ0Z_8\
        );

    \I__7535\ : CascadeMux
    port map (
            O => \N__33397\,
            I => \N__33393\
        );

    \I__7534\ : InMux
    port map (
            O => \N__33396\,
            I => \N__33390\
        );

    \I__7533\ : InMux
    port map (
            O => \N__33393\,
            I => \N__33387\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__33390\,
            I => \b2v_inst20.counterZ0Z_10\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__33387\,
            I => \b2v_inst20.counterZ0Z_10\
        );

    \I__7530\ : InMux
    port map (
            O => \N__33382\,
            I => \N__33378\
        );

    \I__7529\ : InMux
    port map (
            O => \N__33381\,
            I => \N__33375\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__33378\,
            I => \b2v_inst20.counterZ0Z_9\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__33375\,
            I => \b2v_inst20.counterZ0Z_9\
        );

    \I__7526\ : CascadeMux
    port map (
            O => \N__33370\,
            I => \N__33367\
        );

    \I__7525\ : InMux
    port map (
            O => \N__33367\,
            I => \N__33364\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__33364\,
            I => \N__33361\
        );

    \I__7523\ : Span4Mux_v
    port map (
            O => \N__33361\,
            I => \N__33358\
        );

    \I__7522\ : Odrv4
    port map (
            O => \N__33358\,
            I => \b2v_inst20.un4_counter_2_and\
        );

    \I__7521\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33351\
        );

    \I__7520\ : InMux
    port map (
            O => \N__33354\,
            I => \N__33348\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__33351\,
            I => \b2v_inst20.counterZ0Z_12\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__33348\,
            I => \b2v_inst20.counterZ0Z_12\
        );

    \I__7517\ : InMux
    port map (
            O => \N__33343\,
            I => \N__33339\
        );

    \I__7516\ : InMux
    port map (
            O => \N__33342\,
            I => \N__33336\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__33339\,
            I => \b2v_inst20.counterZ0Z_14\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__33336\,
            I => \b2v_inst20.counterZ0Z_14\
        );

    \I__7513\ : CascadeMux
    port map (
            O => \N__33331\,
            I => \N__33327\
        );

    \I__7512\ : InMux
    port map (
            O => \N__33330\,
            I => \N__33324\
        );

    \I__7511\ : InMux
    port map (
            O => \N__33327\,
            I => \N__33321\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__33324\,
            I => \b2v_inst20.counterZ0Z_15\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__33321\,
            I => \b2v_inst20.counterZ0Z_15\
        );

    \I__7508\ : InMux
    port map (
            O => \N__33316\,
            I => \N__33312\
        );

    \I__7507\ : InMux
    port map (
            O => \N__33315\,
            I => \N__33309\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__33312\,
            I => \b2v_inst20.counterZ0Z_13\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__33309\,
            I => \b2v_inst20.counterZ0Z_13\
        );

    \I__7504\ : InMux
    port map (
            O => \N__33304\,
            I => \N__33301\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__33301\,
            I => \N__33298\
        );

    \I__7502\ : Span4Mux_v
    port map (
            O => \N__33298\,
            I => \N__33295\
        );

    \I__7501\ : Odrv4
    port map (
            O => \N__33295\,
            I => \b2v_inst20.un4_counter_3_and\
        );

    \I__7500\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33288\
        );

    \I__7499\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33285\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__33288\,
            I => \b2v_inst20.counterZ0Z_19\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__33285\,
            I => \b2v_inst20.counterZ0Z_19\
        );

    \I__7496\ : InMux
    port map (
            O => \N__33280\,
            I => \N__33276\
        );

    \I__7495\ : InMux
    port map (
            O => \N__33279\,
            I => \N__33273\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__33276\,
            I => \b2v_inst20.counterZ0Z_16\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__33273\,
            I => \b2v_inst20.counterZ0Z_16\
        );

    \I__7492\ : CascadeMux
    port map (
            O => \N__33268\,
            I => \N__33264\
        );

    \I__7491\ : InMux
    port map (
            O => \N__33267\,
            I => \N__33261\
        );

    \I__7490\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33258\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__33261\,
            I => \b2v_inst20.counterZ0Z_17\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__33258\,
            I => \b2v_inst20.counterZ0Z_17\
        );

    \I__7487\ : InMux
    port map (
            O => \N__33253\,
            I => \N__33249\
        );

    \I__7486\ : InMux
    port map (
            O => \N__33252\,
            I => \N__33246\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__33249\,
            I => \b2v_inst20.counterZ0Z_18\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__33246\,
            I => \b2v_inst20.counterZ0Z_18\
        );

    \I__7483\ : CascadeMux
    port map (
            O => \N__33241\,
            I => \N__33238\
        );

    \I__7482\ : InMux
    port map (
            O => \N__33238\,
            I => \N__33235\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__33235\,
            I => \N__33232\
        );

    \I__7480\ : Span4Mux_h
    port map (
            O => \N__33232\,
            I => \N__33229\
        );

    \I__7479\ : Odrv4
    port map (
            O => \N__33229\,
            I => \b2v_inst20.un4_counter_4_and\
        );

    \I__7478\ : InMux
    port map (
            O => \N__33226\,
            I => \N__33222\
        );

    \I__7477\ : InMux
    port map (
            O => \N__33225\,
            I => \N__33219\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__33222\,
            I => \b2v_inst20.counterZ0Z_23\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__33219\,
            I => \b2v_inst20.counterZ0Z_23\
        );

    \I__7474\ : InMux
    port map (
            O => \N__33214\,
            I => \N__33210\
        );

    \I__7473\ : InMux
    port map (
            O => \N__33213\,
            I => \N__33207\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__33210\,
            I => \b2v_inst20.counterZ0Z_22\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__33207\,
            I => \b2v_inst20.counterZ0Z_22\
        );

    \I__7470\ : CascadeMux
    port map (
            O => \N__33202\,
            I => \N__33198\
        );

    \I__7469\ : InMux
    port map (
            O => \N__33201\,
            I => \N__33195\
        );

    \I__7468\ : InMux
    port map (
            O => \N__33198\,
            I => \N__33192\
        );

    \I__7467\ : LocalMux
    port map (
            O => \N__33195\,
            I => \b2v_inst20.counterZ0Z_21\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__33192\,
            I => \b2v_inst20.counterZ0Z_21\
        );

    \I__7465\ : InMux
    port map (
            O => \N__33187\,
            I => \N__33183\
        );

    \I__7464\ : InMux
    port map (
            O => \N__33186\,
            I => \N__33180\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__33183\,
            I => \b2v_inst20.counterZ0Z_20\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__33180\,
            I => \b2v_inst20.counterZ0Z_20\
        );

    \I__7461\ : CascadeMux
    port map (
            O => \N__33175\,
            I => \N__33172\
        );

    \I__7460\ : InMux
    port map (
            O => \N__33172\,
            I => \N__33169\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__33169\,
            I => \N__33166\
        );

    \I__7458\ : Span4Mux_h
    port map (
            O => \N__33166\,
            I => \N__33163\
        );

    \I__7457\ : Odrv4
    port map (
            O => \N__33163\,
            I => \b2v_inst20.un4_counter_5_and\
        );

    \I__7456\ : InMux
    port map (
            O => \N__33160\,
            I => \N__33156\
        );

    \I__7455\ : InMux
    port map (
            O => \N__33159\,
            I => \N__33153\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__33156\,
            I => \b2v_inst20.counterZ0Z_24\
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__33153\,
            I => \b2v_inst20.counterZ0Z_24\
        );

    \I__7452\ : InMux
    port map (
            O => \N__33148\,
            I => \N__33144\
        );

    \I__7451\ : InMux
    port map (
            O => \N__33147\,
            I => \N__33141\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__33144\,
            I => \N__33138\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__33141\,
            I => \b2v_inst20.counterZ0Z_27\
        );

    \I__7448\ : Odrv4
    port map (
            O => \N__33138\,
            I => \b2v_inst20.counterZ0Z_27\
        );

    \I__7447\ : CascadeMux
    port map (
            O => \N__33133\,
            I => \N__33130\
        );

    \I__7446\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33126\
        );

    \I__7445\ : InMux
    port map (
            O => \N__33129\,
            I => \N__33123\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__33126\,
            I => \N__33120\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__33123\,
            I => \b2v_inst20.counterZ0Z_25\
        );

    \I__7442\ : Odrv4
    port map (
            O => \N__33120\,
            I => \b2v_inst20.counterZ0Z_25\
        );

    \I__7441\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33111\
        );

    \I__7440\ : InMux
    port map (
            O => \N__33114\,
            I => \N__33108\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__33111\,
            I => \N__33105\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__33108\,
            I => \b2v_inst20.counterZ0Z_26\
        );

    \I__7437\ : Odrv4
    port map (
            O => \N__33105\,
            I => \b2v_inst20.counterZ0Z_26\
        );

    \I__7436\ : CascadeMux
    port map (
            O => \N__33100\,
            I => \N__33097\
        );

    \I__7435\ : InMux
    port map (
            O => \N__33097\,
            I => \N__33094\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__33094\,
            I => \N__33091\
        );

    \I__7433\ : Span4Mux_h
    port map (
            O => \N__33091\,
            I => \N__33088\
        );

    \I__7432\ : Odrv4
    port map (
            O => \N__33088\,
            I => \b2v_inst20.un4_counter_6_and\
        );

    \I__7431\ : CascadeMux
    port map (
            O => \N__33085\,
            I => \b2v_inst200.curr_stateZ0Z_1_cascade_\
        );

    \I__7430\ : InMux
    port map (
            O => \N__33082\,
            I => \N__33078\
        );

    \I__7429\ : InMux
    port map (
            O => \N__33081\,
            I => \N__33075\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__33078\,
            I => \N__33072\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__33075\,
            I => \N__33069\
        );

    \I__7426\ : Span4Mux_v
    port map (
            O => \N__33072\,
            I => \N__33066\
        );

    \I__7425\ : Span4Mux_h
    port map (
            O => \N__33069\,
            I => \N__33063\
        );

    \I__7424\ : Span4Mux_h
    port map (
            O => \N__33066\,
            I => \N__33060\
        );

    \I__7423\ : Span4Mux_h
    port map (
            O => \N__33063\,
            I => \N__33057\
        );

    \I__7422\ : Span4Mux_h
    port map (
            O => \N__33060\,
            I => \N__33054\
        );

    \I__7421\ : Odrv4
    port map (
            O => \N__33057\,
            I => \N_405\
        );

    \I__7420\ : Odrv4
    port map (
            O => \N__33054\,
            I => \N_405\
        );

    \I__7419\ : CascadeMux
    port map (
            O => \N__33049\,
            I => \b2v_inst5.count_rst_6_cascade_\
        );

    \I__7418\ : InMux
    port map (
            O => \N__33046\,
            I => \N__33041\
        );

    \I__7417\ : InMux
    port map (
            O => \N__33045\,
            I => \N__33038\
        );

    \I__7416\ : InMux
    port map (
            O => \N__33044\,
            I => \N__33035\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__33041\,
            I => \b2v_inst5.countZ0Z_8\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__33038\,
            I => \b2v_inst5.countZ0Z_8\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__33035\,
            I => \b2v_inst5.countZ0Z_8\
        );

    \I__7412\ : InMux
    port map (
            O => \N__33028\,
            I => \N__33022\
        );

    \I__7411\ : InMux
    port map (
            O => \N__33027\,
            I => \N__33022\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__33022\,
            I => \b2v_inst5.un2_count_1_cry_7_THRU_CO\
        );

    \I__7409\ : CascadeMux
    port map (
            O => \N__33019\,
            I => \b2v_inst5.countZ0Z_8_cascade_\
        );

    \I__7408\ : InMux
    port map (
            O => \N__33016\,
            I => \N__33013\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__33013\,
            I => \b2v_inst5.count_0_8\
        );

    \I__7406\ : InMux
    port map (
            O => \N__33010\,
            I => \N__33007\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__33007\,
            I => \b2v_inst5.count_rst_10\
        );

    \I__7404\ : CascadeMux
    port map (
            O => \N__33004\,
            I => \b2v_inst5.count_rst_10_cascade_\
        );

    \I__7403\ : CascadeMux
    port map (
            O => \N__33001\,
            I => \N__32998\
        );

    \I__7402\ : InMux
    port map (
            O => \N__32998\,
            I => \N__32994\
        );

    \I__7401\ : InMux
    port map (
            O => \N__32997\,
            I => \N__32991\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__32994\,
            I => \b2v_inst5.un2_count_1_axb_4\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__32991\,
            I => \b2v_inst5.un2_count_1_axb_4\
        );

    \I__7398\ : InMux
    port map (
            O => \N__32986\,
            I => \N__32980\
        );

    \I__7397\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32980\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__32980\,
            I => \b2v_inst5.un2_count_1_cry_3_THRU_CO\
        );

    \I__7395\ : CascadeMux
    port map (
            O => \N__32977\,
            I => \b2v_inst5.un2_count_1_axb_4_cascade_\
        );

    \I__7394\ : CascadeMux
    port map (
            O => \N__32974\,
            I => \N__32971\
        );

    \I__7393\ : InMux
    port map (
            O => \N__32971\,
            I => \N__32967\
        );

    \I__7392\ : InMux
    port map (
            O => \N__32970\,
            I => \N__32964\
        );

    \I__7391\ : LocalMux
    port map (
            O => \N__32967\,
            I => \b2v_inst5.count_0_4\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__32964\,
            I => \b2v_inst5.count_0_4\
        );

    \I__7389\ : InMux
    port map (
            O => \N__32959\,
            I => \N__32956\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__32956\,
            I => \N__32943\
        );

    \I__7387\ : InMux
    port map (
            O => \N__32955\,
            I => \N__32932\
        );

    \I__7386\ : InMux
    port map (
            O => \N__32954\,
            I => \N__32932\
        );

    \I__7385\ : InMux
    port map (
            O => \N__32953\,
            I => \N__32932\
        );

    \I__7384\ : InMux
    port map (
            O => \N__32952\,
            I => \N__32932\
        );

    \I__7383\ : InMux
    port map (
            O => \N__32951\,
            I => \N__32932\
        );

    \I__7382\ : InMux
    port map (
            O => \N__32950\,
            I => \N__32921\
        );

    \I__7381\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32921\
        );

    \I__7380\ : InMux
    port map (
            O => \N__32948\,
            I => \N__32921\
        );

    \I__7379\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32921\
        );

    \I__7378\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32921\
        );

    \I__7377\ : Span4Mux_v
    port map (
            O => \N__32943\,
            I => \N__32918\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__32932\,
            I => \N__32915\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__32921\,
            I => \b2v_inst5.N_390\
        );

    \I__7374\ : Odrv4
    port map (
            O => \N__32918\,
            I => \b2v_inst5.N_390\
        );

    \I__7373\ : Odrv4
    port map (
            O => \N__32915\,
            I => \b2v_inst5.N_390\
        );

    \I__7372\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32905\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__32905\,
            I => \N__32901\
        );

    \I__7370\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32898\
        );

    \I__7369\ : Odrv4
    port map (
            O => \N__32901\,
            I => \b2v_inst5.un2_count_1_cry_12_THRU_CO\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__32898\,
            I => \b2v_inst5.un2_count_1_cry_12_THRU_CO\
        );

    \I__7367\ : SRMux
    port map (
            O => \N__32893\,
            I => \N__32889\
        );

    \I__7366\ : SRMux
    port map (
            O => \N__32892\,
            I => \N__32886\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__32889\,
            I => \N__32877\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__32886\,
            I => \N__32874\
        );

    \I__7363\ : SRMux
    port map (
            O => \N__32885\,
            I => \N__32871\
        );

    \I__7362\ : CascadeMux
    port map (
            O => \N__32884\,
            I => \N__32862\
        );

    \I__7361\ : CascadeMux
    port map (
            O => \N__32883\,
            I => \N__32858\
        );

    \I__7360\ : SRMux
    port map (
            O => \N__32882\,
            I => \N__32855\
        );

    \I__7359\ : SRMux
    port map (
            O => \N__32881\,
            I => \N__32852\
        );

    \I__7358\ : SRMux
    port map (
            O => \N__32880\,
            I => \N__32849\
        );

    \I__7357\ : Span4Mux_h
    port map (
            O => \N__32877\,
            I => \N__32842\
        );

    \I__7356\ : Span4Mux_v
    port map (
            O => \N__32874\,
            I => \N__32842\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__32871\,
            I => \N__32842\
        );

    \I__7354\ : CascadeMux
    port map (
            O => \N__32870\,
            I => \N__32836\
        );

    \I__7353\ : CascadeMux
    port map (
            O => \N__32869\,
            I => \N__32829\
        );

    \I__7352\ : CascadeMux
    port map (
            O => \N__32868\,
            I => \N__32825\
        );

    \I__7351\ : SRMux
    port map (
            O => \N__32867\,
            I => \N__32822\
        );

    \I__7350\ : InMux
    port map (
            O => \N__32866\,
            I => \N__32819\
        );

    \I__7349\ : InMux
    port map (
            O => \N__32865\,
            I => \N__32810\
        );

    \I__7348\ : InMux
    port map (
            O => \N__32862\,
            I => \N__32810\
        );

    \I__7347\ : InMux
    port map (
            O => \N__32861\,
            I => \N__32810\
        );

    \I__7346\ : InMux
    port map (
            O => \N__32858\,
            I => \N__32810\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__32855\,
            I => \N__32799\
        );

    \I__7344\ : LocalMux
    port map (
            O => \N__32852\,
            I => \N__32794\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__32849\,
            I => \N__32794\
        );

    \I__7342\ : Span4Mux_v
    port map (
            O => \N__32842\,
            I => \N__32791\
        );

    \I__7341\ : InMux
    port map (
            O => \N__32841\,
            I => \N__32786\
        );

    \I__7340\ : InMux
    port map (
            O => \N__32840\,
            I => \N__32786\
        );

    \I__7339\ : InMux
    port map (
            O => \N__32839\,
            I => \N__32779\
        );

    \I__7338\ : InMux
    port map (
            O => \N__32836\,
            I => \N__32779\
        );

    \I__7337\ : InMux
    port map (
            O => \N__32835\,
            I => \N__32779\
        );

    \I__7336\ : InMux
    port map (
            O => \N__32834\,
            I => \N__32772\
        );

    \I__7335\ : InMux
    port map (
            O => \N__32833\,
            I => \N__32772\
        );

    \I__7334\ : InMux
    port map (
            O => \N__32832\,
            I => \N__32772\
        );

    \I__7333\ : InMux
    port map (
            O => \N__32829\,
            I => \N__32765\
        );

    \I__7332\ : InMux
    port map (
            O => \N__32828\,
            I => \N__32765\
        );

    \I__7331\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32765\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__32822\,
            I => \N__32762\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__32819\,
            I => \N__32757\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__32810\,
            I => \N__32757\
        );

    \I__7327\ : InMux
    port map (
            O => \N__32809\,
            I => \N__32752\
        );

    \I__7326\ : InMux
    port map (
            O => \N__32808\,
            I => \N__32752\
        );

    \I__7325\ : InMux
    port map (
            O => \N__32807\,
            I => \N__32747\
        );

    \I__7324\ : InMux
    port map (
            O => \N__32806\,
            I => \N__32747\
        );

    \I__7323\ : InMux
    port map (
            O => \N__32805\,
            I => \N__32742\
        );

    \I__7322\ : InMux
    port map (
            O => \N__32804\,
            I => \N__32742\
        );

    \I__7321\ : InMux
    port map (
            O => \N__32803\,
            I => \N__32737\
        );

    \I__7320\ : InMux
    port map (
            O => \N__32802\,
            I => \N__32737\
        );

    \I__7319\ : Span4Mux_v
    port map (
            O => \N__32799\,
            I => \N__32730\
        );

    \I__7318\ : Span4Mux_v
    port map (
            O => \N__32794\,
            I => \N__32730\
        );

    \I__7317\ : Span4Mux_s0_h
    port map (
            O => \N__32791\,
            I => \N__32730\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__32786\,
            I => \N__32725\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__32779\,
            I => \N__32725\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__32772\,
            I => \N__32720\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__32765\,
            I => \N__32720\
        );

    \I__7312\ : Span4Mux_v
    port map (
            O => \N__32762\,
            I => \N__32707\
        );

    \I__7311\ : Span4Mux_s1_h
    port map (
            O => \N__32757\,
            I => \N__32707\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__32752\,
            I => \N__32707\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__32747\,
            I => \N__32707\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__32742\,
            I => \N__32707\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__32737\,
            I => \N__32707\
        );

    \I__7306\ : Span4Mux_h
    port map (
            O => \N__32730\,
            I => \N__32704\
        );

    \I__7305\ : Span4Mux_s3_h
    port map (
            O => \N__32725\,
            I => \N__32701\
        );

    \I__7304\ : Span4Mux_s3_h
    port map (
            O => \N__32720\,
            I => \N__32698\
        );

    \I__7303\ : Span4Mux_v
    port map (
            O => \N__32707\,
            I => \N__32695\
        );

    \I__7302\ : Odrv4
    port map (
            O => \N__32704\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__7301\ : Odrv4
    port map (
            O => \N__32701\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__7300\ : Odrv4
    port map (
            O => \N__32698\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__7299\ : Odrv4
    port map (
            O => \N__32695\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__7298\ : CEMux
    port map (
            O => \N__32686\,
            I => \N__32683\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__32683\,
            I => \N__32675\
        );

    \I__7296\ : InMux
    port map (
            O => \N__32682\,
            I => \N__32668\
        );

    \I__7295\ : InMux
    port map (
            O => \N__32681\,
            I => \N__32668\
        );

    \I__7294\ : CEMux
    port map (
            O => \N__32680\,
            I => \N__32668\
        );

    \I__7293\ : CEMux
    port map (
            O => \N__32679\,
            I => \N__32665\
        );

    \I__7292\ : CascadeMux
    port map (
            O => \N__32678\,
            I => \N__32661\
        );

    \I__7291\ : Span4Mux_s3_v
    port map (
            O => \N__32675\,
            I => \N__32652\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__32668\,
            I => \N__32652\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__32665\,
            I => \N__32652\
        );

    \I__7288\ : CascadeMux
    port map (
            O => \N__32664\,
            I => \N__32638\
        );

    \I__7287\ : InMux
    port map (
            O => \N__32661\,
            I => \N__32626\
        );

    \I__7286\ : CEMux
    port map (
            O => \N__32660\,
            I => \N__32626\
        );

    \I__7285\ : CEMux
    port map (
            O => \N__32659\,
            I => \N__32623\
        );

    \I__7284\ : Span4Mux_v
    port map (
            O => \N__32652\,
            I => \N__32620\
        );

    \I__7283\ : InMux
    port map (
            O => \N__32651\,
            I => \N__32615\
        );

    \I__7282\ : InMux
    port map (
            O => \N__32650\,
            I => \N__32615\
        );

    \I__7281\ : InMux
    port map (
            O => \N__32649\,
            I => \N__32608\
        );

    \I__7280\ : InMux
    port map (
            O => \N__32648\,
            I => \N__32608\
        );

    \I__7279\ : InMux
    port map (
            O => \N__32647\,
            I => \N__32608\
        );

    \I__7278\ : CEMux
    port map (
            O => \N__32646\,
            I => \N__32599\
        );

    \I__7277\ : InMux
    port map (
            O => \N__32645\,
            I => \N__32599\
        );

    \I__7276\ : InMux
    port map (
            O => \N__32644\,
            I => \N__32599\
        );

    \I__7275\ : InMux
    port map (
            O => \N__32643\,
            I => \N__32599\
        );

    \I__7274\ : InMux
    port map (
            O => \N__32642\,
            I => \N__32596\
        );

    \I__7273\ : InMux
    port map (
            O => \N__32641\,
            I => \N__32589\
        );

    \I__7272\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32589\
        );

    \I__7271\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32589\
        );

    \I__7270\ : InMux
    port map (
            O => \N__32636\,
            I => \N__32584\
        );

    \I__7269\ : CEMux
    port map (
            O => \N__32635\,
            I => \N__32584\
        );

    \I__7268\ : InMux
    port map (
            O => \N__32634\,
            I => \N__32581\
        );

    \I__7267\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32574\
        );

    \I__7266\ : InMux
    port map (
            O => \N__32632\,
            I => \N__32574\
        );

    \I__7265\ : InMux
    port map (
            O => \N__32631\,
            I => \N__32574\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__32626\,
            I => \N__32571\
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__32623\,
            I => \N__32556\
        );

    \I__7262\ : Span4Mux_s0_h
    port map (
            O => \N__32620\,
            I => \N__32556\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__32615\,
            I => \N__32556\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__32608\,
            I => \N__32556\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__32599\,
            I => \N__32556\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__32596\,
            I => \N__32556\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__32589\,
            I => \N__32556\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__32584\,
            I => \N__32553\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__32581\,
            I => \N__32548\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__32574\,
            I => \N__32548\
        );

    \I__7253\ : Span4Mux_s2_h
    port map (
            O => \N__32571\,
            I => \N__32543\
        );

    \I__7252\ : Span4Mux_v
    port map (
            O => \N__32556\,
            I => \N__32540\
        );

    \I__7251\ : Span4Mux_s2_h
    port map (
            O => \N__32553\,
            I => \N__32535\
        );

    \I__7250\ : Span4Mux_s2_h
    port map (
            O => \N__32548\,
            I => \N__32535\
        );

    \I__7249\ : InMux
    port map (
            O => \N__32547\,
            I => \N__32530\
        );

    \I__7248\ : InMux
    port map (
            O => \N__32546\,
            I => \N__32530\
        );

    \I__7247\ : Odrv4
    port map (
            O => \N__32543\,
            I => \b2v_inst5.count_enZ0\
        );

    \I__7246\ : Odrv4
    port map (
            O => \N__32540\,
            I => \b2v_inst5.count_enZ0\
        );

    \I__7245\ : Odrv4
    port map (
            O => \N__32535\,
            I => \b2v_inst5.count_enZ0\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__32530\,
            I => \b2v_inst5.count_enZ0\
        );

    \I__7243\ : CascadeMux
    port map (
            O => \N__32521\,
            I => \b2v_inst5.count_rst_1_cascade_\
        );

    \I__7242\ : InMux
    port map (
            O => \N__32518\,
            I => \N__32515\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__32515\,
            I => \N__32512\
        );

    \I__7240\ : Odrv12
    port map (
            O => \N__32512\,
            I => \b2v_inst5.count_0_13\
        );

    \I__7239\ : InMux
    port map (
            O => \N__32509\,
            I => \N__32506\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__32506\,
            I => \N__32501\
        );

    \I__7237\ : CascadeMux
    port map (
            O => \N__32505\,
            I => \N__32497\
        );

    \I__7236\ : InMux
    port map (
            O => \N__32504\,
            I => \N__32494\
        );

    \I__7235\ : Span4Mux_v
    port map (
            O => \N__32501\,
            I => \N__32491\
        );

    \I__7234\ : InMux
    port map (
            O => \N__32500\,
            I => \N__32488\
        );

    \I__7233\ : InMux
    port map (
            O => \N__32497\,
            I => \N__32485\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__32494\,
            I => \N__32482\
        );

    \I__7231\ : Odrv4
    port map (
            O => \N__32491\,
            I => \b2v_inst5.countZ0Z_13\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__32488\,
            I => \b2v_inst5.countZ0Z_13\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__32485\,
            I => \b2v_inst5.countZ0Z_13\
        );

    \I__7228\ : Odrv12
    port map (
            O => \N__32482\,
            I => \b2v_inst5.countZ0Z_13\
        );

    \I__7227\ : CascadeMux
    port map (
            O => \N__32473\,
            I => \N__32470\
        );

    \I__7226\ : InMux
    port map (
            O => \N__32470\,
            I => \N__32466\
        );

    \I__7225\ : InMux
    port map (
            O => \N__32469\,
            I => \N__32463\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__32466\,
            I => \N__32460\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__32463\,
            I => \b2v_inst5.countZ0Z_3\
        );

    \I__7222\ : Odrv4
    port map (
            O => \N__32460\,
            I => \b2v_inst5.countZ0Z_3\
        );

    \I__7221\ : InMux
    port map (
            O => \N__32455\,
            I => \N__32452\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__32452\,
            I => \N__32449\
        );

    \I__7219\ : Odrv12
    port map (
            O => \N__32449\,
            I => \b2v_inst5.count_1_i_a2_6_0\
        );

    \I__7218\ : CascadeMux
    port map (
            O => \N__32446\,
            I => \b2v_inst5.count_1_i_a2_4_0_cascade_\
        );

    \I__7217\ : InMux
    port map (
            O => \N__32443\,
            I => \N__32438\
        );

    \I__7216\ : InMux
    port map (
            O => \N__32442\,
            I => \N__32433\
        );

    \I__7215\ : InMux
    port map (
            O => \N__32441\,
            I => \N__32433\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__32438\,
            I => \N__32430\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__32433\,
            I => \b2v_inst5.count_1_i_a2_12_0\
        );

    \I__7212\ : Odrv4
    port map (
            O => \N__32430\,
            I => \b2v_inst5.count_1_i_a2_12_0\
        );

    \I__7211\ : InMux
    port map (
            O => \N__32425\,
            I => \N__32419\
        );

    \I__7210\ : InMux
    port map (
            O => \N__32424\,
            I => \N__32419\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__32419\,
            I => \b2v_inst5.count_0_2\
        );

    \I__7208\ : InMux
    port map (
            O => \N__32416\,
            I => \N__32407\
        );

    \I__7207\ : InMux
    port map (
            O => \N__32415\,
            I => \N__32407\
        );

    \I__7206\ : InMux
    port map (
            O => \N__32414\,
            I => \N__32407\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__32407\,
            I => \b2v_inst5.count_rst_12\
        );

    \I__7204\ : InMux
    port map (
            O => \N__32404\,
            I => \N__32401\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__32401\,
            I => \b2v_inst5.un2_count_1_axb_2\
        );

    \I__7202\ : CascadeMux
    port map (
            O => \N__32398\,
            I => \N__32393\
        );

    \I__7201\ : InMux
    port map (
            O => \N__32397\,
            I => \N__32390\
        );

    \I__7200\ : InMux
    port map (
            O => \N__32396\,
            I => \N__32387\
        );

    \I__7199\ : InMux
    port map (
            O => \N__32393\,
            I => \N__32384\
        );

    \I__7198\ : LocalMux
    port map (
            O => \N__32390\,
            I => \b2v_inst5.countZ0Z_1\
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__32387\,
            I => \b2v_inst5.countZ0Z_1\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__32384\,
            I => \b2v_inst5.countZ0Z_1\
        );

    \I__7195\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32374\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__32374\,
            I => \b2v_inst5.count_1_i_a2_3_0\
        );

    \I__7193\ : CascadeMux
    port map (
            O => \N__32371\,
            I => \N__32368\
        );

    \I__7192\ : InMux
    port map (
            O => \N__32368\,
            I => \N__32362\
        );

    \I__7191\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32362\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__32362\,
            I => \b2v_inst5.count_0_11\
        );

    \I__7189\ : InMux
    port map (
            O => \N__32359\,
            I => \N__32350\
        );

    \I__7188\ : InMux
    port map (
            O => \N__32358\,
            I => \N__32350\
        );

    \I__7187\ : InMux
    port map (
            O => \N__32357\,
            I => \N__32350\
        );

    \I__7186\ : LocalMux
    port map (
            O => \N__32350\,
            I => \b2v_inst5.count_rst_3\
        );

    \I__7185\ : InMux
    port map (
            O => \N__32347\,
            I => \N__32344\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__32344\,
            I => \b2v_inst5.un2_count_1_axb_11\
        );

    \I__7183\ : InMux
    port map (
            O => \N__32341\,
            I => \N__32338\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__32338\,
            I => \b2v_inst5.count_1_i_a2_5_0\
        );

    \I__7181\ : CascadeMux
    port map (
            O => \N__32335\,
            I => \b2v_inst5.count_RNIRHC7IZ0Z_2_cascade_\
        );

    \I__7180\ : InMux
    port map (
            O => \N__32332\,
            I => \N__32328\
        );

    \I__7179\ : InMux
    port map (
            O => \N__32331\,
            I => \N__32325\
        );

    \I__7178\ : LocalMux
    port map (
            O => \N__32328\,
            I => \b2v_inst5.countZ0Z_0\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__32325\,
            I => \b2v_inst5.countZ0Z_0\
        );

    \I__7176\ : CascadeMux
    port map (
            O => \N__32320\,
            I => \b2v_inst5.countZ0Z_0_cascade_\
        );

    \I__7175\ : CascadeMux
    port map (
            O => \N__32317\,
            I => \b2v_inst5.count_RNIZ0Z_0_cascade_\
        );

    \I__7174\ : InMux
    port map (
            O => \N__32314\,
            I => \N__32311\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__32311\,
            I => \b2v_inst5.count_RNIZ0Z_0\
        );

    \I__7172\ : InMux
    port map (
            O => \N__32308\,
            I => \N__32305\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__32305\,
            I => \b2v_inst5.count_0_1\
        );

    \I__7170\ : InMux
    port map (
            O => \N__32302\,
            I => \N__32299\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__32299\,
            I => \N__32294\
        );

    \I__7168\ : InMux
    port map (
            O => \N__32298\,
            I => \N__32289\
        );

    \I__7167\ : InMux
    port map (
            O => \N__32297\,
            I => \N__32289\
        );

    \I__7166\ : Odrv4
    port map (
            O => \N__32294\,
            I => \b2v_inst5.count_1_i_a2_11_0\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__32289\,
            I => \b2v_inst5.count_1_i_a2_11_0\
        );

    \I__7164\ : InMux
    port map (
            O => \N__32284\,
            I => \N__32278\
        );

    \I__7163\ : InMux
    port map (
            O => \N__32283\,
            I => \N__32278\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__32278\,
            I => \b2v_inst5.N_2906_i\
        );

    \I__7161\ : InMux
    port map (
            O => \N__32275\,
            I => \N__32272\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__32272\,
            I => \b2v_inst5.count_0_0\
        );

    \I__7159\ : CascadeMux
    port map (
            O => \N__32269\,
            I => \N__32266\
        );

    \I__7158\ : InMux
    port map (
            O => \N__32266\,
            I => \N__32263\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__32263\,
            I => \b2v_inst5.count_0_3\
        );

    \I__7156\ : InMux
    port map (
            O => \N__32260\,
            I => \N__32254\
        );

    \I__7155\ : InMux
    port map (
            O => \N__32259\,
            I => \N__32254\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__32254\,
            I => \b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9\
        );

    \I__7153\ : InMux
    port map (
            O => \N__32251\,
            I => \N__32248\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__32248\,
            I => \b2v_inst36.count_rst_14\
        );

    \I__7151\ : InMux
    port map (
            O => \N__32245\,
            I => \N__32242\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__32242\,
            I => \N__32238\
        );

    \I__7149\ : InMux
    port map (
            O => \N__32241\,
            I => \N__32232\
        );

    \I__7148\ : Span4Mux_s1_v
    port map (
            O => \N__32238\,
            I => \N__32229\
        );

    \I__7147\ : InMux
    port map (
            O => \N__32237\,
            I => \N__32222\
        );

    \I__7146\ : InMux
    port map (
            O => \N__32236\,
            I => \N__32222\
        );

    \I__7145\ : InMux
    port map (
            O => \N__32235\,
            I => \N__32222\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__32232\,
            I => \b2v_inst36.countZ0Z_0\
        );

    \I__7143\ : Odrv4
    port map (
            O => \N__32229\,
            I => \b2v_inst36.countZ0Z_0\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__32222\,
            I => \b2v_inst36.countZ0Z_0\
        );

    \I__7141\ : InMux
    port map (
            O => \N__32215\,
            I => \N__32209\
        );

    \I__7140\ : InMux
    port map (
            O => \N__32214\,
            I => \N__32209\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__32209\,
            I => \N__32202\
        );

    \I__7138\ : InMux
    port map (
            O => \N__32208\,
            I => \N__32190\
        );

    \I__7137\ : InMux
    port map (
            O => \N__32207\,
            I => \N__32183\
        );

    \I__7136\ : InMux
    port map (
            O => \N__32206\,
            I => \N__32183\
        );

    \I__7135\ : InMux
    port map (
            O => \N__32205\,
            I => \N__32183\
        );

    \I__7134\ : Span4Mux_s1_v
    port map (
            O => \N__32202\,
            I => \N__32174\
        );

    \I__7133\ : InMux
    port map (
            O => \N__32201\,
            I => \N__32167\
        );

    \I__7132\ : InMux
    port map (
            O => \N__32200\,
            I => \N__32167\
        );

    \I__7131\ : InMux
    port map (
            O => \N__32199\,
            I => \N__32167\
        );

    \I__7130\ : InMux
    port map (
            O => \N__32198\,
            I => \N__32160\
        );

    \I__7129\ : InMux
    port map (
            O => \N__32197\,
            I => \N__32160\
        );

    \I__7128\ : InMux
    port map (
            O => \N__32196\,
            I => \N__32160\
        );

    \I__7127\ : InMux
    port map (
            O => \N__32195\,
            I => \N__32153\
        );

    \I__7126\ : InMux
    port map (
            O => \N__32194\,
            I => \N__32153\
        );

    \I__7125\ : InMux
    port map (
            O => \N__32193\,
            I => \N__32153\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__32190\,
            I => \N__32148\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__32183\,
            I => \N__32148\
        );

    \I__7122\ : InMux
    port map (
            O => \N__32182\,
            I => \N__32140\
        );

    \I__7121\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32137\
        );

    \I__7120\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32128\
        );

    \I__7119\ : InMux
    port map (
            O => \N__32179\,
            I => \N__32128\
        );

    \I__7118\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32128\
        );

    \I__7117\ : InMux
    port map (
            O => \N__32177\,
            I => \N__32128\
        );

    \I__7116\ : Span4Mux_h
    port map (
            O => \N__32174\,
            I => \N__32125\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__32167\,
            I => \N__32116\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__32160\,
            I => \N__32116\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__32153\,
            I => \N__32116\
        );

    \I__7112\ : Span12Mux_s1_v
    port map (
            O => \N__32148\,
            I => \N__32116\
        );

    \I__7111\ : InMux
    port map (
            O => \N__32147\,
            I => \N__32105\
        );

    \I__7110\ : InMux
    port map (
            O => \N__32146\,
            I => \N__32105\
        );

    \I__7109\ : InMux
    port map (
            O => \N__32145\,
            I => \N__32105\
        );

    \I__7108\ : InMux
    port map (
            O => \N__32144\,
            I => \N__32105\
        );

    \I__7107\ : InMux
    port map (
            O => \N__32143\,
            I => \N__32105\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__32140\,
            I => \b2v_inst36.N_2928_i\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__32137\,
            I => \b2v_inst36.N_2928_i\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__32128\,
            I => \b2v_inst36.N_2928_i\
        );

    \I__7103\ : Odrv4
    port map (
            O => \N__32125\,
            I => \b2v_inst36.N_2928_i\
        );

    \I__7102\ : Odrv12
    port map (
            O => \N__32116\,
            I => \b2v_inst36.N_2928_i\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__32105\,
            I => \b2v_inst36.N_2928_i\
        );

    \I__7100\ : CascadeMux
    port map (
            O => \N__32092\,
            I => \b2v_inst36.countZ0Z_0_cascade_\
        );

    \I__7099\ : CascadeMux
    port map (
            O => \N__32089\,
            I => \N__32077\
        );

    \I__7098\ : InMux
    port map (
            O => \N__32088\,
            I => \N__32066\
        );

    \I__7097\ : InMux
    port map (
            O => \N__32087\,
            I => \N__32066\
        );

    \I__7096\ : InMux
    port map (
            O => \N__32086\,
            I => \N__32066\
        );

    \I__7095\ : InMux
    port map (
            O => \N__32085\,
            I => \N__32066\
        );

    \I__7094\ : InMux
    port map (
            O => \N__32084\,
            I => \N__32066\
        );

    \I__7093\ : InMux
    port map (
            O => \N__32083\,
            I => \N__32057\
        );

    \I__7092\ : InMux
    port map (
            O => \N__32082\,
            I => \N__32057\
        );

    \I__7091\ : InMux
    port map (
            O => \N__32081\,
            I => \N__32057\
        );

    \I__7090\ : InMux
    port map (
            O => \N__32080\,
            I => \N__32057\
        );

    \I__7089\ : InMux
    port map (
            O => \N__32077\,
            I => \N__32048\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__32066\,
            I => \N__32043\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__32057\,
            I => \N__32043\
        );

    \I__7086\ : CascadeMux
    port map (
            O => \N__32056\,
            I => \N__32039\
        );

    \I__7085\ : CascadeMux
    port map (
            O => \N__32055\,
            I => \N__32035\
        );

    \I__7084\ : InMux
    port map (
            O => \N__32054\,
            I => \N__32030\
        );

    \I__7083\ : InMux
    port map (
            O => \N__32053\,
            I => \N__32027\
        );

    \I__7082\ : InMux
    port map (
            O => \N__32052\,
            I => \N__32024\
        );

    \I__7081\ : InMux
    port map (
            O => \N__32051\,
            I => \N__32021\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__32048\,
            I => \N__32018\
        );

    \I__7079\ : Span4Mux_s1_v
    port map (
            O => \N__32043\,
            I => \N__32015\
        );

    \I__7078\ : InMux
    port map (
            O => \N__32042\,
            I => \N__32008\
        );

    \I__7077\ : InMux
    port map (
            O => \N__32039\,
            I => \N__32008\
        );

    \I__7076\ : InMux
    port map (
            O => \N__32038\,
            I => \N__32008\
        );

    \I__7075\ : InMux
    port map (
            O => \N__32035\,
            I => \N__32001\
        );

    \I__7074\ : InMux
    port map (
            O => \N__32034\,
            I => \N__32001\
        );

    \I__7073\ : InMux
    port map (
            O => \N__32033\,
            I => \N__32001\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__32030\,
            I => \b2v_inst36.N_1_i\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__32027\,
            I => \b2v_inst36.N_1_i\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__32024\,
            I => \b2v_inst36.N_1_i\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__32021\,
            I => \b2v_inst36.N_1_i\
        );

    \I__7068\ : Odrv12
    port map (
            O => \N__32018\,
            I => \b2v_inst36.N_1_i\
        );

    \I__7067\ : Odrv4
    port map (
            O => \N__32015\,
            I => \b2v_inst36.N_1_i\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__32008\,
            I => \b2v_inst36.N_1_i\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__32001\,
            I => \b2v_inst36.N_1_i\
        );

    \I__7064\ : InMux
    port map (
            O => \N__31984\,
            I => \N__31981\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__31981\,
            I => \b2v_inst36.count_1_0\
        );

    \I__7062\ : CascadeMux
    port map (
            O => \N__31978\,
            I => \N__31971\
        );

    \I__7061\ : CEMux
    port map (
            O => \N__31977\,
            I => \N__31967\
        );

    \I__7060\ : CEMux
    port map (
            O => \N__31976\,
            I => \N__31955\
        );

    \I__7059\ : CEMux
    port map (
            O => \N__31975\,
            I => \N__31946\
        );

    \I__7058\ : InMux
    port map (
            O => \N__31974\,
            I => \N__31946\
        );

    \I__7057\ : InMux
    port map (
            O => \N__31971\,
            I => \N__31946\
        );

    \I__7056\ : InMux
    port map (
            O => \N__31970\,
            I => \N__31946\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__31967\,
            I => \N__31943\
        );

    \I__7054\ : InMux
    port map (
            O => \N__31966\,
            I => \N__31936\
        );

    \I__7053\ : InMux
    port map (
            O => \N__31965\,
            I => \N__31936\
        );

    \I__7052\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31936\
        );

    \I__7051\ : InMux
    port map (
            O => \N__31963\,
            I => \N__31929\
        );

    \I__7050\ : CEMux
    port map (
            O => \N__31962\,
            I => \N__31926\
        );

    \I__7049\ : InMux
    port map (
            O => \N__31961\,
            I => \N__31921\
        );

    \I__7048\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31921\
        );

    \I__7047\ : InMux
    port map (
            O => \N__31959\,
            I => \N__31916\
        );

    \I__7046\ : CEMux
    port map (
            O => \N__31958\,
            I => \N__31916\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__31955\,
            I => \N__31912\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__31946\,
            I => \N__31909\
        );

    \I__7043\ : Span4Mux_s2_v
    port map (
            O => \N__31943\,
            I => \N__31904\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__31936\,
            I => \N__31901\
        );

    \I__7041\ : CEMux
    port map (
            O => \N__31935\,
            I => \N__31892\
        );

    \I__7040\ : InMux
    port map (
            O => \N__31934\,
            I => \N__31892\
        );

    \I__7039\ : InMux
    port map (
            O => \N__31933\,
            I => \N__31892\
        );

    \I__7038\ : InMux
    port map (
            O => \N__31932\,
            I => \N__31892\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__31929\,
            I => \N__31889\
        );

    \I__7036\ : LocalMux
    port map (
            O => \N__31926\,
            I => \N__31884\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__31921\,
            I => \N__31884\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__31916\,
            I => \N__31881\
        );

    \I__7033\ : InMux
    port map (
            O => \N__31915\,
            I => \N__31878\
        );

    \I__7032\ : Span4Mux_s2_v
    port map (
            O => \N__31912\,
            I => \N__31873\
        );

    \I__7031\ : Span4Mux_s2_v
    port map (
            O => \N__31909\,
            I => \N__31873\
        );

    \I__7030\ : InMux
    port map (
            O => \N__31908\,
            I => \N__31868\
        );

    \I__7029\ : InMux
    port map (
            O => \N__31907\,
            I => \N__31868\
        );

    \I__7028\ : Span4Mux_s1_h
    port map (
            O => \N__31904\,
            I => \N__31863\
        );

    \I__7027\ : Span4Mux_s2_v
    port map (
            O => \N__31901\,
            I => \N__31863\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__31892\,
            I => \N__31860\
        );

    \I__7025\ : Span4Mux_s3_h
    port map (
            O => \N__31889\,
            I => \N__31855\
        );

    \I__7024\ : Span4Mux_s3_h
    port map (
            O => \N__31884\,
            I => \N__31855\
        );

    \I__7023\ : Odrv4
    port map (
            O => \N__31881\,
            I => \b2v_inst36.count_en\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__31878\,
            I => \b2v_inst36.count_en\
        );

    \I__7021\ : Odrv4
    port map (
            O => \N__31873\,
            I => \b2v_inst36.count_en\
        );

    \I__7020\ : LocalMux
    port map (
            O => \N__31868\,
            I => \b2v_inst36.count_en\
        );

    \I__7019\ : Odrv4
    port map (
            O => \N__31863\,
            I => \b2v_inst36.count_en\
        );

    \I__7018\ : Odrv4
    port map (
            O => \N__31860\,
            I => \b2v_inst36.count_en\
        );

    \I__7017\ : Odrv4
    port map (
            O => \N__31855\,
            I => \b2v_inst36.count_en\
        );

    \I__7016\ : SRMux
    port map (
            O => \N__31840\,
            I => \N__31837\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__31837\,
            I => \N__31832\
        );

    \I__7014\ : SRMux
    port map (
            O => \N__31836\,
            I => \N__31829\
        );

    \I__7013\ : SRMux
    port map (
            O => \N__31835\,
            I => \N__31824\
        );

    \I__7012\ : Span4Mux_h
    port map (
            O => \N__31832\,
            I => \N__31819\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__31829\,
            I => \N__31819\
        );

    \I__7010\ : SRMux
    port map (
            O => \N__31828\,
            I => \N__31816\
        );

    \I__7009\ : SRMux
    port map (
            O => \N__31827\,
            I => \N__31812\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__31824\,
            I => \N__31809\
        );

    \I__7007\ : Span4Mux_s1_h
    port map (
            O => \N__31819\,
            I => \N__31804\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__31816\,
            I => \N__31804\
        );

    \I__7005\ : SRMux
    port map (
            O => \N__31815\,
            I => \N__31801\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__31812\,
            I => \N__31797\
        );

    \I__7003\ : Span4Mux_h
    port map (
            O => \N__31809\,
            I => \N__31794\
        );

    \I__7002\ : Span4Mux_s1_v
    port map (
            O => \N__31804\,
            I => \N__31789\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__31801\,
            I => \N__31789\
        );

    \I__7000\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31786\
        );

    \I__6999\ : Span4Mux_s2_v
    port map (
            O => \N__31797\,
            I => \N__31782\
        );

    \I__6998\ : Span4Mux_s2_v
    port map (
            O => \N__31794\,
            I => \N__31779\
        );

    \I__6997\ : Span4Mux_s1_h
    port map (
            O => \N__31789\,
            I => \N__31776\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__31786\,
            I => \N__31773\
        );

    \I__6995\ : InMux
    port map (
            O => \N__31785\,
            I => \N__31770\
        );

    \I__6994\ : Odrv4
    port map (
            O => \N__31782\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__6993\ : Odrv4
    port map (
            O => \N__31779\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__6992\ : Odrv4
    port map (
            O => \N__31776\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__6991\ : Odrv4
    port map (
            O => \N__31773\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__31770\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__6989\ : InMux
    port map (
            O => \N__31759\,
            I => \N__31756\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__31756\,
            I => \b2v_inst5.count_rst_5\
        );

    \I__6987\ : CascadeMux
    port map (
            O => \N__31753\,
            I => \b2v_inst5.count_rst_5_cascade_\
        );

    \I__6986\ : InMux
    port map (
            O => \N__31750\,
            I => \N__31747\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__31747\,
            I => \N__31744\
        );

    \I__6984\ : Span4Mux_v
    port map (
            O => \N__31744\,
            I => \N__31740\
        );

    \I__6983\ : InMux
    port map (
            O => \N__31743\,
            I => \N__31737\
        );

    \I__6982\ : Odrv4
    port map (
            O => \N__31740\,
            I => \b2v_inst5.un2_count_1_axb_9\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__31737\,
            I => \b2v_inst5.un2_count_1_axb_9\
        );

    \I__6980\ : InMux
    port map (
            O => \N__31732\,
            I => \N__31726\
        );

    \I__6979\ : InMux
    port map (
            O => \N__31731\,
            I => \N__31726\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__31726\,
            I => \N__31723\
        );

    \I__6977\ : Odrv4
    port map (
            O => \N__31723\,
            I => \b2v_inst5.un2_count_1_cry_8_THRU_CO\
        );

    \I__6976\ : CascadeMux
    port map (
            O => \N__31720\,
            I => \b2v_inst5.un2_count_1_axb_9_cascade_\
        );

    \I__6975\ : InMux
    port map (
            O => \N__31717\,
            I => \N__31711\
        );

    \I__6974\ : InMux
    port map (
            O => \N__31716\,
            I => \N__31711\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__31711\,
            I => \b2v_inst5.count_0_9\
        );

    \I__6972\ : CascadeMux
    port map (
            O => \N__31708\,
            I => \b2v_inst5.count_rst_4_cascade_\
        );

    \I__6971\ : InMux
    port map (
            O => \N__31705\,
            I => \N__31701\
        );

    \I__6970\ : CascadeMux
    port map (
            O => \N__31704\,
            I => \N__31698\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__31701\,
            I => \N__31694\
        );

    \I__6968\ : InMux
    port map (
            O => \N__31698\,
            I => \N__31689\
        );

    \I__6967\ : InMux
    port map (
            O => \N__31697\,
            I => \N__31689\
        );

    \I__6966\ : Odrv4
    port map (
            O => \N__31694\,
            I => \b2v_inst5.countZ0Z_10\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__31689\,
            I => \b2v_inst5.countZ0Z_10\
        );

    \I__6964\ : CascadeMux
    port map (
            O => \N__31684\,
            I => \b2v_inst5.countZ0Z_10_cascade_\
        );

    \I__6963\ : InMux
    port map (
            O => \N__31681\,
            I => \N__31675\
        );

    \I__6962\ : InMux
    port map (
            O => \N__31680\,
            I => \N__31675\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__31675\,
            I => \N__31672\
        );

    \I__6960\ : Span4Mux_s0_h
    port map (
            O => \N__31672\,
            I => \N__31669\
        );

    \I__6959\ : Odrv4
    port map (
            O => \N__31669\,
            I => \b2v_inst5.un2_count_1_cry_9_THRU_CO\
        );

    \I__6958\ : InMux
    port map (
            O => \N__31666\,
            I => \N__31663\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__31663\,
            I => \b2v_inst5.count_0_10\
        );

    \I__6956\ : CascadeMux
    port map (
            O => \N__31660\,
            I => \b2v_inst6.countZ0Z_8_cascade_\
        );

    \I__6955\ : InMux
    port map (
            O => \N__31657\,
            I => \N__31651\
        );

    \I__6954\ : InMux
    port map (
            O => \N__31656\,
            I => \N__31651\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__31651\,
            I => \N__31648\
        );

    \I__6952\ : Odrv12
    port map (
            O => \N__31648\,
            I => \b2v_inst6.un2_count_1_cry_7_THRU_CO\
        );

    \I__6951\ : InMux
    port map (
            O => \N__31645\,
            I => \N__31642\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__31642\,
            I => \b2v_inst6.count_3_8\
        );

    \I__6949\ : CascadeMux
    port map (
            O => \N__31639\,
            I => \N__31636\
        );

    \I__6948\ : InMux
    port map (
            O => \N__31636\,
            I => \N__31630\
        );

    \I__6947\ : InMux
    port map (
            O => \N__31635\,
            I => \N__31625\
        );

    \I__6946\ : InMux
    port map (
            O => \N__31634\,
            I => \N__31625\
        );

    \I__6945\ : InMux
    port map (
            O => \N__31633\,
            I => \N__31622\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__31630\,
            I => \b2v_inst6.countZ0Z_9\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__31625\,
            I => \b2v_inst6.countZ0Z_9\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__31622\,
            I => \b2v_inst6.countZ0Z_9\
        );

    \I__6941\ : InMux
    port map (
            O => \N__31615\,
            I => \N__31612\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__31612\,
            I => \N__31608\
        );

    \I__6939\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31605\
        );

    \I__6938\ : Odrv4
    port map (
            O => \N__31608\,
            I => \b2v_inst6.un2_count_1_cry_8_THRU_CO\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__31605\,
            I => \b2v_inst6.un2_count_1_cry_8_THRU_CO\
        );

    \I__6936\ : InMux
    port map (
            O => \N__31600\,
            I => \N__31597\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__31597\,
            I => \N__31594\
        );

    \I__6934\ : Odrv4
    port map (
            O => \N__31594\,
            I => \b2v_inst6.count_3_9\
        );

    \I__6933\ : CascadeMux
    port map (
            O => \N__31591\,
            I => \b2v_inst36.N_2928_i_cascade_\
        );

    \I__6932\ : InMux
    port map (
            O => \N__31588\,
            I => \N__31585\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__31585\,
            I => \b2v_inst36.count_1_13\
        );

    \I__6930\ : InMux
    port map (
            O => \N__31582\,
            I => \N__31576\
        );

    \I__6929\ : InMux
    port map (
            O => \N__31581\,
            I => \N__31576\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__31576\,
            I => \N__31573\
        );

    \I__6927\ : Odrv4
    port map (
            O => \N__31573\,
            I => \b2v_inst36.un2_count_1_cry_12_c_RNIS7LZ0Z1\
        );

    \I__6926\ : CascadeMux
    port map (
            O => \N__31570\,
            I => \N__31566\
        );

    \I__6925\ : InMux
    port map (
            O => \N__31569\,
            I => \N__31563\
        );

    \I__6924\ : InMux
    port map (
            O => \N__31566\,
            I => \N__31560\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__31563\,
            I => \N__31557\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__31560\,
            I => \b2v_inst36.countZ0Z_13\
        );

    \I__6921\ : Odrv4
    port map (
            O => \N__31557\,
            I => \b2v_inst36.countZ0Z_13\
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__31552\,
            I => \N__31549\
        );

    \I__6919\ : InMux
    port map (
            O => \N__31549\,
            I => \N__31545\
        );

    \I__6918\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31542\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__31545\,
            I => \N__31539\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__31542\,
            I => \b2v_inst36.countZ0Z_9\
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__31539\,
            I => \b2v_inst36.countZ0Z_9\
        );

    \I__6914\ : CascadeMux
    port map (
            O => \N__31534\,
            I => \N__31531\
        );

    \I__6913\ : InMux
    port map (
            O => \N__31531\,
            I => \N__31525\
        );

    \I__6912\ : InMux
    port map (
            O => \N__31530\,
            I => \N__31525\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__31525\,
            I => \N__31522\
        );

    \I__6910\ : Span4Mux_s1_h
    port map (
            O => \N__31522\,
            I => \N__31519\
        );

    \I__6909\ : Odrv4
    port map (
            O => \N__31519\,
            I => \b2v_inst36.un2_count_1_cry_8_c_RNIH8IZ0Z8\
        );

    \I__6908\ : InMux
    port map (
            O => \N__31516\,
            I => \N__31513\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__31513\,
            I => \b2v_inst36.count_1_9\
        );

    \I__6906\ : CascadeMux
    port map (
            O => \N__31510\,
            I => \b2v_inst6.count_rst_8_cascade_\
        );

    \I__6905\ : InMux
    port map (
            O => \N__31507\,
            I => \N__31501\
        );

    \I__6904\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31501\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__31501\,
            I => \b2v_inst6.count_rst_9\
        );

    \I__6902\ : InMux
    port map (
            O => \N__31498\,
            I => \N__31495\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__31495\,
            I => \N__31492\
        );

    \I__6900\ : Odrv4
    port map (
            O => \N__31492\,
            I => \b2v_inst6.count_3_10\
        );

    \I__6899\ : InMux
    port map (
            O => \N__31489\,
            I => \N__31485\
        );

    \I__6898\ : CascadeMux
    port map (
            O => \N__31488\,
            I => \N__31481\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__31485\,
            I => \N__31478\
        );

    \I__6896\ : InMux
    port map (
            O => \N__31484\,
            I => \N__31475\
        );

    \I__6895\ : InMux
    port map (
            O => \N__31481\,
            I => \N__31472\
        );

    \I__6894\ : Span4Mux_s2_h
    port map (
            O => \N__31478\,
            I => \N__31469\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__31475\,
            I => \N__31466\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__31472\,
            I => \b2v_inst6.countZ0Z_11\
        );

    \I__6891\ : Odrv4
    port map (
            O => \N__31469\,
            I => \b2v_inst6.countZ0Z_11\
        );

    \I__6890\ : Odrv12
    port map (
            O => \N__31466\,
            I => \b2v_inst6.countZ0Z_11\
        );

    \I__6889\ : CascadeMux
    port map (
            O => \N__31459\,
            I => \b2v_inst6.count_rst_6_cascade_\
        );

    \I__6888\ : CascadeMux
    port map (
            O => \N__31456\,
            I => \N__31451\
        );

    \I__6887\ : InMux
    port map (
            O => \N__31455\,
            I => \N__31448\
        );

    \I__6886\ : InMux
    port map (
            O => \N__31454\,
            I => \N__31443\
        );

    \I__6885\ : InMux
    port map (
            O => \N__31451\,
            I => \N__31443\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__31448\,
            I => \N__31440\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__31443\,
            I => \b2v_inst6.countZ0Z_7\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__31440\,
            I => \b2v_inst6.countZ0Z_7\
        );

    \I__6881\ : InMux
    port map (
            O => \N__31435\,
            I => \N__31429\
        );

    \I__6880\ : InMux
    port map (
            O => \N__31434\,
            I => \N__31429\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__31429\,
            I => \N__31426\
        );

    \I__6878\ : Odrv4
    port map (
            O => \N__31426\,
            I => \b2v_inst6.un2_count_1_cry_6_THRU_CO\
        );

    \I__6877\ : CascadeMux
    port map (
            O => \N__31423\,
            I => \b2v_inst6.countZ0Z_7_cascade_\
        );

    \I__6876\ : InMux
    port map (
            O => \N__31420\,
            I => \N__31417\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__31417\,
            I => \b2v_inst6.count_3_7\
        );

    \I__6874\ : CascadeMux
    port map (
            O => \N__31414\,
            I => \b2v_inst6.count_rst_7_cascade_\
        );

    \I__6873\ : CascadeMux
    port map (
            O => \N__31411\,
            I => \N__31407\
        );

    \I__6872\ : InMux
    port map (
            O => \N__31410\,
            I => \N__31403\
        );

    \I__6871\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31398\
        );

    \I__6870\ : InMux
    port map (
            O => \N__31406\,
            I => \N__31398\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__31403\,
            I => \N__31395\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__31398\,
            I => \b2v_inst6.countZ0Z_8\
        );

    \I__6867\ : Odrv4
    port map (
            O => \N__31395\,
            I => \b2v_inst6.countZ0Z_8\
        );

    \I__6866\ : InMux
    port map (
            O => \N__31390\,
            I => \b2v_inst6.un2_count_1_cry_11\
        );

    \I__6865\ : InMux
    port map (
            O => \N__31387\,
            I => \b2v_inst6.un2_count_1_cry_12\
        );

    \I__6864\ : InMux
    port map (
            O => \N__31384\,
            I => \b2v_inst6.un2_count_1_cry_13\
        );

    \I__6863\ : InMux
    port map (
            O => \N__31381\,
            I => \b2v_inst6.un2_count_1_cry_14\
        );

    \I__6862\ : CascadeMux
    port map (
            O => \N__31378\,
            I => \N__31375\
        );

    \I__6861\ : InMux
    port map (
            O => \N__31375\,
            I => \N__31372\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__31372\,
            I => \N__31368\
        );

    \I__6859\ : InMux
    port map (
            O => \N__31371\,
            I => \N__31365\
        );

    \I__6858\ : Span4Mux_s3_v
    port map (
            O => \N__31368\,
            I => \N__31362\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__31365\,
            I => \N__31359\
        );

    \I__6856\ : Odrv4
    port map (
            O => \N__31362\,
            I => \b2v_inst6.un2_count_1_cry_4_THRU_CO\
        );

    \I__6855\ : Odrv12
    port map (
            O => \N__31359\,
            I => \b2v_inst6.un2_count_1_cry_4_THRU_CO\
        );

    \I__6854\ : CascadeMux
    port map (
            O => \N__31354\,
            I => \b2v_inst6.count_rst_4_cascade_\
        );

    \I__6853\ : InMux
    port map (
            O => \N__31351\,
            I => \N__31348\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__31348\,
            I => \N__31345\
        );

    \I__6851\ : Span4Mux_s2_h
    port map (
            O => \N__31345\,
            I => \N__31342\
        );

    \I__6850\ : Odrv4
    port map (
            O => \N__31342\,
            I => \b2v_inst6.count_3_5\
        );

    \I__6849\ : CascadeMux
    port map (
            O => \N__31339\,
            I => \b2v_inst6.count_rst_2_cascade_\
        );

    \I__6848\ : InMux
    port map (
            O => \N__31336\,
            I => \b2v_inst6.un2_count_1_cry_2\
        );

    \I__6847\ : InMux
    port map (
            O => \N__31333\,
            I => \N__31327\
        );

    \I__6846\ : InMux
    port map (
            O => \N__31332\,
            I => \N__31327\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__31327\,
            I => \N__31324\
        );

    \I__6844\ : Span4Mux_h
    port map (
            O => \N__31324\,
            I => \N__31321\
        );

    \I__6843\ : Odrv4
    port map (
            O => \N__31321\,
            I => \b2v_inst6.un2_count_1_cry_3_THRU_CO\
        );

    \I__6842\ : InMux
    port map (
            O => \N__31318\,
            I => \b2v_inst6.un2_count_1_cry_3\
        );

    \I__6841\ : InMux
    port map (
            O => \N__31315\,
            I => \b2v_inst6.un2_count_1_cry_4\
        );

    \I__6840\ : InMux
    port map (
            O => \N__31312\,
            I => \b2v_inst6.un2_count_1_cry_5\
        );

    \I__6839\ : InMux
    port map (
            O => \N__31309\,
            I => \b2v_inst6.un2_count_1_cry_6\
        );

    \I__6838\ : InMux
    port map (
            O => \N__31306\,
            I => \b2v_inst6.un2_count_1_cry_7\
        );

    \I__6837\ : InMux
    port map (
            O => \N__31303\,
            I => \bfn_11_14_0_\
        );

    \I__6836\ : InMux
    port map (
            O => \N__31300\,
            I => \b2v_inst6.un2_count_1_cry_9\
        );

    \I__6835\ : InMux
    port map (
            O => \N__31297\,
            I => \N__31291\
        );

    \I__6834\ : InMux
    port map (
            O => \N__31296\,
            I => \N__31291\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__31291\,
            I => \N__31288\
        );

    \I__6832\ : Odrv4
    port map (
            O => \N__31288\,
            I => \b2v_inst6.un2_count_1_cry_10_THRU_CO\
        );

    \I__6831\ : InMux
    port map (
            O => \N__31285\,
            I => \b2v_inst6.un2_count_1_cry_10\
        );

    \I__6830\ : InMux
    port map (
            O => \N__31282\,
            I => \bfn_11_12_0_\
        );

    \I__6829\ : InMux
    port map (
            O => \N__31279\,
            I => \b2v_inst20.counter_1_cry_25\
        );

    \I__6828\ : InMux
    port map (
            O => \N__31276\,
            I => \b2v_inst20.counter_1_cry_26\
        );

    \I__6827\ : InMux
    port map (
            O => \N__31273\,
            I => \b2v_inst20.counter_1_cry_27\
        );

    \I__6826\ : InMux
    port map (
            O => \N__31270\,
            I => \b2v_inst20.counter_1_cry_28\
        );

    \I__6825\ : InMux
    port map (
            O => \N__31267\,
            I => \b2v_inst20.counter_1_cry_29\
        );

    \I__6824\ : InMux
    port map (
            O => \N__31264\,
            I => \b2v_inst20.counter_1_cry_30\
        );

    \I__6823\ : InMux
    port map (
            O => \N__31261\,
            I => \b2v_inst6.un2_count_1_cry_1\
        );

    \I__6822\ : InMux
    port map (
            O => \N__31258\,
            I => \b2v_inst20.counter_1_cry_15\
        );

    \I__6821\ : InMux
    port map (
            O => \N__31255\,
            I => \bfn_11_11_0_\
        );

    \I__6820\ : InMux
    port map (
            O => \N__31252\,
            I => \b2v_inst20.counter_1_cry_17\
        );

    \I__6819\ : InMux
    port map (
            O => \N__31249\,
            I => \b2v_inst20.counter_1_cry_18\
        );

    \I__6818\ : InMux
    port map (
            O => \N__31246\,
            I => \b2v_inst20.counter_1_cry_19\
        );

    \I__6817\ : InMux
    port map (
            O => \N__31243\,
            I => \b2v_inst20.counter_1_cry_20\
        );

    \I__6816\ : InMux
    port map (
            O => \N__31240\,
            I => \b2v_inst20.counter_1_cry_21\
        );

    \I__6815\ : InMux
    port map (
            O => \N__31237\,
            I => \b2v_inst20.counter_1_cry_22\
        );

    \I__6814\ : InMux
    port map (
            O => \N__31234\,
            I => \b2v_inst20.counter_1_cry_23\
        );

    \I__6813\ : InMux
    port map (
            O => \N__31231\,
            I => \N__31228\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__31228\,
            I => \N__31224\
        );

    \I__6811\ : InMux
    port map (
            O => \N__31227\,
            I => \N__31221\
        );

    \I__6810\ : Span4Mux_h
    port map (
            O => \N__31224\,
            I => \N__31218\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__31221\,
            I => \b2v_inst20.counterZ0Z_7\
        );

    \I__6808\ : Odrv4
    port map (
            O => \N__31218\,
            I => \b2v_inst20.counterZ0Z_7\
        );

    \I__6807\ : InMux
    port map (
            O => \N__31213\,
            I => \b2v_inst20.counter_1_cry_6\
        );

    \I__6806\ : InMux
    port map (
            O => \N__31210\,
            I => \b2v_inst20.counter_1_cry_7\
        );

    \I__6805\ : InMux
    port map (
            O => \N__31207\,
            I => \bfn_11_10_0_\
        );

    \I__6804\ : InMux
    port map (
            O => \N__31204\,
            I => \b2v_inst20.counter_1_cry_9\
        );

    \I__6803\ : InMux
    port map (
            O => \N__31201\,
            I => \b2v_inst20.counter_1_cry_10\
        );

    \I__6802\ : InMux
    port map (
            O => \N__31198\,
            I => \b2v_inst20.counter_1_cry_11\
        );

    \I__6801\ : InMux
    port map (
            O => \N__31195\,
            I => \b2v_inst20.counter_1_cry_12\
        );

    \I__6800\ : InMux
    port map (
            O => \N__31192\,
            I => \b2v_inst20.counter_1_cry_13\
        );

    \I__6799\ : InMux
    port map (
            O => \N__31189\,
            I => \b2v_inst20.counter_1_cry_14\
        );

    \I__6798\ : InMux
    port map (
            O => \N__31186\,
            I => \N__31183\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__31183\,
            I => \N__31179\
        );

    \I__6796\ : InMux
    port map (
            O => \N__31182\,
            I => \N__31176\
        );

    \I__6795\ : Odrv4
    port map (
            O => \N__31179\,
            I => \b2v_inst5.countZ0Z_15\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__31176\,
            I => \b2v_inst5.countZ0Z_15\
        );

    \I__6793\ : InMux
    port map (
            O => \N__31171\,
            I => \b2v_inst5.un2_count_1_cry_14\
        );

    \I__6792\ : InMux
    port map (
            O => \N__31168\,
            I => \N__31164\
        );

    \I__6791\ : InMux
    port map (
            O => \N__31167\,
            I => \N__31161\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__31164\,
            I => \N__31158\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__31161\,
            I => \b2v_inst5.count_rst\
        );

    \I__6788\ : Odrv12
    port map (
            O => \N__31158\,
            I => \b2v_inst5.count_rst\
        );

    \I__6787\ : InMux
    port map (
            O => \N__31153\,
            I => \N__31150\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__31150\,
            I => \N__31147\
        );

    \I__6785\ : Odrv12
    port map (
            O => \N__31147\,
            I => \b2v_inst5.count_0_15\
        );

    \I__6784\ : InMux
    port map (
            O => \N__31144\,
            I => \N__31141\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__31141\,
            I => \N__31137\
        );

    \I__6782\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31133\
        );

    \I__6781\ : Span4Mux_s2_h
    port map (
            O => \N__31137\,
            I => \N__31130\
        );

    \I__6780\ : InMux
    port map (
            O => \N__31136\,
            I => \N__31127\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__31133\,
            I => \b2v_inst20.counterZ0Z_1\
        );

    \I__6778\ : Odrv4
    port map (
            O => \N__31130\,
            I => \b2v_inst20.counterZ0Z_1\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__31127\,
            I => \b2v_inst20.counterZ0Z_1\
        );

    \I__6776\ : CascadeMux
    port map (
            O => \N__31120\,
            I => \N__31117\
        );

    \I__6775\ : InMux
    port map (
            O => \N__31117\,
            I => \N__31114\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__31114\,
            I => \N__31109\
        );

    \I__6773\ : InMux
    port map (
            O => \N__31113\,
            I => \N__31105\
        );

    \I__6772\ : InMux
    port map (
            O => \N__31112\,
            I => \N__31102\
        );

    \I__6771\ : Span4Mux_s2_h
    port map (
            O => \N__31109\,
            I => \N__31099\
        );

    \I__6770\ : InMux
    port map (
            O => \N__31108\,
            I => \N__31096\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__31105\,
            I => \b2v_inst20.counterZ0Z_0\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__31102\,
            I => \b2v_inst20.counterZ0Z_0\
        );

    \I__6767\ : Odrv4
    port map (
            O => \N__31099\,
            I => \b2v_inst20.counterZ0Z_0\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__31096\,
            I => \b2v_inst20.counterZ0Z_0\
        );

    \I__6765\ : InMux
    port map (
            O => \N__31087\,
            I => \N__31084\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__31084\,
            I => \N__31080\
        );

    \I__6763\ : InMux
    port map (
            O => \N__31083\,
            I => \N__31076\
        );

    \I__6762\ : Span4Mux_s2_h
    port map (
            O => \N__31080\,
            I => \N__31073\
        );

    \I__6761\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31070\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__31076\,
            I => \b2v_inst20.counterZ0Z_2\
        );

    \I__6759\ : Odrv4
    port map (
            O => \N__31073\,
            I => \b2v_inst20.counterZ0Z_2\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__31070\,
            I => \b2v_inst20.counterZ0Z_2\
        );

    \I__6757\ : InMux
    port map (
            O => \N__31063\,
            I => \N__31060\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__31060\,
            I => \N__31057\
        );

    \I__6755\ : Span4Mux_h
    port map (
            O => \N__31057\,
            I => \N__31054\
        );

    \I__6754\ : Odrv4
    port map (
            O => \N__31054\,
            I => \b2v_inst20.counter_1_cry_1_THRU_CO\
        );

    \I__6753\ : InMux
    port map (
            O => \N__31051\,
            I => \b2v_inst20.counter_1_cry_1\
        );

    \I__6752\ : InMux
    port map (
            O => \N__31048\,
            I => \N__31045\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__31045\,
            I => \N__31040\
        );

    \I__6750\ : CascadeMux
    port map (
            O => \N__31044\,
            I => \N__31037\
        );

    \I__6749\ : InMux
    port map (
            O => \N__31043\,
            I => \N__31034\
        );

    \I__6748\ : Span4Mux_s2_h
    port map (
            O => \N__31040\,
            I => \N__31031\
        );

    \I__6747\ : InMux
    port map (
            O => \N__31037\,
            I => \N__31028\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__31034\,
            I => \b2v_inst20.counterZ0Z_3\
        );

    \I__6745\ : Odrv4
    port map (
            O => \N__31031\,
            I => \b2v_inst20.counterZ0Z_3\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__31028\,
            I => \b2v_inst20.counterZ0Z_3\
        );

    \I__6743\ : InMux
    port map (
            O => \N__31021\,
            I => \N__31018\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__31018\,
            I => \N__31015\
        );

    \I__6741\ : Span4Mux_h
    port map (
            O => \N__31015\,
            I => \N__31012\
        );

    \I__6740\ : Odrv4
    port map (
            O => \N__31012\,
            I => \b2v_inst20.counter_1_cry_2_THRU_CO\
        );

    \I__6739\ : InMux
    port map (
            O => \N__31009\,
            I => \b2v_inst20.counter_1_cry_2\
        );

    \I__6738\ : InMux
    port map (
            O => \N__31006\,
            I => \N__31002\
        );

    \I__6737\ : InMux
    port map (
            O => \N__31005\,
            I => \N__30998\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__31002\,
            I => \N__30995\
        );

    \I__6735\ : InMux
    port map (
            O => \N__31001\,
            I => \N__30992\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__30998\,
            I => \b2v_inst20.counterZ0Z_4\
        );

    \I__6733\ : Odrv12
    port map (
            O => \N__30995\,
            I => \b2v_inst20.counterZ0Z_4\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__30992\,
            I => \b2v_inst20.counterZ0Z_4\
        );

    \I__6731\ : InMux
    port map (
            O => \N__30985\,
            I => \N__30982\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__30982\,
            I => \N__30979\
        );

    \I__6729\ : Odrv12
    port map (
            O => \N__30979\,
            I => \b2v_inst20.counter_1_cry_3_THRU_CO\
        );

    \I__6728\ : InMux
    port map (
            O => \N__30976\,
            I => \b2v_inst20.counter_1_cry_3\
        );

    \I__6727\ : InMux
    port map (
            O => \N__30973\,
            I => \N__30970\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__30970\,
            I => \N__30967\
        );

    \I__6725\ : Span4Mux_s3_h
    port map (
            O => \N__30967\,
            I => \N__30962\
        );

    \I__6724\ : InMux
    port map (
            O => \N__30966\,
            I => \N__30957\
        );

    \I__6723\ : InMux
    port map (
            O => \N__30965\,
            I => \N__30957\
        );

    \I__6722\ : Odrv4
    port map (
            O => \N__30962\,
            I => \b2v_inst20.counterZ0Z_5\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__30957\,
            I => \b2v_inst20.counterZ0Z_5\
        );

    \I__6720\ : InMux
    port map (
            O => \N__30952\,
            I => \N__30949\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__30949\,
            I => \N__30946\
        );

    \I__6718\ : Span4Mux_v
    port map (
            O => \N__30946\,
            I => \N__30943\
        );

    \I__6717\ : Odrv4
    port map (
            O => \N__30943\,
            I => \b2v_inst20.counter_1_cry_4_THRU_CO\
        );

    \I__6716\ : InMux
    port map (
            O => \N__30940\,
            I => \b2v_inst20.counter_1_cry_4\
        );

    \I__6715\ : InMux
    port map (
            O => \N__30937\,
            I => \N__30934\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__30934\,
            I => \N__30930\
        );

    \I__6713\ : CascadeMux
    port map (
            O => \N__30933\,
            I => \N__30926\
        );

    \I__6712\ : Span4Mux_v
    port map (
            O => \N__30930\,
            I => \N__30923\
        );

    \I__6711\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30918\
        );

    \I__6710\ : InMux
    port map (
            O => \N__30926\,
            I => \N__30918\
        );

    \I__6709\ : Odrv4
    port map (
            O => \N__30923\,
            I => \b2v_inst20.counterZ0Z_6\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__30918\,
            I => \b2v_inst20.counterZ0Z_6\
        );

    \I__6707\ : InMux
    port map (
            O => \N__30913\,
            I => \N__30910\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__30910\,
            I => \N__30907\
        );

    \I__6705\ : Span4Mux_v
    port map (
            O => \N__30907\,
            I => \N__30904\
        );

    \I__6704\ : Span4Mux_h
    port map (
            O => \N__30904\,
            I => \N__30901\
        );

    \I__6703\ : Odrv4
    port map (
            O => \N__30901\,
            I => \b2v_inst20.counter_1_cry_5_THRU_CO\
        );

    \I__6702\ : InMux
    port map (
            O => \N__30898\,
            I => \b2v_inst20.counter_1_cry_5\
        );

    \I__6701\ : CascadeMux
    port map (
            O => \N__30895\,
            I => \N__30892\
        );

    \I__6700\ : InMux
    port map (
            O => \N__30892\,
            I => \N__30888\
        );

    \I__6699\ : InMux
    port map (
            O => \N__30891\,
            I => \N__30885\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__30888\,
            I => \N__30882\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__30885\,
            I => \N__30879\
        );

    \I__6696\ : Span4Mux_v
    port map (
            O => \N__30882\,
            I => \N__30876\
        );

    \I__6695\ : Span4Mux_s2_h
    port map (
            O => \N__30879\,
            I => \N__30873\
        );

    \I__6694\ : Odrv4
    port map (
            O => \N__30876\,
            I => \b2v_inst5.countZ0Z_7\
        );

    \I__6693\ : Odrv4
    port map (
            O => \N__30873\,
            I => \b2v_inst5.countZ0Z_7\
        );

    \I__6692\ : InMux
    port map (
            O => \N__30868\,
            I => \N__30864\
        );

    \I__6691\ : InMux
    port map (
            O => \N__30867\,
            I => \N__30861\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__30864\,
            I => \N__30858\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__30861\,
            I => \N__30855\
        );

    \I__6688\ : Span4Mux_h
    port map (
            O => \N__30858\,
            I => \N__30852\
        );

    \I__6687\ : Odrv12
    port map (
            O => \N__30855\,
            I => \b2v_inst5.count_rst_7\
        );

    \I__6686\ : Odrv4
    port map (
            O => \N__30852\,
            I => \b2v_inst5.count_rst_7\
        );

    \I__6685\ : InMux
    port map (
            O => \N__30847\,
            I => \b2v_inst5.un2_count_1_cry_6\
        );

    \I__6684\ : InMux
    port map (
            O => \N__30844\,
            I => \b2v_inst5.un2_count_1_cry_7\
        );

    \I__6683\ : InMux
    port map (
            O => \N__30841\,
            I => \bfn_11_8_0_\
        );

    \I__6682\ : InMux
    port map (
            O => \N__30838\,
            I => \b2v_inst5.un2_count_1_cry_9\
        );

    \I__6681\ : InMux
    port map (
            O => \N__30835\,
            I => \b2v_inst5.un2_count_1_cry_10\
        );

    \I__6680\ : CascadeMux
    port map (
            O => \N__30832\,
            I => \N__30829\
        );

    \I__6679\ : InMux
    port map (
            O => \N__30829\,
            I => \N__30826\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__30826\,
            I => \N__30823\
        );

    \I__6677\ : Odrv4
    port map (
            O => \N__30823\,
            I => \b2v_inst5.un2_count_1_axb_12\
        );

    \I__6676\ : InMux
    port map (
            O => \N__30820\,
            I => \N__30811\
        );

    \I__6675\ : InMux
    port map (
            O => \N__30819\,
            I => \N__30811\
        );

    \I__6674\ : InMux
    port map (
            O => \N__30818\,
            I => \N__30811\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__30811\,
            I => \N__30808\
        );

    \I__6672\ : Odrv4
    port map (
            O => \N__30808\,
            I => \b2v_inst5.count_rst_2\
        );

    \I__6671\ : InMux
    port map (
            O => \N__30805\,
            I => \b2v_inst5.un2_count_1_cry_11\
        );

    \I__6670\ : InMux
    port map (
            O => \N__30802\,
            I => \b2v_inst5.un2_count_1_cry_12\
        );

    \I__6669\ : CascadeMux
    port map (
            O => \N__30799\,
            I => \N__30796\
        );

    \I__6668\ : InMux
    port map (
            O => \N__30796\,
            I => \N__30793\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__30793\,
            I => \N__30789\
        );

    \I__6666\ : InMux
    port map (
            O => \N__30792\,
            I => \N__30786\
        );

    \I__6665\ : Span4Mux_v
    port map (
            O => \N__30789\,
            I => \N__30783\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__30786\,
            I => \N__30780\
        );

    \I__6663\ : Odrv4
    port map (
            O => \N__30783\,
            I => \b2v_inst5.countZ0Z_14\
        );

    \I__6662\ : Odrv12
    port map (
            O => \N__30780\,
            I => \b2v_inst5.countZ0Z_14\
        );

    \I__6661\ : InMux
    port map (
            O => \N__30775\,
            I => \N__30771\
        );

    \I__6660\ : InMux
    port map (
            O => \N__30774\,
            I => \N__30768\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__30771\,
            I => \N__30765\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__30768\,
            I => \N__30762\
        );

    \I__6657\ : Odrv12
    port map (
            O => \N__30765\,
            I => \b2v_inst5.count_rst_0\
        );

    \I__6656\ : Odrv4
    port map (
            O => \N__30762\,
            I => \b2v_inst5.count_rst_0\
        );

    \I__6655\ : InMux
    port map (
            O => \N__30757\,
            I => \b2v_inst5.un2_count_1_cry_13\
        );

    \I__6654\ : InMux
    port map (
            O => \N__30754\,
            I => \N__30748\
        );

    \I__6653\ : InMux
    port map (
            O => \N__30753\,
            I => \N__30748\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__30748\,
            I => \b2v_inst5.count_0_5\
        );

    \I__6651\ : InMux
    port map (
            O => \N__30745\,
            I => \N__30741\
        );

    \I__6650\ : InMux
    port map (
            O => \N__30744\,
            I => \N__30738\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__30741\,
            I => \N__30735\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__30738\,
            I => \N__30732\
        );

    \I__6647\ : Span4Mux_v
    port map (
            O => \N__30735\,
            I => \N__30729\
        );

    \I__6646\ : Odrv4
    port map (
            O => \N__30732\,
            I => \b2v_inst5.count_0_6\
        );

    \I__6645\ : Odrv4
    port map (
            O => \N__30729\,
            I => \b2v_inst5.count_0_6\
        );

    \I__6644\ : InMux
    port map (
            O => \N__30724\,
            I => \N__30721\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__30721\,
            I => \b2v_inst5.count_1_i_a2_2_0\
        );

    \I__6642\ : InMux
    port map (
            O => \N__30718\,
            I => \b2v_inst5.un2_count_1_cry_1\
        );

    \I__6641\ : InMux
    port map (
            O => \N__30715\,
            I => \b2v_inst5.un2_count_1_cry_2\
        );

    \I__6640\ : InMux
    port map (
            O => \N__30712\,
            I => \b2v_inst5.un2_count_1_cry_3\
        );

    \I__6639\ : InMux
    port map (
            O => \N__30709\,
            I => \N__30706\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__30706\,
            I => \b2v_inst5.un2_count_1_axb_5\
        );

    \I__6637\ : InMux
    port map (
            O => \N__30703\,
            I => \N__30694\
        );

    \I__6636\ : InMux
    port map (
            O => \N__30702\,
            I => \N__30694\
        );

    \I__6635\ : InMux
    port map (
            O => \N__30701\,
            I => \N__30694\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__30694\,
            I => \b2v_inst5.count_rst_9\
        );

    \I__6633\ : InMux
    port map (
            O => \N__30691\,
            I => \b2v_inst5.un2_count_1_cry_4\
        );

    \I__6632\ : InMux
    port map (
            O => \N__30688\,
            I => \N__30685\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__30685\,
            I => \N__30682\
        );

    \I__6630\ : Span4Mux_s2_h
    port map (
            O => \N__30682\,
            I => \N__30679\
        );

    \I__6629\ : Odrv4
    port map (
            O => \N__30679\,
            I => \b2v_inst5.un2_count_1_axb_6\
        );

    \I__6628\ : InMux
    port map (
            O => \N__30676\,
            I => \N__30673\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__30673\,
            I => \N__30670\
        );

    \I__6626\ : Span4Mux_v
    port map (
            O => \N__30670\,
            I => \N__30666\
        );

    \I__6625\ : InMux
    port map (
            O => \N__30669\,
            I => \N__30662\
        );

    \I__6624\ : Sp12to4
    port map (
            O => \N__30666\,
            I => \N__30659\
        );

    \I__6623\ : InMux
    port map (
            O => \N__30665\,
            I => \N__30656\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__30662\,
            I => \N__30653\
        );

    \I__6621\ : Odrv12
    port map (
            O => \N__30659\,
            I => \b2v_inst5.count_rst_8\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__30656\,
            I => \b2v_inst5.count_rst_8\
        );

    \I__6619\ : Odrv4
    port map (
            O => \N__30653\,
            I => \b2v_inst5.count_rst_8\
        );

    \I__6618\ : InMux
    port map (
            O => \N__30646\,
            I => \b2v_inst5.un2_count_1_cry_5\
        );

    \I__6617\ : CascadeMux
    port map (
            O => \N__30643\,
            I => \N__30640\
        );

    \I__6616\ : InMux
    port map (
            O => \N__30640\,
            I => \N__30634\
        );

    \I__6615\ : CEMux
    port map (
            O => \N__30639\,
            I => \N__30634\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__30634\,
            I => \N__30619\
        );

    \I__6613\ : InMux
    port map (
            O => \N__30633\,
            I => \N__30610\
        );

    \I__6612\ : InMux
    port map (
            O => \N__30632\,
            I => \N__30610\
        );

    \I__6611\ : InMux
    port map (
            O => \N__30631\,
            I => \N__30610\
        );

    \I__6610\ : InMux
    port map (
            O => \N__30630\,
            I => \N__30610\
        );

    \I__6609\ : CEMux
    port map (
            O => \N__30629\,
            I => \N__30606\
        );

    \I__6608\ : CEMux
    port map (
            O => \N__30628\,
            I => \N__30599\
        );

    \I__6607\ : InMux
    port map (
            O => \N__30627\,
            I => \N__30589\
        );

    \I__6606\ : InMux
    port map (
            O => \N__30626\,
            I => \N__30589\
        );

    \I__6605\ : InMux
    port map (
            O => \N__30625\,
            I => \N__30589\
        );

    \I__6604\ : InMux
    port map (
            O => \N__30624\,
            I => \N__30589\
        );

    \I__6603\ : CEMux
    port map (
            O => \N__30623\,
            I => \N__30586\
        );

    \I__6602\ : CEMux
    port map (
            O => \N__30622\,
            I => \N__30583\
        );

    \I__6601\ : Span4Mux_s2_v
    port map (
            O => \N__30619\,
            I => \N__30578\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__30610\,
            I => \N__30578\
        );

    \I__6599\ : InMux
    port map (
            O => \N__30609\,
            I => \N__30575\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__30606\,
            I => \N__30568\
        );

    \I__6597\ : CEMux
    port map (
            O => \N__30605\,
            I => \N__30564\
        );

    \I__6596\ : CEMux
    port map (
            O => \N__30604\,
            I => \N__30561\
        );

    \I__6595\ : InMux
    port map (
            O => \N__30603\,
            I => \N__30556\
        );

    \I__6594\ : InMux
    port map (
            O => \N__30602\,
            I => \N__30556\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__30599\,
            I => \N__30553\
        );

    \I__6592\ : CEMux
    port map (
            O => \N__30598\,
            I => \N__30550\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__30589\,
            I => \N__30547\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__30586\,
            I => \N__30538\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__30583\,
            I => \N__30538\
        );

    \I__6588\ : Span4Mux_v
    port map (
            O => \N__30578\,
            I => \N__30538\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__30575\,
            I => \N__30538\
        );

    \I__6586\ : InMux
    port map (
            O => \N__30574\,
            I => \N__30529\
        );

    \I__6585\ : InMux
    port map (
            O => \N__30573\,
            I => \N__30529\
        );

    \I__6584\ : InMux
    port map (
            O => \N__30572\,
            I => \N__30529\
        );

    \I__6583\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30529\
        );

    \I__6582\ : Span4Mux_s2_h
    port map (
            O => \N__30568\,
            I => \N__30526\
        );

    \I__6581\ : InMux
    port map (
            O => \N__30567\,
            I => \N__30523\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__30564\,
            I => \N__30520\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__30561\,
            I => \N__30515\
        );

    \I__6578\ : LocalMux
    port map (
            O => \N__30556\,
            I => \N__30515\
        );

    \I__6577\ : Span4Mux_s1_h
    port map (
            O => \N__30553\,
            I => \N__30512\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__30550\,
            I => \N__30503\
        );

    \I__6575\ : Span4Mux_s2_v
    port map (
            O => \N__30547\,
            I => \N__30503\
        );

    \I__6574\ : Span4Mux_s2_v
    port map (
            O => \N__30538\,
            I => \N__30503\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__30529\,
            I => \N__30503\
        );

    \I__6572\ : Span4Mux_v
    port map (
            O => \N__30526\,
            I => \N__30498\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__30523\,
            I => \N__30498\
        );

    \I__6570\ : Span4Mux_h
    port map (
            O => \N__30520\,
            I => \N__30493\
        );

    \I__6569\ : Span4Mux_s1_h
    port map (
            O => \N__30515\,
            I => \N__30493\
        );

    \I__6568\ : Span4Mux_h
    port map (
            O => \N__30512\,
            I => \N__30490\
        );

    \I__6567\ : Span4Mux_h
    port map (
            O => \N__30503\,
            I => \N__30487\
        );

    \I__6566\ : Span4Mux_h
    port map (
            O => \N__30498\,
            I => \N__30482\
        );

    \I__6565\ : Span4Mux_h
    port map (
            O => \N__30493\,
            I => \N__30482\
        );

    \I__6564\ : Odrv4
    port map (
            O => \N__30490\,
            I => \b2v_inst16.count_en\
        );

    \I__6563\ : Odrv4
    port map (
            O => \N__30487\,
            I => \b2v_inst16.count_en\
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__30482\,
            I => \b2v_inst16.count_en\
        );

    \I__6561\ : InMux
    port map (
            O => \N__30475\,
            I => \N__30472\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__30472\,
            I => \N__30469\
        );

    \I__6559\ : Span4Mux_v
    port map (
            O => \N__30469\,
            I => \N__30466\
        );

    \I__6558\ : Odrv4
    port map (
            O => \N__30466\,
            I => \b2v_inst36.count_1_4\
        );

    \I__6557\ : InMux
    port map (
            O => \N__30463\,
            I => \N__30459\
        );

    \I__6556\ : InMux
    port map (
            O => \N__30462\,
            I => \N__30456\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__30459\,
            I => \N__30453\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__30456\,
            I => \N__30450\
        );

    \I__6553\ : Span4Mux_v
    port map (
            O => \N__30453\,
            I => \N__30447\
        );

    \I__6552\ : Odrv12
    port map (
            O => \N__30450\,
            I => \b2v_inst36.count_rst_10\
        );

    \I__6551\ : Odrv4
    port map (
            O => \N__30447\,
            I => \b2v_inst36.count_rst_10\
        );

    \I__6550\ : InMux
    port map (
            O => \N__30442\,
            I => \N__30438\
        );

    \I__6549\ : InMux
    port map (
            O => \N__30441\,
            I => \N__30435\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__30438\,
            I => \N__30432\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__30435\,
            I => \N__30427\
        );

    \I__6546\ : Span4Mux_h
    port map (
            O => \N__30432\,
            I => \N__30427\
        );

    \I__6545\ : Odrv4
    port map (
            O => \N__30427\,
            I => \b2v_inst36.countZ0Z_4\
        );

    \I__6544\ : CascadeMux
    port map (
            O => \N__30424\,
            I => \b2v_inst5.N_2906_i_cascade_\
        );

    \I__6543\ : CascadeMux
    port map (
            O => \N__30421\,
            I => \b2v_inst5.count_1_i_a2_1_0_cascade_\
        );

    \I__6542\ : InMux
    port map (
            O => \N__30418\,
            I => \N__30412\
        );

    \I__6541\ : InMux
    port map (
            O => \N__30417\,
            I => \N__30412\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__30412\,
            I => \b2v_inst5.count_0_12\
        );

    \I__6539\ : InMux
    port map (
            O => \N__30409\,
            I => \N__30406\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__30406\,
            I => \b2v_inst5.count_1_i_a2_0_0\
        );

    \I__6537\ : InMux
    port map (
            O => \N__30403\,
            I => \N__30399\
        );

    \I__6536\ : InMux
    port map (
            O => \N__30402\,
            I => \N__30396\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__30399\,
            I => \N__30393\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__30396\,
            I => \N__30390\
        );

    \I__6533\ : Sp12to4
    port map (
            O => \N__30393\,
            I => \N__30385\
        );

    \I__6532\ : Span4Mux_v
    port map (
            O => \N__30390\,
            I => \N__30382\
        );

    \I__6531\ : InMux
    port map (
            O => \N__30389\,
            I => \N__30379\
        );

    \I__6530\ : InMux
    port map (
            O => \N__30388\,
            I => \N__30376\
        );

    \I__6529\ : Span12Mux_v
    port map (
            O => \N__30385\,
            I => \N__30373\
        );

    \I__6528\ : Odrv4
    port map (
            O => \N__30382\,
            I => \b2v_inst36.curr_stateZ0Z_0\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__30379\,
            I => \b2v_inst36.curr_stateZ0Z_0\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__30376\,
            I => \b2v_inst36.curr_stateZ0Z_0\
        );

    \I__6525\ : Odrv12
    port map (
            O => \N__30373\,
            I => \b2v_inst36.curr_stateZ0Z_0\
        );

    \I__6524\ : InMux
    port map (
            O => \N__30364\,
            I => \N__30361\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__30361\,
            I => \b2v_inst36.curr_state_4_0\
        );

    \I__6522\ : InMux
    port map (
            O => \N__30358\,
            I => \N__30354\
        );

    \I__6521\ : CascadeMux
    port map (
            O => \N__30357\,
            I => \N__30350\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__30354\,
            I => \N__30346\
        );

    \I__6519\ : CascadeMux
    port map (
            O => \N__30353\,
            I => \N__30343\
        );

    \I__6518\ : InMux
    port map (
            O => \N__30350\,
            I => \N__30340\
        );

    \I__6517\ : CascadeMux
    port map (
            O => \N__30349\,
            I => \N__30337\
        );

    \I__6516\ : Span12Mux_v
    port map (
            O => \N__30346\,
            I => \N__30331\
        );

    \I__6515\ : InMux
    port map (
            O => \N__30343\,
            I => \N__30328\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__30340\,
            I => \N__30325\
        );

    \I__6513\ : InMux
    port map (
            O => \N__30337\,
            I => \N__30316\
        );

    \I__6512\ : InMux
    port map (
            O => \N__30336\,
            I => \N__30316\
        );

    \I__6511\ : InMux
    port map (
            O => \N__30335\,
            I => \N__30316\
        );

    \I__6510\ : InMux
    port map (
            O => \N__30334\,
            I => \N__30316\
        );

    \I__6509\ : Odrv12
    port map (
            O => \N__30331\,
            I => \b2v_inst36.curr_stateZ0Z_1\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__30328\,
            I => \b2v_inst36.curr_stateZ0Z_1\
        );

    \I__6507\ : Odrv4
    port map (
            O => \N__30325\,
            I => \b2v_inst36.curr_stateZ0Z_1\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__30316\,
            I => \b2v_inst36.curr_stateZ0Z_1\
        );

    \I__6505\ : CascadeMux
    port map (
            O => \N__30307\,
            I => \N__30303\
        );

    \I__6504\ : InMux
    port map (
            O => \N__30306\,
            I => \N__30295\
        );

    \I__6503\ : InMux
    port map (
            O => \N__30303\,
            I => \N__30282\
        );

    \I__6502\ : InMux
    port map (
            O => \N__30302\,
            I => \N__30282\
        );

    \I__6501\ : InMux
    port map (
            O => \N__30301\,
            I => \N__30282\
        );

    \I__6500\ : InMux
    port map (
            O => \N__30300\,
            I => \N__30282\
        );

    \I__6499\ : InMux
    port map (
            O => \N__30299\,
            I => \N__30282\
        );

    \I__6498\ : InMux
    port map (
            O => \N__30298\,
            I => \N__30282\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__30295\,
            I => \N__30279\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__30282\,
            I => \N__30276\
        );

    \I__6495\ : Span4Mux_v
    port map (
            O => \N__30279\,
            I => \N__30273\
        );

    \I__6494\ : Span4Mux_v
    port map (
            O => \N__30276\,
            I => \N__30270\
        );

    \I__6493\ : Span4Mux_h
    port map (
            O => \N__30273\,
            I => \N__30265\
        );

    \I__6492\ : Span4Mux_v
    port map (
            O => \N__30270\,
            I => \N__30265\
        );

    \I__6491\ : Span4Mux_v
    port map (
            O => \N__30265\,
            I => \N__30262\
        );

    \I__6490\ : Odrv4
    port map (
            O => \N__30262\,
            I => \V33DSW_OK_c\
        );

    \I__6489\ : InMux
    port map (
            O => \N__30259\,
            I => \N__30253\
        );

    \I__6488\ : InMux
    port map (
            O => \N__30258\,
            I => \N__30246\
        );

    \I__6487\ : InMux
    port map (
            O => \N__30257\,
            I => \N__30246\
        );

    \I__6486\ : InMux
    port map (
            O => \N__30256\,
            I => \N__30246\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__30253\,
            I => \N__30241\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__30246\,
            I => \N__30241\
        );

    \I__6483\ : Span4Mux_s3_h
    port map (
            O => \N__30241\,
            I => \N__30238\
        );

    \I__6482\ : Span4Mux_v
    port map (
            O => \N__30238\,
            I => \N__30235\
        );

    \I__6481\ : Span4Mux_h
    port map (
            O => \N__30235\,
            I => \N__30232\
        );

    \I__6480\ : Odrv4
    port map (
            O => \N__30232\,
            I => \b2v_inst36.N_2925_i\
        );

    \I__6479\ : InMux
    port map (
            O => \N__30229\,
            I => \N__30226\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__30226\,
            I => \N__30223\
        );

    \I__6477\ : IoSpan4Mux
    port map (
            O => \N__30223\,
            I => \N__30220\
        );

    \I__6476\ : IoSpan4Mux
    port map (
            O => \N__30220\,
            I => \N__30217\
        );

    \I__6475\ : Odrv4
    port map (
            O => \N__30217\,
            I => \b2v_inst5.count_0_14\
        );

    \I__6474\ : InMux
    port map (
            O => \N__30214\,
            I => \N__30211\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__30211\,
            I => \N__30208\
        );

    \I__6472\ : Span4Mux_v
    port map (
            O => \N__30208\,
            I => \N__30205\
        );

    \I__6471\ : Span4Mux_h
    port map (
            O => \N__30205\,
            I => \N__30202\
        );

    \I__6470\ : Odrv4
    port map (
            O => \N__30202\,
            I => \b2v_inst5.count_0_7\
        );

    \I__6469\ : InMux
    port map (
            O => \N__30199\,
            I => \N__30195\
        );

    \I__6468\ : InMux
    port map (
            O => \N__30198\,
            I => \N__30192\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__30195\,
            I => \N__30187\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__30192\,
            I => \N__30187\
        );

    \I__6465\ : Span4Mux_s2_h
    port map (
            O => \N__30187\,
            I => \N__30184\
        );

    \I__6464\ : Span4Mux_h
    port map (
            O => \N__30184\,
            I => \N__30181\
        );

    \I__6463\ : Span4Mux_h
    port map (
            O => \N__30181\,
            I => \N__30178\
        );

    \I__6462\ : Odrv4
    port map (
            O => \N__30178\,
            I => \b2v_inst16.countZ0Z_8\
        );

    \I__6461\ : InMux
    port map (
            O => \N__30175\,
            I => \N__30169\
        );

    \I__6460\ : InMux
    port map (
            O => \N__30174\,
            I => \N__30169\
        );

    \I__6459\ : LocalMux
    port map (
            O => \N__30169\,
            I => \N__30166\
        );

    \I__6458\ : Span4Mux_v
    port map (
            O => \N__30166\,
            I => \N__30163\
        );

    \I__6457\ : Sp12to4
    port map (
            O => \N__30163\,
            I => \N__30160\
        );

    \I__6456\ : Odrv12
    port map (
            O => \N__30160\,
            I => \b2v_inst16.count_rst_13\
        );

    \I__6455\ : InMux
    port map (
            O => \N__30157\,
            I => \N__30154\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__30154\,
            I => \b2v_inst16.count_4_8\
        );

    \I__6453\ : InMux
    port map (
            O => \N__30151\,
            I => \N__30147\
        );

    \I__6452\ : CascadeMux
    port map (
            O => \N__30150\,
            I => \N__30144\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__30147\,
            I => \N__30141\
        );

    \I__6450\ : InMux
    port map (
            O => \N__30144\,
            I => \N__30138\
        );

    \I__6449\ : Span4Mux_s1_v
    port map (
            O => \N__30141\,
            I => \N__30135\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__30138\,
            I => \N__30132\
        );

    \I__6447\ : Span4Mux_h
    port map (
            O => \N__30135\,
            I => \N__30129\
        );

    \I__6446\ : Span12Mux_s10_h
    port map (
            O => \N__30132\,
            I => \N__30126\
        );

    \I__6445\ : Span4Mux_h
    port map (
            O => \N__30129\,
            I => \N__30123\
        );

    \I__6444\ : Odrv12
    port map (
            O => \N__30126\,
            I => \b2v_inst16.countZ0Z_9\
        );

    \I__6443\ : Odrv4
    port map (
            O => \N__30123\,
            I => \b2v_inst16.countZ0Z_9\
        );

    \I__6442\ : InMux
    port map (
            O => \N__30118\,
            I => \N__30112\
        );

    \I__6441\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30112\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__30112\,
            I => \N__30109\
        );

    \I__6439\ : Span4Mux_s2_h
    port map (
            O => \N__30109\,
            I => \N__30106\
        );

    \I__6438\ : Span4Mux_h
    port map (
            O => \N__30106\,
            I => \N__30103\
        );

    \I__6437\ : Span4Mux_h
    port map (
            O => \N__30103\,
            I => \N__30100\
        );

    \I__6436\ : Odrv4
    port map (
            O => \N__30100\,
            I => \b2v_inst16.count_rst_14\
        );

    \I__6435\ : InMux
    port map (
            O => \N__30097\,
            I => \N__30094\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__30094\,
            I => \b2v_inst16.count_4_9\
        );

    \I__6433\ : InMux
    port map (
            O => \N__30091\,
            I => \N__30088\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__30088\,
            I => \N__30085\
        );

    \I__6431\ : Span4Mux_s1_v
    port map (
            O => \N__30085\,
            I => \N__30081\
        );

    \I__6430\ : InMux
    port map (
            O => \N__30084\,
            I => \N__30078\
        );

    \I__6429\ : Odrv4
    port map (
            O => \N__30081\,
            I => \b2v_inst36.un2_count_1_cry_10_THRU_CO\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__30078\,
            I => \b2v_inst36.un2_count_1_cry_10_THRU_CO\
        );

    \I__6427\ : CascadeMux
    port map (
            O => \N__30073\,
            I => \b2v_inst36.countZ0Z_11_cascade_\
        );

    \I__6426\ : InMux
    port map (
            O => \N__30070\,
            I => \N__30067\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__30067\,
            I => \b2v_inst36.count_1_11\
        );

    \I__6424\ : CascadeMux
    port map (
            O => \N__30064\,
            I => \N__30061\
        );

    \I__6423\ : InMux
    port map (
            O => \N__30061\,
            I => \N__30052\
        );

    \I__6422\ : InMux
    port map (
            O => \N__30060\,
            I => \N__30052\
        );

    \I__6421\ : InMux
    port map (
            O => \N__30059\,
            I => \N__30052\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__30052\,
            I => \N__30049\
        );

    \I__6419\ : Span4Mux_v
    port map (
            O => \N__30049\,
            I => \N__30046\
        );

    \I__6418\ : Odrv4
    port map (
            O => \N__30046\,
            I => \b2v_inst36.count_rst_8\
        );

    \I__6417\ : InMux
    port map (
            O => \N__30043\,
            I => \N__30037\
        );

    \I__6416\ : InMux
    port map (
            O => \N__30042\,
            I => \N__30037\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__30037\,
            I => \b2v_inst36.count_1_6\
        );

    \I__6414\ : InMux
    port map (
            O => \N__30034\,
            I => \N__30031\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__30031\,
            I => \N__30028\
        );

    \I__6412\ : Span4Mux_s2_v
    port map (
            O => \N__30028\,
            I => \N__30024\
        );

    \I__6411\ : InMux
    port map (
            O => \N__30027\,
            I => \N__30021\
        );

    \I__6410\ : Odrv4
    port map (
            O => \N__30024\,
            I => \b2v_inst36.countZ0Z_12\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__30021\,
            I => \b2v_inst36.countZ0Z_12\
        );

    \I__6408\ : CascadeMux
    port map (
            O => \N__30016\,
            I => \b2v_inst36.countZ0Z_6_cascade_\
        );

    \I__6407\ : InMux
    port map (
            O => \N__30013\,
            I => \N__30010\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__30010\,
            I => \b2v_inst36.un12_clk_100khz_9\
        );

    \I__6405\ : CascadeMux
    port map (
            O => \N__30007\,
            I => \b2v_inst36.curr_stateZ0Z_1_cascade_\
        );

    \I__6404\ : CascadeMux
    port map (
            O => \N__30004\,
            I => \b2v_inst36.curr_state_7_0_cascade_\
        );

    \I__6403\ : CascadeMux
    port map (
            O => \N__30001\,
            I => \b2v_inst36.curr_stateZ0Z_0_cascade_\
        );

    \I__6402\ : InMux
    port map (
            O => \N__29998\,
            I => \N__29995\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__29995\,
            I => \N__29992\
        );

    \I__6400\ : Span4Mux_h
    port map (
            O => \N__29992\,
            I => \N__29989\
        );

    \I__6399\ : Span4Mux_v
    port map (
            O => \N__29989\,
            I => \N__29986\
        );

    \I__6398\ : Odrv4
    port map (
            O => \N__29986\,
            I => \b2v_inst36.DSW_PWROK_0\
        );

    \I__6397\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29980\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__29980\,
            I => \b2v_inst36.curr_state_3_1\
        );

    \I__6395\ : InMux
    port map (
            O => \N__29977\,
            I => \N__29974\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__29974\,
            I => \b2v_inst36.curr_state_7_1\
        );

    \I__6393\ : CascadeMux
    port map (
            O => \N__29971\,
            I => \b2v_inst36.count_rst_12_cascade_\
        );

    \I__6392\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29964\
        );

    \I__6391\ : InMux
    port map (
            O => \N__29967\,
            I => \N__29960\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__29964\,
            I => \N__29957\
        );

    \I__6389\ : InMux
    port map (
            O => \N__29963\,
            I => \N__29954\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__29960\,
            I => \N__29951\
        );

    \I__6387\ : Odrv4
    port map (
            O => \N__29957\,
            I => \b2v_inst36.countZ0Z_2\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__29954\,
            I => \b2v_inst36.countZ0Z_2\
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__29951\,
            I => \b2v_inst36.countZ0Z_2\
        );

    \I__6384\ : CascadeMux
    port map (
            O => \N__29944\,
            I => \b2v_inst36.countZ0Z_2_cascade_\
        );

    \I__6383\ : CascadeMux
    port map (
            O => \N__29941\,
            I => \N__29937\
        );

    \I__6382\ : InMux
    port map (
            O => \N__29940\,
            I => \N__29934\
        );

    \I__6381\ : InMux
    port map (
            O => \N__29937\,
            I => \N__29931\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__29934\,
            I => \N__29926\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__29931\,
            I => \N__29926\
        );

    \I__6378\ : Span4Mux_s1_h
    port map (
            O => \N__29926\,
            I => \N__29923\
        );

    \I__6377\ : Odrv4
    port map (
            O => \N__29923\,
            I => \b2v_inst36.un2_count_1_cry_1_THRU_CO\
        );

    \I__6376\ : InMux
    port map (
            O => \N__29920\,
            I => \N__29917\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__29917\,
            I => \b2v_inst36.count_1_2\
        );

    \I__6374\ : CascadeMux
    port map (
            O => \N__29914\,
            I => \N__29910\
        );

    \I__6373\ : InMux
    port map (
            O => \N__29913\,
            I => \N__29906\
        );

    \I__6372\ : InMux
    port map (
            O => \N__29910\,
            I => \N__29900\
        );

    \I__6371\ : InMux
    port map (
            O => \N__29909\,
            I => \N__29900\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__29906\,
            I => \N__29897\
        );

    \I__6369\ : InMux
    port map (
            O => \N__29905\,
            I => \N__29894\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__29900\,
            I => \b2v_inst36.countZ0Z_3\
        );

    \I__6367\ : Odrv12
    port map (
            O => \N__29897\,
            I => \b2v_inst36.countZ0Z_3\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__29894\,
            I => \b2v_inst36.countZ0Z_3\
        );

    \I__6365\ : InMux
    port map (
            O => \N__29887\,
            I => \N__29884\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__29884\,
            I => \N__29880\
        );

    \I__6363\ : InMux
    port map (
            O => \N__29883\,
            I => \N__29877\
        );

    \I__6362\ : Odrv4
    port map (
            O => \N__29880\,
            I => \b2v_inst36.un2_count_1_cry_2_THRU_CO\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__29877\,
            I => \b2v_inst36.un2_count_1_cry_2_THRU_CO\
        );

    \I__6360\ : InMux
    port map (
            O => \N__29872\,
            I => \N__29869\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__29869\,
            I => \N__29866\
        );

    \I__6358\ : Odrv12
    port map (
            O => \N__29866\,
            I => \b2v_inst36.count_1_3\
        );

    \I__6357\ : InMux
    port map (
            O => \N__29863\,
            I => \N__29860\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__29860\,
            I => \N__29855\
        );

    \I__6355\ : InMux
    port map (
            O => \N__29859\,
            I => \N__29852\
        );

    \I__6354\ : InMux
    port map (
            O => \N__29858\,
            I => \N__29849\
        );

    \I__6353\ : Odrv12
    port map (
            O => \N__29855\,
            I => \b2v_inst36.countZ0Z_8\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__29852\,
            I => \b2v_inst36.countZ0Z_8\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__29849\,
            I => \b2v_inst36.countZ0Z_8\
        );

    \I__6350\ : InMux
    port map (
            O => \N__29842\,
            I => \N__29838\
        );

    \I__6349\ : CascadeMux
    port map (
            O => \N__29841\,
            I => \N__29835\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__29838\,
            I => \N__29831\
        );

    \I__6347\ : InMux
    port map (
            O => \N__29835\,
            I => \N__29828\
        );

    \I__6346\ : InMux
    port map (
            O => \N__29834\,
            I => \N__29825\
        );

    \I__6345\ : Odrv12
    port map (
            O => \N__29831\,
            I => \b2v_inst36.countZ0Z_10\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__29828\,
            I => \b2v_inst36.countZ0Z_10\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__29825\,
            I => \b2v_inst36.countZ0Z_10\
        );

    \I__6342\ : CascadeMux
    port map (
            O => \N__29818\,
            I => \N__29814\
        );

    \I__6341\ : CascadeMux
    port map (
            O => \N__29817\,
            I => \N__29811\
        );

    \I__6340\ : InMux
    port map (
            O => \N__29814\,
            I => \N__29807\
        );

    \I__6339\ : InMux
    port map (
            O => \N__29811\,
            I => \N__29804\
        );

    \I__6338\ : InMux
    port map (
            O => \N__29810\,
            I => \N__29801\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__29807\,
            I => \N__29798\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__29804\,
            I => \b2v_inst36.countZ0Z_1\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__29801\,
            I => \b2v_inst36.countZ0Z_1\
        );

    \I__6334\ : Odrv4
    port map (
            O => \N__29798\,
            I => \b2v_inst36.countZ0Z_1\
        );

    \I__6333\ : InMux
    port map (
            O => \N__29791\,
            I => \N__29788\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__29788\,
            I => \N__29785\
        );

    \I__6331\ : Span4Mux_v
    port map (
            O => \N__29785\,
            I => \N__29782\
        );

    \I__6330\ : Odrv4
    port map (
            O => \N__29782\,
            I => \b2v_inst36.un12_clk_100khz_11\
        );

    \I__6329\ : CascadeMux
    port map (
            O => \N__29779\,
            I => \b2v_inst36.un12_clk_100khz_10_cascade_\
        );

    \I__6328\ : InMux
    port map (
            O => \N__29776\,
            I => \N__29773\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__29773\,
            I => \b2v_inst36.un12_clk_100khz_8\
        );

    \I__6326\ : InMux
    port map (
            O => \N__29770\,
            I => \N__29767\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__29767\,
            I => \N__29764\
        );

    \I__6324\ : Span4Mux_s1_v
    port map (
            O => \N__29764\,
            I => \N__29761\
        );

    \I__6323\ : Odrv4
    port map (
            O => \N__29761\,
            I => \b2v_inst36.un2_count_1_axb_6\
        );

    \I__6322\ : InMux
    port map (
            O => \N__29758\,
            I => \N__29755\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__29755\,
            I => \N__29752\
        );

    \I__6320\ : Odrv4
    port map (
            O => \N__29752\,
            I => \b2v_inst36.count_rst_3\
        );

    \I__6319\ : CascadeMux
    port map (
            O => \N__29749\,
            I => \N__29746\
        );

    \I__6318\ : InMux
    port map (
            O => \N__29746\,
            I => \N__29742\
        );

    \I__6317\ : InMux
    port map (
            O => \N__29745\,
            I => \N__29738\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__29742\,
            I => \N__29735\
        );

    \I__6315\ : InMux
    port map (
            O => \N__29741\,
            I => \N__29732\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__29738\,
            I => \N__29729\
        );

    \I__6313\ : Odrv4
    port map (
            O => \N__29735\,
            I => \b2v_inst36.countZ0Z_11\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__29732\,
            I => \b2v_inst36.countZ0Z_11\
        );

    \I__6311\ : Odrv4
    port map (
            O => \N__29729\,
            I => \b2v_inst36.countZ0Z_11\
        );

    \I__6310\ : InMux
    port map (
            O => \N__29722\,
            I => \N__29718\
        );

    \I__6309\ : InMux
    port map (
            O => \N__29721\,
            I => \N__29715\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__29718\,
            I => \N__29710\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__29715\,
            I => \N__29710\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__29710\,
            I => \VR_READY_VCCIN_c\
        );

    \I__6305\ : CascadeMux
    port map (
            O => \N__29707\,
            I => \N__29703\
        );

    \I__6304\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29700\
        );

    \I__6303\ : InMux
    port map (
            O => \N__29703\,
            I => \N__29697\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__29700\,
            I => \N__29694\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__29697\,
            I => \N__29691\
        );

    \I__6300\ : Odrv4
    port map (
            O => \N__29694\,
            I => \VR_READY_VCCINAUX_c\
        );

    \I__6299\ : Odrv4
    port map (
            O => \N__29691\,
            I => \VR_READY_VCCINAUX_c\
        );

    \I__6298\ : IoInMux
    port map (
            O => \N__29686\,
            I => \N__29682\
        );

    \I__6297\ : IoInMux
    port map (
            O => \N__29685\,
            I => \N__29679\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__29682\,
            I => \N__29673\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__29679\,
            I => \N__29673\
        );

    \I__6294\ : CascadeMux
    port map (
            O => \N__29678\,
            I => \N__29667\
        );

    \I__6293\ : IoSpan4Mux
    port map (
            O => \N__29673\,
            I => \N__29664\
        );

    \I__6292\ : InMux
    port map (
            O => \N__29672\,
            I => \N__29661\
        );

    \I__6291\ : CascadeMux
    port map (
            O => \N__29671\,
            I => \N__29655\
        );

    \I__6290\ : CascadeMux
    port map (
            O => \N__29670\,
            I => \N__29649\
        );

    \I__6289\ : InMux
    port map (
            O => \N__29667\,
            I => \N__29646\
        );

    \I__6288\ : IoSpan4Mux
    port map (
            O => \N__29664\,
            I => \N__29643\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__29661\,
            I => \N__29640\
        );

    \I__6286\ : InMux
    port map (
            O => \N__29660\,
            I => \N__29635\
        );

    \I__6285\ : InMux
    port map (
            O => \N__29659\,
            I => \N__29630\
        );

    \I__6284\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29627\
        );

    \I__6283\ : InMux
    port map (
            O => \N__29655\,
            I => \N__29620\
        );

    \I__6282\ : InMux
    port map (
            O => \N__29654\,
            I => \N__29620\
        );

    \I__6281\ : InMux
    port map (
            O => \N__29653\,
            I => \N__29620\
        );

    \I__6280\ : InMux
    port map (
            O => \N__29652\,
            I => \N__29616\
        );

    \I__6279\ : InMux
    port map (
            O => \N__29649\,
            I => \N__29612\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__29646\,
            I => \N__29609\
        );

    \I__6277\ : Span4Mux_s2_h
    port map (
            O => \N__29643\,
            I => \N__29604\
        );

    \I__6276\ : Span4Mux_v
    port map (
            O => \N__29640\,
            I => \N__29604\
        );

    \I__6275\ : InMux
    port map (
            O => \N__29639\,
            I => \N__29601\
        );

    \I__6274\ : InMux
    port map (
            O => \N__29638\,
            I => \N__29598\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__29635\,
            I => \N__29595\
        );

    \I__6272\ : InMux
    port map (
            O => \N__29634\,
            I => \N__29590\
        );

    \I__6271\ : InMux
    port map (
            O => \N__29633\,
            I => \N__29590\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__29630\,
            I => \N__29583\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__29627\,
            I => \N__29583\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__29620\,
            I => \N__29583\
        );

    \I__6267\ : InMux
    port map (
            O => \N__29619\,
            I => \N__29580\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__29616\,
            I => \N__29577\
        );

    \I__6265\ : InMux
    port map (
            O => \N__29615\,
            I => \N__29574\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__29612\,
            I => \N__29571\
        );

    \I__6263\ : Span4Mux_v
    port map (
            O => \N__29609\,
            I => \N__29566\
        );

    \I__6262\ : Span4Mux_h
    port map (
            O => \N__29604\,
            I => \N__29566\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__29601\,
            I => \N__29553\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__29598\,
            I => \N__29553\
        );

    \I__6259\ : Span4Mux_h
    port map (
            O => \N__29595\,
            I => \N__29553\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__29590\,
            I => \N__29553\
        );

    \I__6257\ : Span4Mux_s3_v
    port map (
            O => \N__29583\,
            I => \N__29553\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__29580\,
            I => \N__29553\
        );

    \I__6255\ : Odrv12
    port map (
            O => \N__29577\,
            I => \SYNTHESIZED_WIRE_48_i_0_o3_2\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__29574\,
            I => \SYNTHESIZED_WIRE_48_i_0_o3_2\
        );

    \I__6253\ : Odrv12
    port map (
            O => \N__29571\,
            I => \SYNTHESIZED_WIRE_48_i_0_o3_2\
        );

    \I__6252\ : Odrv4
    port map (
            O => \N__29566\,
            I => \SYNTHESIZED_WIRE_48_i_0_o3_2\
        );

    \I__6251\ : Odrv4
    port map (
            O => \N__29553\,
            I => \SYNTHESIZED_WIRE_48_i_0_o3_2\
        );

    \I__6250\ : CascadeMux
    port map (
            O => \N__29542\,
            I => \b2v_inst6.N_413_cascade_\
        );

    \I__6249\ : CascadeMux
    port map (
            O => \N__29539\,
            I => \b2v_inst6.curr_state_7_1_cascade_\
        );

    \I__6248\ : InMux
    port map (
            O => \N__29536\,
            I => \N__29529\
        );

    \I__6247\ : InMux
    port map (
            O => \N__29535\,
            I => \N__29520\
        );

    \I__6246\ : InMux
    port map (
            O => \N__29534\,
            I => \N__29520\
        );

    \I__6245\ : InMux
    port map (
            O => \N__29533\,
            I => \N__29520\
        );

    \I__6244\ : InMux
    port map (
            O => \N__29532\,
            I => \N__29520\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__29529\,
            I => \b2v_inst6.curr_stateZ0Z_1\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__29520\,
            I => \b2v_inst6.curr_stateZ0Z_1\
        );

    \I__6241\ : CascadeMux
    port map (
            O => \N__29515\,
            I => \N__29507\
        );

    \I__6240\ : InMux
    port map (
            O => \N__29514\,
            I => \N__29502\
        );

    \I__6239\ : InMux
    port map (
            O => \N__29513\,
            I => \N__29493\
        );

    \I__6238\ : InMux
    port map (
            O => \N__29512\,
            I => \N__29493\
        );

    \I__6237\ : InMux
    port map (
            O => \N__29511\,
            I => \N__29493\
        );

    \I__6236\ : InMux
    port map (
            O => \N__29510\,
            I => \N__29493\
        );

    \I__6235\ : InMux
    port map (
            O => \N__29507\,
            I => \N__29486\
        );

    \I__6234\ : InMux
    port map (
            O => \N__29506\,
            I => \N__29486\
        );

    \I__6233\ : InMux
    port map (
            O => \N__29505\,
            I => \N__29486\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__29502\,
            I => \b2v_inst6.curr_stateZ0Z_0\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__29493\,
            I => \b2v_inst6.curr_stateZ0Z_0\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__29486\,
            I => \b2v_inst6.curr_stateZ0Z_0\
        );

    \I__6229\ : CascadeMux
    port map (
            O => \N__29479\,
            I => \b2v_inst6.curr_stateZ0Z_1_cascade_\
        );

    \I__6228\ : InMux
    port map (
            O => \N__29476\,
            I => \N__29466\
        );

    \I__6227\ : InMux
    port map (
            O => \N__29475\,
            I => \N__29466\
        );

    \I__6226\ : InMux
    port map (
            O => \N__29474\,
            I => \N__29457\
        );

    \I__6225\ : InMux
    port map (
            O => \N__29473\,
            I => \N__29457\
        );

    \I__6224\ : InMux
    port map (
            O => \N__29472\,
            I => \N__29457\
        );

    \I__6223\ : InMux
    port map (
            O => \N__29471\,
            I => \N__29457\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__29466\,
            I => \b2v_inst6.N_413\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__29457\,
            I => \b2v_inst6.N_413\
        );

    \I__6220\ : InMux
    port map (
            O => \N__29452\,
            I => \N__29449\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__29449\,
            I => \b2v_inst6.curr_state_1_1\
        );

    \I__6218\ : CascadeMux
    port map (
            O => \N__29446\,
            I => \b2v_inst36.countZ0Z_1_cascade_\
        );

    \I__6217\ : InMux
    port map (
            O => \N__29443\,
            I => \N__29440\
        );

    \I__6216\ : LocalMux
    port map (
            O => \N__29440\,
            I => \b2v_inst36.count_rst_13\
        );

    \I__6215\ : InMux
    port map (
            O => \N__29437\,
            I => \N__29434\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__29434\,
            I => \N__29431\
        );

    \I__6213\ : Span4Mux_s1_v
    port map (
            O => \N__29431\,
            I => \N__29427\
        );

    \I__6212\ : InMux
    port map (
            O => \N__29430\,
            I => \N__29424\
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__29427\,
            I => \b2v_inst36.countZ0Z_14\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__29424\,
            I => \b2v_inst36.countZ0Z_14\
        );

    \I__6209\ : InMux
    port map (
            O => \N__29419\,
            I => \N__29416\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__29416\,
            I => \N__29412\
        );

    \I__6207\ : InMux
    port map (
            O => \N__29415\,
            I => \N__29409\
        );

    \I__6206\ : Span4Mux_s3_h
    port map (
            O => \N__29412\,
            I => \N__29404\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__29409\,
            I => \N__29404\
        );

    \I__6204\ : Odrv4
    port map (
            O => \N__29404\,
            I => \b2v_inst36.countZ0Z_15\
        );

    \I__6203\ : InMux
    port map (
            O => \N__29401\,
            I => \N__29398\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__29398\,
            I => \b2v_inst36.count_1_1\
        );

    \I__6201\ : InMux
    port map (
            O => \N__29395\,
            I => \N__29392\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__29392\,
            I => \b2v_inst6.count_rst_10\
        );

    \I__6199\ : CascadeMux
    port map (
            O => \N__29389\,
            I => \b2v_inst6.count_rst_3_cascade_\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__29386\,
            I => \b2v_inst6.countZ0Z_4_cascade_\
        );

    \I__6197\ : InMux
    port map (
            O => \N__29383\,
            I => \N__29380\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__29380\,
            I => \b2v_inst6.count_3_4\
        );

    \I__6195\ : CascadeMux
    port map (
            O => \N__29377\,
            I => \G_2746_cascade_\
        );

    \I__6194\ : CascadeMux
    port map (
            O => \N__29374\,
            I => \b2v_inst6.curr_stateZ0Z_0_cascade_\
        );

    \I__6193\ : InMux
    port map (
            O => \N__29371\,
            I => \N__29368\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__29368\,
            I => \b2v_inst6.curr_state_2_0\
        );

    \I__6191\ : InMux
    port map (
            O => \N__29365\,
            I => \N__29355\
        );

    \I__6190\ : InMux
    port map (
            O => \N__29364\,
            I => \N__29355\
        );

    \I__6189\ : InMux
    port map (
            O => \N__29363\,
            I => \N__29355\
        );

    \I__6188\ : CascadeMux
    port map (
            O => \N__29362\,
            I => \N__29350\
        );

    \I__6187\ : LocalMux
    port map (
            O => \N__29355\,
            I => \N__29347\
        );

    \I__6186\ : InMux
    port map (
            O => \N__29354\,
            I => \N__29344\
        );

    \I__6185\ : CascadeMux
    port map (
            O => \N__29353\,
            I => \N__29341\
        );

    \I__6184\ : InMux
    port map (
            O => \N__29350\,
            I => \N__29338\
        );

    \I__6183\ : Span4Mux_v
    port map (
            O => \N__29347\,
            I => \N__29335\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__29344\,
            I => \N__29332\
        );

    \I__6181\ : InMux
    port map (
            O => \N__29341\,
            I => \N__29329\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__29338\,
            I => \N__29325\
        );

    \I__6179\ : Span4Mux_h
    port map (
            O => \N__29335\,
            I => \N__29318\
        );

    \I__6178\ : Span4Mux_v
    port map (
            O => \N__29332\,
            I => \N__29318\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__29329\,
            I => \N__29318\
        );

    \I__6176\ : InMux
    port map (
            O => \N__29328\,
            I => \N__29315\
        );

    \I__6175\ : Span4Mux_v
    port map (
            O => \N__29325\,
            I => \N__29311\
        );

    \I__6174\ : Span4Mux_h
    port map (
            O => \N__29318\,
            I => \N__29308\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__29315\,
            I => \N__29305\
        );

    \I__6172\ : InMux
    port map (
            O => \N__29314\,
            I => \N__29302\
        );

    \I__6171\ : Odrv4
    port map (
            O => \N__29311\,
            I => \b2v_inst11.N_158\
        );

    \I__6170\ : Odrv4
    port map (
            O => \N__29308\,
            I => \b2v_inst11.N_158\
        );

    \I__6169\ : Odrv12
    port map (
            O => \N__29305\,
            I => \b2v_inst11.N_158\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__29302\,
            I => \b2v_inst11.N_158\
        );

    \I__6167\ : CascadeMux
    port map (
            O => \N__29293\,
            I => \N__29290\
        );

    \I__6166\ : InMux
    port map (
            O => \N__29290\,
            I => \N__29287\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__29287\,
            I => \N__29281\
        );

    \I__6164\ : InMux
    port map (
            O => \N__29286\,
            I => \N__29278\
        );

    \I__6163\ : InMux
    port map (
            O => \N__29285\,
            I => \N__29274\
        );

    \I__6162\ : InMux
    port map (
            O => \N__29284\,
            I => \N__29269\
        );

    \I__6161\ : Span4Mux_v
    port map (
            O => \N__29281\,
            I => \N__29265\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__29278\,
            I => \N__29262\
        );

    \I__6159\ : InMux
    port map (
            O => \N__29277\,
            I => \N__29259\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__29274\,
            I => \N__29256\
        );

    \I__6157\ : InMux
    port map (
            O => \N__29273\,
            I => \N__29251\
        );

    \I__6156\ : InMux
    port map (
            O => \N__29272\,
            I => \N__29251\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__29269\,
            I => \N__29243\
        );

    \I__6154\ : InMux
    port map (
            O => \N__29268\,
            I => \N__29240\
        );

    \I__6153\ : Span4Mux_s1_v
    port map (
            O => \N__29265\,
            I => \N__29228\
        );

    \I__6152\ : Span4Mux_v
    port map (
            O => \N__29262\,
            I => \N__29228\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__29259\,
            I => \N__29228\
        );

    \I__6150\ : Span4Mux_s3_h
    port map (
            O => \N__29256\,
            I => \N__29223\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__29251\,
            I => \N__29223\
        );

    \I__6148\ : CascadeMux
    port map (
            O => \N__29250\,
            I => \N__29218\
        );

    \I__6147\ : CascadeMux
    port map (
            O => \N__29249\,
            I => \N__29211\
        );

    \I__6146\ : CascadeMux
    port map (
            O => \N__29248\,
            I => \N__29208\
        );

    \I__6145\ : CascadeMux
    port map (
            O => \N__29247\,
            I => \N__29205\
        );

    \I__6144\ : CascadeMux
    port map (
            O => \N__29246\,
            I => \N__29202\
        );

    \I__6143\ : Span4Mux_s2_v
    port map (
            O => \N__29243\,
            I => \N__29197\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__29240\,
            I => \N__29194\
        );

    \I__6141\ : InMux
    port map (
            O => \N__29239\,
            I => \N__29191\
        );

    \I__6140\ : InMux
    port map (
            O => \N__29238\,
            I => \N__29186\
        );

    \I__6139\ : InMux
    port map (
            O => \N__29237\,
            I => \N__29186\
        );

    \I__6138\ : InMux
    port map (
            O => \N__29236\,
            I => \N__29183\
        );

    \I__6137\ : InMux
    port map (
            O => \N__29235\,
            I => \N__29180\
        );

    \I__6136\ : Span4Mux_h
    port map (
            O => \N__29228\,
            I => \N__29175\
        );

    \I__6135\ : Span4Mux_h
    port map (
            O => \N__29223\,
            I => \N__29175\
        );

    \I__6134\ : InMux
    port map (
            O => \N__29222\,
            I => \N__29164\
        );

    \I__6133\ : InMux
    port map (
            O => \N__29221\,
            I => \N__29164\
        );

    \I__6132\ : InMux
    port map (
            O => \N__29218\,
            I => \N__29164\
        );

    \I__6131\ : InMux
    port map (
            O => \N__29217\,
            I => \N__29164\
        );

    \I__6130\ : InMux
    port map (
            O => \N__29216\,
            I => \N__29164\
        );

    \I__6129\ : InMux
    port map (
            O => \N__29215\,
            I => \N__29147\
        );

    \I__6128\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29147\
        );

    \I__6127\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29147\
        );

    \I__6126\ : InMux
    port map (
            O => \N__29208\,
            I => \N__29147\
        );

    \I__6125\ : InMux
    port map (
            O => \N__29205\,
            I => \N__29147\
        );

    \I__6124\ : InMux
    port map (
            O => \N__29202\,
            I => \N__29147\
        );

    \I__6123\ : InMux
    port map (
            O => \N__29201\,
            I => \N__29147\
        );

    \I__6122\ : InMux
    port map (
            O => \N__29200\,
            I => \N__29147\
        );

    \I__6121\ : Odrv4
    port map (
            O => \N__29197\,
            I => \b2v_inst11.N_3046_i\
        );

    \I__6120\ : Odrv12
    port map (
            O => \N__29194\,
            I => \b2v_inst11.N_3046_i\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__29191\,
            I => \b2v_inst11.N_3046_i\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__29186\,
            I => \b2v_inst11.N_3046_i\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__29183\,
            I => \b2v_inst11.N_3046_i\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__29180\,
            I => \b2v_inst11.N_3046_i\
        );

    \I__6115\ : Odrv4
    port map (
            O => \N__29175\,
            I => \b2v_inst11.N_3046_i\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__29164\,
            I => \b2v_inst11.N_3046_i\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__29147\,
            I => \b2v_inst11.N_3046_i\
        );

    \I__6112\ : InMux
    port map (
            O => \N__29128\,
            I => \N__29125\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__29125\,
            I => \b2v_inst11.g3_0\
        );

    \I__6110\ : CascadeMux
    port map (
            O => \N__29122\,
            I => \b2v_inst11.g2_0_cascade_\
        );

    \I__6109\ : IoInMux
    port map (
            O => \N__29119\,
            I => \N__29116\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__29116\,
            I => \N__29113\
        );

    \I__6107\ : IoSpan4Mux
    port map (
            O => \N__29113\,
            I => \N__29108\
        );

    \I__6106\ : InMux
    port map (
            O => \N__29112\,
            I => \N__29103\
        );

    \I__6105\ : InMux
    port map (
            O => \N__29111\,
            I => \N__29103\
        );

    \I__6104\ : Span4Mux_s3_h
    port map (
            O => \N__29108\,
            I => \N__29100\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__29103\,
            I => \N__29096\
        );

    \I__6102\ : Span4Mux_v
    port map (
            O => \N__29100\,
            I => \N__29089\
        );

    \I__6101\ : InMux
    port map (
            O => \N__29099\,
            I => \N__29086\
        );

    \I__6100\ : Sp12to4
    port map (
            O => \N__29096\,
            I => \N__29082\
        );

    \I__6099\ : InMux
    port map (
            O => \N__29095\,
            I => \N__29079\
        );

    \I__6098\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29076\
        );

    \I__6097\ : InMux
    port map (
            O => \N__29093\,
            I => \N__29073\
        );

    \I__6096\ : InMux
    port map (
            O => \N__29092\,
            I => \N__29068\
        );

    \I__6095\ : Span4Mux_v
    port map (
            O => \N__29089\,
            I => \N__29063\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__29086\,
            I => \N__29063\
        );

    \I__6093\ : InMux
    port map (
            O => \N__29085\,
            I => \N__29060\
        );

    \I__6092\ : Span12Mux_s7_h
    port map (
            O => \N__29082\,
            I => \N__29055\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__29079\,
            I => \N__29055\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__29076\,
            I => \N__29050\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__29073\,
            I => \N__29050\
        );

    \I__6088\ : InMux
    port map (
            O => \N__29072\,
            I => \N__29047\
        );

    \I__6087\ : InMux
    port map (
            O => \N__29071\,
            I => \N__29044\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__29068\,
            I => \N__29037\
        );

    \I__6085\ : Span4Mux_h
    port map (
            O => \N__29063\,
            I => \N__29037\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__29060\,
            I => \N__29037\
        );

    \I__6083\ : Span12Mux_s2_v
    port map (
            O => \N__29055\,
            I => \N__29034\
        );

    \I__6082\ : Odrv4
    port map (
            O => \N__29050\,
            I => \RSMRSTn_RNI8DFE\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__29047\,
            I => \RSMRSTn_RNI8DFE\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__29044\,
            I => \RSMRSTn_RNI8DFE\
        );

    \I__6079\ : Odrv4
    port map (
            O => \N__29037\,
            I => \RSMRSTn_RNI8DFE\
        );

    \I__6078\ : Odrv12
    port map (
            O => \N__29034\,
            I => \RSMRSTn_RNI8DFE\
        );

    \I__6077\ : InMux
    port map (
            O => \N__29023\,
            I => \N__29020\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__29020\,
            I => \N__29017\
        );

    \I__6075\ : Span4Mux_s3_v
    port map (
            O => \N__29017\,
            I => \N__29014\
        );

    \I__6074\ : Odrv4
    port map (
            O => \N__29014\,
            I => \b2v_inst11.N_228_N_0\
        );

    \I__6073\ : InMux
    port map (
            O => \N__29011\,
            I => \N__29008\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__29008\,
            I => \N__29005\
        );

    \I__6071\ : Odrv4
    port map (
            O => \N__29005\,
            I => \b2v_inst6.delayed_vccin_vccinaux_okZ0\
        );

    \I__6070\ : InMux
    port map (
            O => \N__29002\,
            I => \N__28999\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__28999\,
            I => \b2v_inst11.g1_4_2_0\
        );

    \I__6068\ : CascadeMux
    port map (
            O => \N__28996\,
            I => \N__28987\
        );

    \I__6067\ : CascadeMux
    port map (
            O => \N__28995\,
            I => \N__28984\
        );

    \I__6066\ : InMux
    port map (
            O => \N__28994\,
            I => \N__28981\
        );

    \I__6065\ : InMux
    port map (
            O => \N__28993\,
            I => \N__28978\
        );

    \I__6064\ : CascadeMux
    port map (
            O => \N__28992\,
            I => \N__28975\
        );

    \I__6063\ : InMux
    port map (
            O => \N__28991\,
            I => \N__28966\
        );

    \I__6062\ : InMux
    port map (
            O => \N__28990\,
            I => \N__28966\
        );

    \I__6061\ : InMux
    port map (
            O => \N__28987\,
            I => \N__28963\
        );

    \I__6060\ : InMux
    port map (
            O => \N__28984\,
            I => \N__28959\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__28981\,
            I => \N__28950\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__28978\,
            I => \N__28947\
        );

    \I__6057\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28944\
        );

    \I__6056\ : CascadeMux
    port map (
            O => \N__28974\,
            I => \N__28941\
        );

    \I__6055\ : CascadeMux
    port map (
            O => \N__28973\,
            I => \N__28937\
        );

    \I__6054\ : InMux
    port map (
            O => \N__28972\,
            I => \N__28931\
        );

    \I__6053\ : InMux
    port map (
            O => \N__28971\,
            I => \N__28927\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__28966\,
            I => \N__28924\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__28963\,
            I => \N__28921\
        );

    \I__6050\ : CascadeMux
    port map (
            O => \N__28962\,
            I => \N__28918\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__28959\,
            I => \N__28915\
        );

    \I__6048\ : InMux
    port map (
            O => \N__28958\,
            I => \N__28910\
        );

    \I__6047\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28910\
        );

    \I__6046\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28901\
        );

    \I__6045\ : InMux
    port map (
            O => \N__28955\,
            I => \N__28901\
        );

    \I__6044\ : InMux
    port map (
            O => \N__28954\,
            I => \N__28901\
        );

    \I__6043\ : InMux
    port map (
            O => \N__28953\,
            I => \N__28901\
        );

    \I__6042\ : Span4Mux_v
    port map (
            O => \N__28950\,
            I => \N__28896\
        );

    \I__6041\ : Span4Mux_v
    port map (
            O => \N__28947\,
            I => \N__28896\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__28944\,
            I => \N__28893\
        );

    \I__6039\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28888\
        );

    \I__6038\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28888\
        );

    \I__6037\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28879\
        );

    \I__6036\ : InMux
    port map (
            O => \N__28936\,
            I => \N__28879\
        );

    \I__6035\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28879\
        );

    \I__6034\ : InMux
    port map (
            O => \N__28934\,
            I => \N__28879\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__28931\,
            I => \N__28876\
        );

    \I__6032\ : InMux
    port map (
            O => \N__28930\,
            I => \N__28873\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__28927\,
            I => \N__28866\
        );

    \I__6030\ : Span4Mux_v
    port map (
            O => \N__28924\,
            I => \N__28866\
        );

    \I__6029\ : Span4Mux_s3_v
    port map (
            O => \N__28921\,
            I => \N__28866\
        );

    \I__6028\ : InMux
    port map (
            O => \N__28918\,
            I => \N__28863\
        );

    \I__6027\ : Span4Mux_v
    port map (
            O => \N__28915\,
            I => \N__28856\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__28910\,
            I => \N__28856\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__28901\,
            I => \N__28856\
        );

    \I__6024\ : Odrv4
    port map (
            O => \N__28896\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__6023\ : Odrv12
    port map (
            O => \N__28893\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__28888\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__28879\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__6020\ : Odrv4
    port map (
            O => \N__28876\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__28873\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__6018\ : Odrv4
    port map (
            O => \N__28866\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__28863\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__28856\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__6015\ : CascadeMux
    port map (
            O => \N__28837\,
            I => \N__28833\
        );

    \I__6014\ : InMux
    port map (
            O => \N__28836\,
            I => \N__28825\
        );

    \I__6013\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28822\
        );

    \I__6012\ : InMux
    port map (
            O => \N__28832\,
            I => \N__28819\
        );

    \I__6011\ : InMux
    port map (
            O => \N__28831\,
            I => \N__28814\
        );

    \I__6010\ : InMux
    port map (
            O => \N__28830\,
            I => \N__28814\
        );

    \I__6009\ : InMux
    port map (
            O => \N__28829\,
            I => \N__28811\
        );

    \I__6008\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28808\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__28825\,
            I => \N__28805\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__28822\,
            I => \N__28802\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__28819\,
            I => \N__28799\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__28814\,
            I => \N__28795\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__28811\,
            I => \N__28792\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__28808\,
            I => \N__28789\
        );

    \I__6001\ : Span4Mux_h
    port map (
            O => \N__28805\,
            I => \N__28784\
        );

    \I__6000\ : Span4Mux_h
    port map (
            O => \N__28802\,
            I => \N__28784\
        );

    \I__5999\ : Span4Mux_v
    port map (
            O => \N__28799\,
            I => \N__28781\
        );

    \I__5998\ : InMux
    port map (
            O => \N__28798\,
            I => \N__28778\
        );

    \I__5997\ : Span4Mux_v
    port map (
            O => \N__28795\,
            I => \N__28773\
        );

    \I__5996\ : Span4Mux_v
    port map (
            O => \N__28792\,
            I => \N__28773\
        );

    \I__5995\ : Odrv4
    port map (
            O => \N__28789\,
            I => \N_19_i\
        );

    \I__5994\ : Odrv4
    port map (
            O => \N__28784\,
            I => \N_19_i\
        );

    \I__5993\ : Odrv4
    port map (
            O => \N__28781\,
            I => \N_19_i\
        );

    \I__5992\ : LocalMux
    port map (
            O => \N__28778\,
            I => \N_19_i\
        );

    \I__5991\ : Odrv4
    port map (
            O => \N__28773\,
            I => \N_19_i\
        );

    \I__5990\ : InMux
    port map (
            O => \N__28762\,
            I => \N__28756\
        );

    \I__5989\ : InMux
    port map (
            O => \N__28761\,
            I => \N__28756\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__28756\,
            I => \b2v_inst11.g0_8_0_0\
        );

    \I__5987\ : CascadeMux
    port map (
            O => \N__28753\,
            I => \N__28748\
        );

    \I__5986\ : CascadeMux
    port map (
            O => \N__28752\,
            I => \N__28741\
        );

    \I__5985\ : CascadeMux
    port map (
            O => \N__28751\,
            I => \N__28736\
        );

    \I__5984\ : InMux
    port map (
            O => \N__28748\,
            I => \N__28733\
        );

    \I__5983\ : InMux
    port map (
            O => \N__28747\,
            I => \N__28728\
        );

    \I__5982\ : InMux
    port map (
            O => \N__28746\,
            I => \N__28725\
        );

    \I__5981\ : InMux
    port map (
            O => \N__28745\,
            I => \N__28722\
        );

    \I__5980\ : InMux
    port map (
            O => \N__28744\,
            I => \N__28717\
        );

    \I__5979\ : InMux
    port map (
            O => \N__28741\,
            I => \N__28717\
        );

    \I__5978\ : InMux
    port map (
            O => \N__28740\,
            I => \N__28712\
        );

    \I__5977\ : InMux
    port map (
            O => \N__28739\,
            I => \N__28712\
        );

    \I__5976\ : InMux
    port map (
            O => \N__28736\,
            I => \N__28709\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__28733\,
            I => \N__28702\
        );

    \I__5974\ : InMux
    port map (
            O => \N__28732\,
            I => \N__28697\
        );

    \I__5973\ : InMux
    port map (
            O => \N__28731\,
            I => \N__28697\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__28728\,
            I => \N__28692\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__28725\,
            I => \N__28692\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__28722\,
            I => \N__28685\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__28717\,
            I => \N__28685\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__28712\,
            I => \N__28685\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__28709\,
            I => \N__28682\
        );

    \I__5966\ : InMux
    port map (
            O => \N__28708\,
            I => \N__28679\
        );

    \I__5965\ : InMux
    port map (
            O => \N__28707\,
            I => \N__28675\
        );

    \I__5964\ : InMux
    port map (
            O => \N__28706\,
            I => \N__28669\
        );

    \I__5963\ : InMux
    port map (
            O => \N__28705\,
            I => \N__28669\
        );

    \I__5962\ : Span4Mux_v
    port map (
            O => \N__28702\,
            I => \N__28663\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__28697\,
            I => \N__28663\
        );

    \I__5960\ : Span4Mux_v
    port map (
            O => \N__28692\,
            I => \N__28654\
        );

    \I__5959\ : Span4Mux_h
    port map (
            O => \N__28685\,
            I => \N__28654\
        );

    \I__5958\ : Span4Mux_v
    port map (
            O => \N__28682\,
            I => \N__28654\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__28679\,
            I => \N__28654\
        );

    \I__5956\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28651\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__28675\,
            I => \N__28648\
        );

    \I__5954\ : InMux
    port map (
            O => \N__28674\,
            I => \N__28645\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__28669\,
            I => \N__28642\
        );

    \I__5952\ : InMux
    port map (
            O => \N__28668\,
            I => \N__28639\
        );

    \I__5951\ : IoSpan4Mux
    port map (
            O => \N__28663\,
            I => \N__28636\
        );

    \I__5950\ : Span4Mux_h
    port map (
            O => \N__28654\,
            I => \N__28633\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__28651\,
            I => \N__28630\
        );

    \I__5948\ : Span4Mux_h
    port map (
            O => \N__28648\,
            I => \N__28625\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__28645\,
            I => \N__28625\
        );

    \I__5946\ : Span4Mux_h
    port map (
            O => \N__28642\,
            I => \N__28620\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__28639\,
            I => \N__28620\
        );

    \I__5944\ : IoSpan4Mux
    port map (
            O => \N__28636\,
            I => \N__28617\
        );

    \I__5943\ : Span4Mux_v
    port map (
            O => \N__28633\,
            I => \N__28614\
        );

    \I__5942\ : IoSpan4Mux
    port map (
            O => \N__28630\,
            I => \N__28611\
        );

    \I__5941\ : IoSpan4Mux
    port map (
            O => \N__28625\,
            I => \N__28606\
        );

    \I__5940\ : IoSpan4Mux
    port map (
            O => \N__28620\,
            I => \N__28606\
        );

    \I__5939\ : Odrv4
    port map (
            O => \N__28617\,
            I => \SLP_S4n_c\
        );

    \I__5938\ : Odrv4
    port map (
            O => \N__28614\,
            I => \SLP_S4n_c\
        );

    \I__5937\ : Odrv4
    port map (
            O => \N__28611\,
            I => \SLP_S4n_c\
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__28606\,
            I => \SLP_S4n_c\
        );

    \I__5935\ : InMux
    port map (
            O => \N__28597\,
            I => \N__28594\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__28594\,
            I => \N__28588\
        );

    \I__5933\ : InMux
    port map (
            O => \N__28593\,
            I => \N__28583\
        );

    \I__5932\ : InMux
    port map (
            O => \N__28592\,
            I => \N__28583\
        );

    \I__5931\ : InMux
    port map (
            O => \N__28591\,
            I => \N__28578\
        );

    \I__5930\ : Span4Mux_h
    port map (
            O => \N__28588\,
            I => \N__28567\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__28583\,
            I => \N__28567\
        );

    \I__5928\ : InMux
    port map (
            O => \N__28582\,
            I => \N__28564\
        );

    \I__5927\ : InMux
    port map (
            O => \N__28581\,
            I => \N__28561\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__28578\,
            I => \N__28556\
        );

    \I__5925\ : InMux
    port map (
            O => \N__28577\,
            I => \N__28553\
        );

    \I__5924\ : InMux
    port map (
            O => \N__28576\,
            I => \N__28550\
        );

    \I__5923\ : InMux
    port map (
            O => \N__28575\,
            I => \N__28545\
        );

    \I__5922\ : InMux
    port map (
            O => \N__28574\,
            I => \N__28542\
        );

    \I__5921\ : InMux
    port map (
            O => \N__28573\,
            I => \N__28539\
        );

    \I__5920\ : InMux
    port map (
            O => \N__28572\,
            I => \N__28536\
        );

    \I__5919\ : Span4Mux_v
    port map (
            O => \N__28567\,
            I => \N__28529\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__28564\,
            I => \N__28529\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__28561\,
            I => \N__28529\
        );

    \I__5916\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28524\
        );

    \I__5915\ : InMux
    port map (
            O => \N__28559\,
            I => \N__28524\
        );

    \I__5914\ : Span4Mux_v
    port map (
            O => \N__28556\,
            I => \N__28519\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__28553\,
            I => \N__28519\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__28550\,
            I => \N__28516\
        );

    \I__5911\ : InMux
    port map (
            O => \N__28549\,
            I => \N__28511\
        );

    \I__5910\ : InMux
    port map (
            O => \N__28548\,
            I => \N__28511\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__28545\,
            I => \N__28504\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__28542\,
            I => \N__28504\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__28539\,
            I => \N__28504\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__28536\,
            I => \N__28501\
        );

    \I__5905\ : Span4Mux_h
    port map (
            O => \N__28529\,
            I => \N__28496\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__28524\,
            I => \N__28496\
        );

    \I__5903\ : Span4Mux_v
    port map (
            O => \N__28519\,
            I => \N__28489\
        );

    \I__5902\ : Span4Mux_h
    port map (
            O => \N__28516\,
            I => \N__28489\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__28511\,
            I => \N__28489\
        );

    \I__5900\ : Span12Mux_s9_h
    port map (
            O => \N__28504\,
            I => \N__28485\
        );

    \I__5899\ : Span4Mux_v
    port map (
            O => \N__28501\,
            I => \N__28482\
        );

    \I__5898\ : IoSpan4Mux
    port map (
            O => \N__28496\,
            I => \N__28479\
        );

    \I__5897\ : Span4Mux_h
    port map (
            O => \N__28489\,
            I => \N__28476\
        );

    \I__5896\ : InMux
    port map (
            O => \N__28488\,
            I => \N__28473\
        );

    \I__5895\ : Odrv12
    port map (
            O => \N__28485\,
            I => \GPIO_FPGA_PCH_5_c\
        );

    \I__5894\ : Odrv4
    port map (
            O => \N__28482\,
            I => \GPIO_FPGA_PCH_5_c\
        );

    \I__5893\ : Odrv4
    port map (
            O => \N__28479\,
            I => \GPIO_FPGA_PCH_5_c\
        );

    \I__5892\ : Odrv4
    port map (
            O => \N__28476\,
            I => \GPIO_FPGA_PCH_5_c\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__28473\,
            I => \GPIO_FPGA_PCH_5_c\
        );

    \I__5890\ : InMux
    port map (
            O => \N__28462\,
            I => \N__28447\
        );

    \I__5889\ : InMux
    port map (
            O => \N__28461\,
            I => \N__28447\
        );

    \I__5888\ : InMux
    port map (
            O => \N__28460\,
            I => \N__28447\
        );

    \I__5887\ : InMux
    port map (
            O => \N__28459\,
            I => \N__28440\
        );

    \I__5886\ : InMux
    port map (
            O => \N__28458\,
            I => \N__28440\
        );

    \I__5885\ : InMux
    port map (
            O => \N__28457\,
            I => \N__28440\
        );

    \I__5884\ : InMux
    port map (
            O => \N__28456\,
            I => \N__28435\
        );

    \I__5883\ : InMux
    port map (
            O => \N__28455\,
            I => \N__28435\
        );

    \I__5882\ : InMux
    port map (
            O => \N__28454\,
            I => \N__28430\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__28447\,
            I => \N__28426\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__28440\,
            I => \N__28423\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__28435\,
            I => \N__28420\
        );

    \I__5878\ : InMux
    port map (
            O => \N__28434\,
            I => \N__28417\
        );

    \I__5877\ : CascadeMux
    port map (
            O => \N__28433\,
            I => \N__28414\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__28430\,
            I => \N__28409\
        );

    \I__5875\ : InMux
    port map (
            O => \N__28429\,
            I => \N__28406\
        );

    \I__5874\ : Span4Mux_s3_v
    port map (
            O => \N__28426\,
            I => \N__28396\
        );

    \I__5873\ : Span4Mux_s3_h
    port map (
            O => \N__28423\,
            I => \N__28396\
        );

    \I__5872\ : Span4Mux_v
    port map (
            O => \N__28420\,
            I => \N__28396\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__28417\,
            I => \N__28392\
        );

    \I__5870\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28389\
        );

    \I__5869\ : InMux
    port map (
            O => \N__28413\,
            I => \N__28386\
        );

    \I__5868\ : InMux
    port map (
            O => \N__28412\,
            I => \N__28383\
        );

    \I__5867\ : Span4Mux_s3_v
    port map (
            O => \N__28409\,
            I => \N__28378\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__28406\,
            I => \N__28378\
        );

    \I__5865\ : InMux
    port map (
            O => \N__28405\,
            I => \N__28371\
        );

    \I__5864\ : InMux
    port map (
            O => \N__28404\,
            I => \N__28371\
        );

    \I__5863\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28371\
        );

    \I__5862\ : Span4Mux_h
    port map (
            O => \N__28396\,
            I => \N__28368\
        );

    \I__5861\ : InMux
    port map (
            O => \N__28395\,
            I => \N__28365\
        );

    \I__5860\ : Odrv4
    port map (
            O => \N__28392\,
            I => \b2v_inst11.func_state\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__28389\,
            I => \b2v_inst11.func_state\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__28386\,
            I => \b2v_inst11.func_state\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__28383\,
            I => \b2v_inst11.func_state\
        );

    \I__5856\ : Odrv4
    port map (
            O => \N__28378\,
            I => \b2v_inst11.func_state\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__28371\,
            I => \b2v_inst11.func_state\
        );

    \I__5854\ : Odrv4
    port map (
            O => \N__28368\,
            I => \b2v_inst11.func_state\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__28365\,
            I => \b2v_inst11.func_state\
        );

    \I__5852\ : InMux
    port map (
            O => \N__28348\,
            I => \N__28340\
        );

    \I__5851\ : InMux
    port map (
            O => \N__28347\,
            I => \N__28337\
        );

    \I__5850\ : CascadeMux
    port map (
            O => \N__28346\,
            I => \N__28333\
        );

    \I__5849\ : CascadeMux
    port map (
            O => \N__28345\,
            I => \N__28329\
        );

    \I__5848\ : CascadeMux
    port map (
            O => \N__28344\,
            I => \N__28326\
        );

    \I__5847\ : CascadeMux
    port map (
            O => \N__28343\,
            I => \N__28323\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__28340\,
            I => \N__28317\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__28337\,
            I => \N__28317\
        );

    \I__5844\ : InMux
    port map (
            O => \N__28336\,
            I => \N__28312\
        );

    \I__5843\ : InMux
    port map (
            O => \N__28333\,
            I => \N__28312\
        );

    \I__5842\ : InMux
    port map (
            O => \N__28332\,
            I => \N__28304\
        );

    \I__5841\ : InMux
    port map (
            O => \N__28329\,
            I => \N__28301\
        );

    \I__5840\ : InMux
    port map (
            O => \N__28326\,
            I => \N__28298\
        );

    \I__5839\ : InMux
    port map (
            O => \N__28323\,
            I => \N__28293\
        );

    \I__5838\ : InMux
    port map (
            O => \N__28322\,
            I => \N__28293\
        );

    \I__5837\ : Span4Mux_h
    port map (
            O => \N__28317\,
            I => \N__28287\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__28312\,
            I => \N__28284\
        );

    \I__5835\ : InMux
    port map (
            O => \N__28311\,
            I => \N__28277\
        );

    \I__5834\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28277\
        );

    \I__5833\ : InMux
    port map (
            O => \N__28309\,
            I => \N__28277\
        );

    \I__5832\ : CascadeMux
    port map (
            O => \N__28308\,
            I => \N__28273\
        );

    \I__5831\ : InMux
    port map (
            O => \N__28307\,
            I => \N__28270\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__28304\,
            I => \N__28265\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__28301\,
            I => \N__28265\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__28298\,
            I => \N__28260\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__28293\,
            I => \N__28260\
        );

    \I__5826\ : InMux
    port map (
            O => \N__28292\,
            I => \N__28257\
        );

    \I__5825\ : InMux
    port map (
            O => \N__28291\,
            I => \N__28254\
        );

    \I__5824\ : CascadeMux
    port map (
            O => \N__28290\,
            I => \N__28249\
        );

    \I__5823\ : Span4Mux_v
    port map (
            O => \N__28287\,
            I => \N__28244\
        );

    \I__5822\ : Span4Mux_h
    port map (
            O => \N__28284\,
            I => \N__28244\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__28277\,
            I => \N__28241\
        );

    \I__5820\ : InMux
    port map (
            O => \N__28276\,
            I => \N__28238\
        );

    \I__5819\ : InMux
    port map (
            O => \N__28273\,
            I => \N__28235\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__28270\,
            I => \N__28232\
        );

    \I__5817\ : Span4Mux_h
    port map (
            O => \N__28265\,
            I => \N__28223\
        );

    \I__5816\ : Span4Mux_h
    port map (
            O => \N__28260\,
            I => \N__28223\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__28257\,
            I => \N__28223\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__28254\,
            I => \N__28223\
        );

    \I__5813\ : InMux
    port map (
            O => \N__28253\,
            I => \N__28220\
        );

    \I__5812\ : InMux
    port map (
            O => \N__28252\,
            I => \N__28216\
        );

    \I__5811\ : InMux
    port map (
            O => \N__28249\,
            I => \N__28213\
        );

    \I__5810\ : IoSpan4Mux
    port map (
            O => \N__28244\,
            I => \N__28210\
        );

    \I__5809\ : Span4Mux_v
    port map (
            O => \N__28241\,
            I => \N__28203\
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__28238\,
            I => \N__28203\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__28235\,
            I => \N__28203\
        );

    \I__5806\ : Span4Mux_v
    port map (
            O => \N__28232\,
            I => \N__28196\
        );

    \I__5805\ : Span4Mux_h
    port map (
            O => \N__28223\,
            I => \N__28196\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__28220\,
            I => \N__28196\
        );

    \I__5803\ : InMux
    port map (
            O => \N__28219\,
            I => \N__28193\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__28216\,
            I => \N__28188\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__28213\,
            I => \N__28188\
        );

    \I__5800\ : Span4Mux_s0_v
    port map (
            O => \N__28210\,
            I => \N__28179\
        );

    \I__5799\ : Span4Mux_h
    port map (
            O => \N__28203\,
            I => \N__28179\
        );

    \I__5798\ : Span4Mux_v
    port map (
            O => \N__28196\,
            I => \N__28179\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__28193\,
            I => \N__28179\
        );

    \I__5796\ : Span12Mux_s10_h
    port map (
            O => \N__28188\,
            I => \N__28176\
        );

    \I__5795\ : Span4Mux_h
    port map (
            O => \N__28179\,
            I => \N__28173\
        );

    \I__5794\ : Odrv12
    port map (
            O => \N__28176\,
            I => \SLP_S3n_c\
        );

    \I__5793\ : Odrv4
    port map (
            O => \N__28173\,
            I => \SLP_S3n_c\
        );

    \I__5792\ : InMux
    port map (
            O => \N__28168\,
            I => \N__28160\
        );

    \I__5791\ : InMux
    port map (
            O => \N__28167\,
            I => \N__28154\
        );

    \I__5790\ : InMux
    port map (
            O => \N__28166\,
            I => \N__28148\
        );

    \I__5789\ : InMux
    port map (
            O => \N__28165\,
            I => \N__28148\
        );

    \I__5788\ : InMux
    port map (
            O => \N__28164\,
            I => \N__28143\
        );

    \I__5787\ : InMux
    port map (
            O => \N__28163\,
            I => \N__28143\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__28160\,
            I => \N__28137\
        );

    \I__5785\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28130\
        );

    \I__5784\ : InMux
    port map (
            O => \N__28158\,
            I => \N__28130\
        );

    \I__5783\ : InMux
    port map (
            O => \N__28157\,
            I => \N__28130\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__28154\,
            I => \N__28127\
        );

    \I__5781\ : InMux
    port map (
            O => \N__28153\,
            I => \N__28124\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__28148\,
            I => \N__28119\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__28143\,
            I => \N__28119\
        );

    \I__5778\ : InMux
    port map (
            O => \N__28142\,
            I => \N__28114\
        );

    \I__5777\ : InMux
    port map (
            O => \N__28141\,
            I => \N__28111\
        );

    \I__5776\ : InMux
    port map (
            O => \N__28140\,
            I => \N__28108\
        );

    \I__5775\ : Span4Mux_v
    port map (
            O => \N__28137\,
            I => \N__28102\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__28130\,
            I => \N__28102\
        );

    \I__5773\ : Span4Mux_v
    port map (
            O => \N__28127\,
            I => \N__28097\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__28124\,
            I => \N__28097\
        );

    \I__5771\ : Span4Mux_v
    port map (
            O => \N__28119\,
            I => \N__28093\
        );

    \I__5770\ : InMux
    port map (
            O => \N__28118\,
            I => \N__28090\
        );

    \I__5769\ : InMux
    port map (
            O => \N__28117\,
            I => \N__28087\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__28114\,
            I => \N__28080\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__28111\,
            I => \N__28080\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__28108\,
            I => \N__28080\
        );

    \I__5765\ : InMux
    port map (
            O => \N__28107\,
            I => \N__28077\
        );

    \I__5764\ : Span4Mux_s2_v
    port map (
            O => \N__28102\,
            I => \N__28074\
        );

    \I__5763\ : Span4Mux_h
    port map (
            O => \N__28097\,
            I => \N__28071\
        );

    \I__5762\ : InMux
    port map (
            O => \N__28096\,
            I => \N__28068\
        );

    \I__5761\ : Sp12to4
    port map (
            O => \N__28093\,
            I => \N__28063\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__28090\,
            I => \N__28063\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__28087\,
            I => \N__28056\
        );

    \I__5758\ : Span4Mux_v
    port map (
            O => \N__28080\,
            I => \N__28056\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__28077\,
            I => \N__28056\
        );

    \I__5756\ : Span4Mux_h
    port map (
            O => \N__28074\,
            I => \N__28053\
        );

    \I__5755\ : Span4Mux_h
    port map (
            O => \N__28071\,
            I => \N__28048\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__28068\,
            I => \N__28048\
        );

    \I__5753\ : Odrv12
    port map (
            O => \N__28063\,
            I => \b2v_inst11.count_clk_RNIZ0Z_3\
        );

    \I__5752\ : Odrv4
    port map (
            O => \N__28056\,
            I => \b2v_inst11.count_clk_RNIZ0Z_3\
        );

    \I__5751\ : Odrv4
    port map (
            O => \N__28053\,
            I => \b2v_inst11.count_clk_RNIZ0Z_3\
        );

    \I__5750\ : Odrv4
    port map (
            O => \N__28048\,
            I => \b2v_inst11.count_clk_RNIZ0Z_3\
        );

    \I__5749\ : CascadeMux
    port map (
            O => \N__28039\,
            I => \b2v_inst11.g1_2_1_cascade_\
        );

    \I__5748\ : CascadeMux
    port map (
            O => \N__28036\,
            I => \N__28033\
        );

    \I__5747\ : InMux
    port map (
            O => \N__28033\,
            I => \N__28025\
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__28032\,
            I => \N__28021\
        );

    \I__5745\ : InMux
    port map (
            O => \N__28031\,
            I => \N__28003\
        );

    \I__5744\ : InMux
    port map (
            O => \N__28030\,
            I => \N__28003\
        );

    \I__5743\ : InMux
    port map (
            O => \N__28029\,
            I => \N__28003\
        );

    \I__5742\ : CascadeMux
    port map (
            O => \N__28028\,
            I => \N__28000\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__28025\,
            I => \N__27996\
        );

    \I__5740\ : InMux
    port map (
            O => \N__28024\,
            I => \N__27991\
        );

    \I__5739\ : InMux
    port map (
            O => \N__28021\,
            I => \N__27991\
        );

    \I__5738\ : CascadeMux
    port map (
            O => \N__28020\,
            I => \N__27988\
        );

    \I__5737\ : InMux
    port map (
            O => \N__28019\,
            I => \N__27982\
        );

    \I__5736\ : InMux
    port map (
            O => \N__28018\,
            I => \N__27975\
        );

    \I__5735\ : InMux
    port map (
            O => \N__28017\,
            I => \N__27975\
        );

    \I__5734\ : InMux
    port map (
            O => \N__28016\,
            I => \N__27975\
        );

    \I__5733\ : InMux
    port map (
            O => \N__28015\,
            I => \N__27972\
        );

    \I__5732\ : InMux
    port map (
            O => \N__28014\,
            I => \N__27969\
        );

    \I__5731\ : CascadeMux
    port map (
            O => \N__28013\,
            I => \N__27966\
        );

    \I__5730\ : InMux
    port map (
            O => \N__28012\,
            I => \N__27958\
        );

    \I__5729\ : InMux
    port map (
            O => \N__28011\,
            I => \N__27958\
        );

    \I__5728\ : InMux
    port map (
            O => \N__28010\,
            I => \N__27958\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__28003\,
            I => \N__27953\
        );

    \I__5726\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27950\
        );

    \I__5725\ : InMux
    port map (
            O => \N__27999\,
            I => \N__27947\
        );

    \I__5724\ : Span4Mux_v
    port map (
            O => \N__27996\,
            I => \N__27942\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__27991\,
            I => \N__27942\
        );

    \I__5722\ : InMux
    port map (
            O => \N__27988\,
            I => \N__27939\
        );

    \I__5721\ : InMux
    port map (
            O => \N__27987\,
            I => \N__27936\
        );

    \I__5720\ : InMux
    port map (
            O => \N__27986\,
            I => \N__27931\
        );

    \I__5719\ : InMux
    port map (
            O => \N__27985\,
            I => \N__27931\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__27982\,
            I => \N__27928\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__27975\,
            I => \N__27921\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__27972\,
            I => \N__27921\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__27969\,
            I => \N__27921\
        );

    \I__5714\ : InMux
    port map (
            O => \N__27966\,
            I => \N__27916\
        );

    \I__5713\ : InMux
    port map (
            O => \N__27965\,
            I => \N__27916\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__27958\,
            I => \N__27913\
        );

    \I__5711\ : InMux
    port map (
            O => \N__27957\,
            I => \N__27909\
        );

    \I__5710\ : InMux
    port map (
            O => \N__27956\,
            I => \N__27906\
        );

    \I__5709\ : Span4Mux_v
    port map (
            O => \N__27953\,
            I => \N__27897\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__27950\,
            I => \N__27897\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__27947\,
            I => \N__27897\
        );

    \I__5706\ : Span4Mux_v
    port map (
            O => \N__27942\,
            I => \N__27897\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__27939\,
            I => \N__27890\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__27936\,
            I => \N__27890\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__27931\,
            I => \N__27890\
        );

    \I__5702\ : Span4Mux_v
    port map (
            O => \N__27928\,
            I => \N__27883\
        );

    \I__5701\ : Span4Mux_h
    port map (
            O => \N__27921\,
            I => \N__27883\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__27916\,
            I => \N__27883\
        );

    \I__5699\ : Span4Mux_h
    port map (
            O => \N__27913\,
            I => \N__27880\
        );

    \I__5698\ : InMux
    port map (
            O => \N__27912\,
            I => \N__27877\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__27909\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__27906\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__5695\ : Odrv4
    port map (
            O => \N__27897\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__5694\ : Odrv4
    port map (
            O => \N__27890\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__5693\ : Odrv4
    port map (
            O => \N__27883\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__5692\ : Odrv4
    port map (
            O => \N__27880\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__27877\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__5690\ : InMux
    port map (
            O => \N__27862\,
            I => \N__27859\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__27859\,
            I => \N__27856\
        );

    \I__5688\ : Odrv4
    port map (
            O => \N__27856\,
            I => \b2v_inst11.g1_2\
        );

    \I__5687\ : CascadeMux
    port map (
            O => \N__27853\,
            I => \b2v_inst6.countZ0Z_11_cascade_\
        );

    \I__5686\ : InMux
    port map (
            O => \N__27850\,
            I => \N__27847\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__27847\,
            I => \b2v_inst6.count_3_11\
        );

    \I__5684\ : CascadeMux
    port map (
            O => \N__27844\,
            I => \N__27840\
        );

    \I__5683\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27835\
        );

    \I__5682\ : InMux
    port map (
            O => \N__27840\,
            I => \N__27835\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__27835\,
            I => \b2v_inst6.curr_state_RNIDMSJ1Z0Z_1\
        );

    \I__5680\ : InMux
    port map (
            O => \N__27832\,
            I => \N__27829\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__27829\,
            I => b2v_inst11_count_off_1_sqmuxa_0_0_0
        );

    \I__5678\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27823\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__27823\,
            I => \G_26_0_a5_1_0\
        );

    \I__5676\ : CascadeMux
    port map (
            O => \N__27820\,
            I => \G_26_0_a5_2_1_cascade_\
        );

    \I__5675\ : InMux
    port map (
            O => \N__27817\,
            I => \N__27814\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__27814\,
            I => \G_26_0_0\
        );

    \I__5673\ : InMux
    port map (
            O => \N__27811\,
            I => \N__27808\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__27808\,
            I => \N__27805\
        );

    \I__5671\ : Span4Mux_h
    port map (
            O => \N__27805\,
            I => \N__27802\
        );

    \I__5670\ : Odrv4
    port map (
            O => \N__27802\,
            I => \b2v_inst11.g2_0_1\
        );

    \I__5669\ : InMux
    port map (
            O => \N__27799\,
            I => \N__27796\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__27796\,
            I => \b2v_inst11.un1_dutycycle_172_m4\
        );

    \I__5667\ : CascadeMux
    port map (
            O => \N__27793\,
            I => \b2v_inst11_un1_dutycycle_172_m3_0_0_0_cascade_\
        );

    \I__5666\ : InMux
    port map (
            O => \N__27790\,
            I => \N__27787\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__27787\,
            I => \N__27784\
        );

    \I__5664\ : Odrv4
    port map (
            O => \N__27784\,
            I => \b2v_inst11.g2_1\
        );

    \I__5663\ : CascadeMux
    port map (
            O => \N__27781\,
            I => \N__27773\
        );

    \I__5662\ : InMux
    port map (
            O => \N__27780\,
            I => \N__27767\
        );

    \I__5661\ : InMux
    port map (
            O => \N__27779\,
            I => \N__27764\
        );

    \I__5660\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27761\
        );

    \I__5659\ : InMux
    port map (
            O => \N__27777\,
            I => \N__27755\
        );

    \I__5658\ : InMux
    port map (
            O => \N__27776\,
            I => \N__27747\
        );

    \I__5657\ : InMux
    port map (
            O => \N__27773\,
            I => \N__27742\
        );

    \I__5656\ : InMux
    port map (
            O => \N__27772\,
            I => \N__27742\
        );

    \I__5655\ : InMux
    port map (
            O => \N__27771\,
            I => \N__27738\
        );

    \I__5654\ : InMux
    port map (
            O => \N__27770\,
            I => \N__27735\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__27767\,
            I => \N__27728\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__27764\,
            I => \N__27728\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__27761\,
            I => \N__27728\
        );

    \I__5650\ : InMux
    port map (
            O => \N__27760\,
            I => \N__27721\
        );

    \I__5649\ : InMux
    port map (
            O => \N__27759\,
            I => \N__27721\
        );

    \I__5648\ : InMux
    port map (
            O => \N__27758\,
            I => \N__27721\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__27755\,
            I => \N__27718\
        );

    \I__5646\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27715\
        );

    \I__5645\ : InMux
    port map (
            O => \N__27753\,
            I => \N__27710\
        );

    \I__5644\ : InMux
    port map (
            O => \N__27752\,
            I => \N__27710\
        );

    \I__5643\ : InMux
    port map (
            O => \N__27751\,
            I => \N__27707\
        );

    \I__5642\ : InMux
    port map (
            O => \N__27750\,
            I => \N__27704\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__27747\,
            I => \N__27699\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__27742\,
            I => \N__27699\
        );

    \I__5639\ : CascadeMux
    port map (
            O => \N__27741\,
            I => \N__27696\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__27738\,
            I => \N__27689\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__27735\,
            I => \N__27686\
        );

    \I__5636\ : Span4Mux_v
    port map (
            O => \N__27728\,
            I => \N__27681\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__27721\,
            I => \N__27681\
        );

    \I__5634\ : Span4Mux_h
    port map (
            O => \N__27718\,
            I => \N__27676\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__27715\,
            I => \N__27676\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__27710\,
            I => \N__27667\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__27707\,
            I => \N__27667\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__27704\,
            I => \N__27667\
        );

    \I__5629\ : Span4Mux_s2_v
    port map (
            O => \N__27699\,
            I => \N__27667\
        );

    \I__5628\ : InMux
    port map (
            O => \N__27696\,
            I => \N__27664\
        );

    \I__5627\ : InMux
    port map (
            O => \N__27695\,
            I => \N__27661\
        );

    \I__5626\ : InMux
    port map (
            O => \N__27694\,
            I => \N__27654\
        );

    \I__5625\ : InMux
    port map (
            O => \N__27693\,
            I => \N__27654\
        );

    \I__5624\ : InMux
    port map (
            O => \N__27692\,
            I => \N__27654\
        );

    \I__5623\ : Span4Mux_s3_v
    port map (
            O => \N__27689\,
            I => \N__27645\
        );

    \I__5622\ : Span4Mux_s3_v
    port map (
            O => \N__27686\,
            I => \N__27645\
        );

    \I__5621\ : Span4Mux_h
    port map (
            O => \N__27681\,
            I => \N__27645\
        );

    \I__5620\ : Span4Mux_h
    port map (
            O => \N__27676\,
            I => \N__27645\
        );

    \I__5619\ : Span4Mux_v
    port map (
            O => \N__27667\,
            I => \N__27642\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__27664\,
            I => \N__27637\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__27661\,
            I => \N__27637\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__27654\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z2\
        );

    \I__5615\ : Odrv4
    port map (
            O => \N__27645\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z2\
        );

    \I__5614\ : Odrv4
    port map (
            O => \N__27642\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z2\
        );

    \I__5613\ : Odrv4
    port map (
            O => \N__27637\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z2\
        );

    \I__5612\ : CascadeMux
    port map (
            O => \N__27628\,
            I => \b2v_inst11.g4_cascade_\
        );

    \I__5611\ : IoInMux
    port map (
            O => \N__27625\,
            I => \N__27621\
        );

    \I__5610\ : InMux
    port map (
            O => \N__27624\,
            I => \N__27614\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__27621\,
            I => \N__27611\
        );

    \I__5608\ : CascadeMux
    port map (
            O => \N__27620\,
            I => \N__27607\
        );

    \I__5607\ : InMux
    port map (
            O => \N__27619\,
            I => \N__27600\
        );

    \I__5606\ : InMux
    port map (
            O => \N__27618\,
            I => \N__27588\
        );

    \I__5605\ : InMux
    port map (
            O => \N__27617\,
            I => \N__27588\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__27614\,
            I => \N__27582\
        );

    \I__5603\ : IoSpan4Mux
    port map (
            O => \N__27611\,
            I => \N__27582\
        );

    \I__5602\ : InMux
    port map (
            O => \N__27610\,
            I => \N__27575\
        );

    \I__5601\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27575\
        );

    \I__5600\ : InMux
    port map (
            O => \N__27606\,
            I => \N__27575\
        );

    \I__5599\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27570\
        );

    \I__5598\ : InMux
    port map (
            O => \N__27604\,
            I => \N__27570\
        );

    \I__5597\ : InMux
    port map (
            O => \N__27603\,
            I => \N__27567\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__27600\,
            I => \N__27564\
        );

    \I__5595\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27561\
        );

    \I__5594\ : InMux
    port map (
            O => \N__27598\,
            I => \N__27558\
        );

    \I__5593\ : InMux
    port map (
            O => \N__27597\,
            I => \N__27551\
        );

    \I__5592\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27551\
        );

    \I__5591\ : InMux
    port map (
            O => \N__27595\,
            I => \N__27551\
        );

    \I__5590\ : InMux
    port map (
            O => \N__27594\,
            I => \N__27540\
        );

    \I__5589\ : InMux
    port map (
            O => \N__27593\,
            I => \N__27540\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__27588\,
            I => \N__27537\
        );

    \I__5587\ : InMux
    port map (
            O => \N__27587\,
            I => \N__27532\
        );

    \I__5586\ : Span4Mux_s3_v
    port map (
            O => \N__27582\,
            I => \N__27529\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__27575\,
            I => \N__27524\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__27570\,
            I => \N__27524\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__27567\,
            I => \N__27521\
        );

    \I__5582\ : Span4Mux_s3_v
    port map (
            O => \N__27564\,
            I => \N__27514\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__27561\,
            I => \N__27514\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__27558\,
            I => \N__27514\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__27551\,
            I => \N__27511\
        );

    \I__5578\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27504\
        );

    \I__5577\ : InMux
    port map (
            O => \N__27549\,
            I => \N__27504\
        );

    \I__5576\ : InMux
    port map (
            O => \N__27548\,
            I => \N__27504\
        );

    \I__5575\ : InMux
    port map (
            O => \N__27547\,
            I => \N__27499\
        );

    \I__5574\ : InMux
    port map (
            O => \N__27546\,
            I => \N__27499\
        );

    \I__5573\ : InMux
    port map (
            O => \N__27545\,
            I => \N__27496\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__27540\,
            I => \N__27493\
        );

    \I__5571\ : Span4Mux_h
    port map (
            O => \N__27537\,
            I => \N__27490\
        );

    \I__5570\ : InMux
    port map (
            O => \N__27536\,
            I => \N__27485\
        );

    \I__5569\ : InMux
    port map (
            O => \N__27535\,
            I => \N__27485\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__27532\,
            I => \N__27482\
        );

    \I__5567\ : Span4Mux_h
    port map (
            O => \N__27529\,
            I => \N__27467\
        );

    \I__5566\ : Span4Mux_s3_v
    port map (
            O => \N__27524\,
            I => \N__27467\
        );

    \I__5565\ : Span4Mux_s3_v
    port map (
            O => \N__27521\,
            I => \N__27467\
        );

    \I__5564\ : Span4Mux_h
    port map (
            O => \N__27514\,
            I => \N__27467\
        );

    \I__5563\ : Span4Mux_h
    port map (
            O => \N__27511\,
            I => \N__27467\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__27504\,
            I => \N__27467\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__27499\,
            I => \N__27467\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__27496\,
            I => \N__27464\
        );

    \I__5559\ : Odrv4
    port map (
            O => \N__27493\,
            I => b2v_inst16_delayed_vddq_pwrgd_en
        );

    \I__5558\ : Odrv4
    port map (
            O => \N__27490\,
            I => b2v_inst16_delayed_vddq_pwrgd_en
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__27485\,
            I => b2v_inst16_delayed_vddq_pwrgd_en
        );

    \I__5556\ : Odrv12
    port map (
            O => \N__27482\,
            I => b2v_inst16_delayed_vddq_pwrgd_en
        );

    \I__5555\ : Odrv4
    port map (
            O => \N__27467\,
            I => b2v_inst16_delayed_vddq_pwrgd_en
        );

    \I__5554\ : Odrv4
    port map (
            O => \N__27464\,
            I => b2v_inst16_delayed_vddq_pwrgd_en
        );

    \I__5553\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27445\
        );

    \I__5552\ : InMux
    port map (
            O => \N__27450\,
            I => \N__27445\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__27445\,
            I => \b2v_inst11.N_5\
        );

    \I__5550\ : InMux
    port map (
            O => \N__27442\,
            I => \N__27439\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__27439\,
            I => \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_xZ0\
        );

    \I__5548\ : CascadeMux
    port map (
            O => \N__27436\,
            I => \N__27432\
        );

    \I__5547\ : CascadeMux
    port map (
            O => \N__27435\,
            I => \N__27429\
        );

    \I__5546\ : InMux
    port map (
            O => \N__27432\,
            I => \N__27423\
        );

    \I__5545\ : InMux
    port map (
            O => \N__27429\,
            I => \N__27418\
        );

    \I__5544\ : InMux
    port map (
            O => \N__27428\,
            I => \N__27418\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__27427\,
            I => \N__27414\
        );

    \I__5542\ : InMux
    port map (
            O => \N__27426\,
            I => \N__27410\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__27423\,
            I => \N__27403\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__27418\,
            I => \N__27403\
        );

    \I__5539\ : InMux
    port map (
            O => \N__27417\,
            I => \N__27400\
        );

    \I__5538\ : InMux
    port map (
            O => \N__27414\,
            I => \N__27397\
        );

    \I__5537\ : CascadeMux
    port map (
            O => \N__27413\,
            I => \N__27394\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__27410\,
            I => \N__27391\
        );

    \I__5535\ : InMux
    port map (
            O => \N__27409\,
            I => \N__27386\
        );

    \I__5534\ : InMux
    port map (
            O => \N__27408\,
            I => \N__27383\
        );

    \I__5533\ : Span4Mux_v
    port map (
            O => \N__27403\,
            I => \N__27379\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__27400\,
            I => \N__27374\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__27397\,
            I => \N__27374\
        );

    \I__5530\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27371\
        );

    \I__5529\ : Span12Mux_v
    port map (
            O => \N__27391\,
            I => \N__27368\
        );

    \I__5528\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27365\
        );

    \I__5527\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27362\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__27386\,
            I => \N__27359\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__27383\,
            I => \N__27356\
        );

    \I__5524\ : InMux
    port map (
            O => \N__27382\,
            I => \N__27353\
        );

    \I__5523\ : Span4Mux_v
    port map (
            O => \N__27379\,
            I => \N__27346\
        );

    \I__5522\ : Span4Mux_s3_v
    port map (
            O => \N__27374\,
            I => \N__27346\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__27371\,
            I => \N__27346\
        );

    \I__5520\ : Odrv12
    port map (
            O => \N__27368\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__27365\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__27362\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__5517\ : Odrv4
    port map (
            O => \N__27359\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__5516\ : Odrv4
    port map (
            O => \N__27356\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__27353\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__5514\ : Odrv4
    port map (
            O => \N__27346\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__5513\ : InMux
    port map (
            O => \N__27331\,
            I => \N__27325\
        );

    \I__5512\ : InMux
    port map (
            O => \N__27330\,
            I => \N__27325\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__27325\,
            I => \b2v_inst11.N_12\
        );

    \I__5510\ : CascadeMux
    port map (
            O => \N__27322\,
            I => \N__27319\
        );

    \I__5509\ : InMux
    port map (
            O => \N__27319\,
            I => \N__27308\
        );

    \I__5508\ : InMux
    port map (
            O => \N__27318\,
            I => \N__27297\
        );

    \I__5507\ : InMux
    port map (
            O => \N__27317\,
            I => \N__27297\
        );

    \I__5506\ : InMux
    port map (
            O => \N__27316\,
            I => \N__27289\
        );

    \I__5505\ : InMux
    port map (
            O => \N__27315\,
            I => \N__27284\
        );

    \I__5504\ : InMux
    port map (
            O => \N__27314\,
            I => \N__27284\
        );

    \I__5503\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27279\
        );

    \I__5502\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27279\
        );

    \I__5501\ : InMux
    port map (
            O => \N__27311\,
            I => \N__27276\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__27308\,
            I => \N__27271\
        );

    \I__5499\ : InMux
    port map (
            O => \N__27307\,
            I => \N__27266\
        );

    \I__5498\ : InMux
    port map (
            O => \N__27306\,
            I => \N__27266\
        );

    \I__5497\ : InMux
    port map (
            O => \N__27305\,
            I => \N__27263\
        );

    \I__5496\ : InMux
    port map (
            O => \N__27304\,
            I => \N__27259\
        );

    \I__5495\ : InMux
    port map (
            O => \N__27303\,
            I => \N__27252\
        );

    \I__5494\ : InMux
    port map (
            O => \N__27302\,
            I => \N__27252\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__27297\,
            I => \N__27249\
        );

    \I__5492\ : InMux
    port map (
            O => \N__27296\,
            I => \N__27240\
        );

    \I__5491\ : InMux
    port map (
            O => \N__27295\,
            I => \N__27240\
        );

    \I__5490\ : InMux
    port map (
            O => \N__27294\,
            I => \N__27240\
        );

    \I__5489\ : InMux
    port map (
            O => \N__27293\,
            I => \N__27240\
        );

    \I__5488\ : InMux
    port map (
            O => \N__27292\,
            I => \N__27237\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__27289\,
            I => \N__27221\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__27284\,
            I => \N__27221\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__27279\,
            I => \N__27221\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__27276\,
            I => \N__27218\
        );

    \I__5483\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27213\
        );

    \I__5482\ : InMux
    port map (
            O => \N__27274\,
            I => \N__27213\
        );

    \I__5481\ : Span4Mux_v
    port map (
            O => \N__27271\,
            I => \N__27206\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__27266\,
            I => \N__27206\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__27263\,
            I => \N__27206\
        );

    \I__5478\ : InMux
    port map (
            O => \N__27262\,
            I => \N__27203\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__27259\,
            I => \N__27200\
        );

    \I__5476\ : InMux
    port map (
            O => \N__27258\,
            I => \N__27195\
        );

    \I__5475\ : InMux
    port map (
            O => \N__27257\,
            I => \N__27195\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__27252\,
            I => \N__27188\
        );

    \I__5473\ : Span4Mux_v
    port map (
            O => \N__27249\,
            I => \N__27188\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__27240\,
            I => \N__27188\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__27237\,
            I => \N__27185\
        );

    \I__5470\ : InMux
    port map (
            O => \N__27236\,
            I => \N__27182\
        );

    \I__5469\ : InMux
    port map (
            O => \N__27235\,
            I => \N__27179\
        );

    \I__5468\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27168\
        );

    \I__5467\ : InMux
    port map (
            O => \N__27233\,
            I => \N__27168\
        );

    \I__5466\ : InMux
    port map (
            O => \N__27232\,
            I => \N__27168\
        );

    \I__5465\ : InMux
    port map (
            O => \N__27231\,
            I => \N__27168\
        );

    \I__5464\ : InMux
    port map (
            O => \N__27230\,
            I => \N__27168\
        );

    \I__5463\ : InMux
    port map (
            O => \N__27229\,
            I => \N__27163\
        );

    \I__5462\ : InMux
    port map (
            O => \N__27228\,
            I => \N__27163\
        );

    \I__5461\ : Span4Mux_v
    port map (
            O => \N__27221\,
            I => \N__27160\
        );

    \I__5460\ : Span4Mux_v
    port map (
            O => \N__27218\,
            I => \N__27153\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__27213\,
            I => \N__27153\
        );

    \I__5458\ : Span4Mux_v
    port map (
            O => \N__27206\,
            I => \N__27153\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__27203\,
            I => \N__27148\
        );

    \I__5456\ : Span4Mux_h
    port map (
            O => \N__27200\,
            I => \N__27148\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__27195\,
            I => \N__27141\
        );

    \I__5454\ : Span4Mux_h
    port map (
            O => \N__27188\,
            I => \N__27141\
        );

    \I__5453\ : Span4Mux_h
    port map (
            O => \N__27185\,
            I => \N__27141\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__27182\,
            I => \b2v_inst11.func_state_RNINJ641_0Z0Z_1\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__27179\,
            I => \b2v_inst11.func_state_RNINJ641_0Z0Z_1\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__27168\,
            I => \b2v_inst11.func_state_RNINJ641_0Z0Z_1\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__27163\,
            I => \b2v_inst11.func_state_RNINJ641_0Z0Z_1\
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__27160\,
            I => \b2v_inst11.func_state_RNINJ641_0Z0Z_1\
        );

    \I__5447\ : Odrv4
    port map (
            O => \N__27153\,
            I => \b2v_inst11.func_state_RNINJ641_0Z0Z_1\
        );

    \I__5446\ : Odrv4
    port map (
            O => \N__27148\,
            I => \b2v_inst11.func_state_RNINJ641_0Z0Z_1\
        );

    \I__5445\ : Odrv4
    port map (
            O => \N__27141\,
            I => \b2v_inst11.func_state_RNINJ641_0Z0Z_1\
        );

    \I__5444\ : InMux
    port map (
            O => \N__27124\,
            I => \N__27121\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__27121\,
            I => \N_4\
        );

    \I__5442\ : InMux
    port map (
            O => \N__27118\,
            I => \N__27115\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__27115\,
            I => \N__27112\
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__27112\,
            I => \G_26_0_a5_2\
        );

    \I__5439\ : CascadeMux
    port map (
            O => \N__27109\,
            I => \N__27104\
        );

    \I__5438\ : InMux
    port map (
            O => \N__27108\,
            I => \N__27098\
        );

    \I__5437\ : InMux
    port map (
            O => \N__27107\,
            I => \N__27098\
        );

    \I__5436\ : InMux
    port map (
            O => \N__27104\,
            I => \N__27093\
        );

    \I__5435\ : InMux
    port map (
            O => \N__27103\,
            I => \N__27093\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__27098\,
            I => \N__27084\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__27093\,
            I => \N__27081\
        );

    \I__5432\ : InMux
    port map (
            O => \N__27092\,
            I => \N__27078\
        );

    \I__5431\ : InMux
    port map (
            O => \N__27091\,
            I => \N__27075\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__27090\,
            I => \N__27072\
        );

    \I__5429\ : InMux
    port map (
            O => \N__27089\,
            I => \N__27065\
        );

    \I__5428\ : InMux
    port map (
            O => \N__27088\,
            I => \N__27065\
        );

    \I__5427\ : InMux
    port map (
            O => \N__27087\,
            I => \N__27062\
        );

    \I__5426\ : Span4Mux_v
    port map (
            O => \N__27084\,
            I => \N__27053\
        );

    \I__5425\ : Span4Mux_h
    port map (
            O => \N__27081\,
            I => \N__27053\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__27078\,
            I => \N__27053\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__27075\,
            I => \N__27053\
        );

    \I__5422\ : InMux
    port map (
            O => \N__27072\,
            I => \N__27050\
        );

    \I__5421\ : InMux
    port map (
            O => \N__27071\,
            I => \N__27045\
        );

    \I__5420\ : InMux
    port map (
            O => \N__27070\,
            I => \N__27045\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__27065\,
            I => \curr_state_RNI5VS71_0_1\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__27062\,
            I => \curr_state_RNI5VS71_0_1\
        );

    \I__5417\ : Odrv4
    port map (
            O => \N__27053\,
            I => \curr_state_RNI5VS71_0_1\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__27050\,
            I => \curr_state_RNI5VS71_0_1\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__27045\,
            I => \curr_state_RNI5VS71_0_1\
        );

    \I__5414\ : InMux
    port map (
            O => \N__27034\,
            I => \N__27031\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__27031\,
            I => \N__27022\
        );

    \I__5412\ : InMux
    port map (
            O => \N__27030\,
            I => \N__27016\
        );

    \I__5411\ : InMux
    port map (
            O => \N__27029\,
            I => \N__27016\
        );

    \I__5410\ : InMux
    port map (
            O => \N__27028\,
            I => \N__27013\
        );

    \I__5409\ : InMux
    port map (
            O => \N__27027\,
            I => \N__27008\
        );

    \I__5408\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27008\
        );

    \I__5407\ : CascadeMux
    port map (
            O => \N__27025\,
            I => \N__27005\
        );

    \I__5406\ : Span12Mux_s7_v
    port map (
            O => \N__27022\,
            I => \N__27001\
        );

    \I__5405\ : InMux
    port map (
            O => \N__27021\,
            I => \N__26998\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__27016\,
            I => \N__26995\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__27013\,
            I => \N__26990\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__27008\,
            I => \N__26990\
        );

    \I__5401\ : InMux
    port map (
            O => \N__27005\,
            I => \N__26987\
        );

    \I__5400\ : InMux
    port map (
            O => \N__27004\,
            I => \N__26984\
        );

    \I__5399\ : Odrv12
    port map (
            O => \N__27001\,
            I => \RSMRSTn_0\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__26998\,
            I => \RSMRSTn_0\
        );

    \I__5397\ : Odrv4
    port map (
            O => \N__26995\,
            I => \RSMRSTn_0\
        );

    \I__5396\ : Odrv12
    port map (
            O => \N__26990\,
            I => \RSMRSTn_0\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__26987\,
            I => \RSMRSTn_0\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__26984\,
            I => \RSMRSTn_0\
        );

    \I__5393\ : CascadeMux
    port map (
            O => \N__26971\,
            I => \b2v_inst11.N_234_cascade_\
        );

    \I__5392\ : CascadeMux
    port map (
            O => \N__26968\,
            I => \b2v_inst11.un1_clk_100khz_52_and_i_0_0_cascade_\
        );

    \I__5391\ : CascadeMux
    port map (
            O => \N__26965\,
            I => \N__26961\
        );

    \I__5390\ : InMux
    port map (
            O => \N__26964\,
            I => \N__26956\
        );

    \I__5389\ : InMux
    port map (
            O => \N__26961\,
            I => \N__26951\
        );

    \I__5388\ : InMux
    port map (
            O => \N__26960\,
            I => \N__26946\
        );

    \I__5387\ : InMux
    port map (
            O => \N__26959\,
            I => \N__26946\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__26956\,
            I => \N__26943\
        );

    \I__5385\ : InMux
    port map (
            O => \N__26955\,
            I => \N__26937\
        );

    \I__5384\ : InMux
    port map (
            O => \N__26954\,
            I => \N__26937\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__26951\,
            I => \N__26934\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__26946\,
            I => \N__26931\
        );

    \I__5381\ : Span4Mux_v
    port map (
            O => \N__26943\,
            I => \N__26928\
        );

    \I__5380\ : InMux
    port map (
            O => \N__26942\,
            I => \N__26920\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__26937\,
            I => \N__26917\
        );

    \I__5378\ : Span4Mux_v
    port map (
            O => \N__26934\,
            I => \N__26912\
        );

    \I__5377\ : Span4Mux_v
    port map (
            O => \N__26931\,
            I => \N__26912\
        );

    \I__5376\ : Span4Mux_h
    port map (
            O => \N__26928\,
            I => \N__26909\
        );

    \I__5375\ : InMux
    port map (
            O => \N__26927\,
            I => \N__26906\
        );

    \I__5374\ : InMux
    port map (
            O => \N__26926\,
            I => \N__26899\
        );

    \I__5373\ : InMux
    port map (
            O => \N__26925\,
            I => \N__26899\
        );

    \I__5372\ : InMux
    port map (
            O => \N__26924\,
            I => \N__26899\
        );

    \I__5371\ : InMux
    port map (
            O => \N__26923\,
            I => \N__26896\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__26920\,
            I => \SYNTHESIZED_WIRE_47keep_rep1\
        );

    \I__5369\ : Odrv12
    port map (
            O => \N__26917\,
            I => \SYNTHESIZED_WIRE_47keep_rep1\
        );

    \I__5368\ : Odrv4
    port map (
            O => \N__26912\,
            I => \SYNTHESIZED_WIRE_47keep_rep1\
        );

    \I__5367\ : Odrv4
    port map (
            O => \N__26909\,
            I => \SYNTHESIZED_WIRE_47keep_rep1\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__26906\,
            I => \SYNTHESIZED_WIRE_47keep_rep1\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__26899\,
            I => \SYNTHESIZED_WIRE_47keep_rep1\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__26896\,
            I => \SYNTHESIZED_WIRE_47keep_rep1\
        );

    \I__5363\ : CascadeMux
    port map (
            O => \N__26881\,
            I => \N__26874\
        );

    \I__5362\ : InMux
    port map (
            O => \N__26880\,
            I => \N__26868\
        );

    \I__5361\ : InMux
    port map (
            O => \N__26879\,
            I => \N__26868\
        );

    \I__5360\ : InMux
    port map (
            O => \N__26878\,
            I => \N__26863\
        );

    \I__5359\ : InMux
    port map (
            O => \N__26877\,
            I => \N__26860\
        );

    \I__5358\ : InMux
    port map (
            O => \N__26874\,
            I => \N__26855\
        );

    \I__5357\ : InMux
    port map (
            O => \N__26873\,
            I => \N__26855\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__26868\,
            I => \N__26852\
        );

    \I__5355\ : CascadeMux
    port map (
            O => \N__26867\,
            I => \N__26845\
        );

    \I__5354\ : InMux
    port map (
            O => \N__26866\,
            I => \N__26840\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__26863\,
            I => \N__26837\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__26860\,
            I => \N__26834\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__26855\,
            I => \N__26831\
        );

    \I__5350\ : Span4Mux_h
    port map (
            O => \N__26852\,
            I => \N__26828\
        );

    \I__5349\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26822\
        );

    \I__5348\ : InMux
    port map (
            O => \N__26850\,
            I => \N__26822\
        );

    \I__5347\ : InMux
    port map (
            O => \N__26849\,
            I => \N__26811\
        );

    \I__5346\ : InMux
    port map (
            O => \N__26848\,
            I => \N__26811\
        );

    \I__5345\ : InMux
    port map (
            O => \N__26845\,
            I => \N__26811\
        );

    \I__5344\ : InMux
    port map (
            O => \N__26844\,
            I => \N__26811\
        );

    \I__5343\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26811\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__26840\,
            I => \N__26806\
        );

    \I__5341\ : Span4Mux_v
    port map (
            O => \N__26837\,
            I => \N__26806\
        );

    \I__5340\ : Span4Mux_v
    port map (
            O => \N__26834\,
            I => \N__26801\
        );

    \I__5339\ : Span4Mux_h
    port map (
            O => \N__26831\,
            I => \N__26801\
        );

    \I__5338\ : Span4Mux_h
    port map (
            O => \N__26828\,
            I => \N__26798\
        );

    \I__5337\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26795\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__26822\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__26811\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__5334\ : Odrv4
    port map (
            O => \N__26806\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__5333\ : Odrv4
    port map (
            O => \N__26801\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__5332\ : Odrv4
    port map (
            O => \N__26798\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__26795\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__5330\ : CascadeMux
    port map (
            O => \N__26782\,
            I => \N__26776\
        );

    \I__5329\ : CascadeMux
    port map (
            O => \N__26781\,
            I => \N__26773\
        );

    \I__5328\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26770\
        );

    \I__5327\ : CascadeMux
    port map (
            O => \N__26779\,
            I => \N__26767\
        );

    \I__5326\ : InMux
    port map (
            O => \N__26776\,
            I => \N__26761\
        );

    \I__5325\ : InMux
    port map (
            O => \N__26773\,
            I => \N__26758\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__26770\,
            I => \N__26754\
        );

    \I__5323\ : InMux
    port map (
            O => \N__26767\,
            I => \N__26749\
        );

    \I__5322\ : InMux
    port map (
            O => \N__26766\,
            I => \N__26749\
        );

    \I__5321\ : InMux
    port map (
            O => \N__26765\,
            I => \N__26746\
        );

    \I__5320\ : CascadeMux
    port map (
            O => \N__26764\,
            I => \N__26743\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__26761\,
            I => \N__26739\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__26758\,
            I => \N__26736\
        );

    \I__5317\ : CascadeMux
    port map (
            O => \N__26757\,
            I => \N__26733\
        );

    \I__5316\ : Span4Mux_h
    port map (
            O => \N__26754\,
            I => \N__26729\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__26749\,
            I => \N__26724\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__26746\,
            I => \N__26724\
        );

    \I__5313\ : InMux
    port map (
            O => \N__26743\,
            I => \N__26721\
        );

    \I__5312\ : InMux
    port map (
            O => \N__26742\,
            I => \N__26718\
        );

    \I__5311\ : Span4Mux_v
    port map (
            O => \N__26739\,
            I => \N__26713\
        );

    \I__5310\ : Span4Mux_v
    port map (
            O => \N__26736\,
            I => \N__26713\
        );

    \I__5309\ : InMux
    port map (
            O => \N__26733\,
            I => \N__26708\
        );

    \I__5308\ : InMux
    port map (
            O => \N__26732\,
            I => \N__26708\
        );

    \I__5307\ : Span4Mux_v
    port map (
            O => \N__26729\,
            I => \N__26703\
        );

    \I__5306\ : Span4Mux_h
    port map (
            O => \N__26724\,
            I => \N__26703\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__26721\,
            I => \dutycycle_RNIIOE3D_0_5\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__26718\,
            I => \dutycycle_RNIIOE3D_0_5\
        );

    \I__5303\ : Odrv4
    port map (
            O => \N__26713\,
            I => \dutycycle_RNIIOE3D_0_5\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__26708\,
            I => \dutycycle_RNIIOE3D_0_5\
        );

    \I__5301\ : Odrv4
    port map (
            O => \N__26703\,
            I => \dutycycle_RNIIOE3D_0_5\
        );

    \I__5300\ : InMux
    port map (
            O => \N__26692\,
            I => \bfn_9_10_0_\
        );

    \I__5299\ : CascadeMux
    port map (
            O => \N__26689\,
            I => \N__26686\
        );

    \I__5298\ : InMux
    port map (
            O => \N__26686\,
            I => \N__26683\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__26683\,
            I => \b2v_inst20.un4_counter_1_and\
        );

    \I__5296\ : InMux
    port map (
            O => \N__26680\,
            I => \N__26677\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__26677\,
            I => \N__26674\
        );

    \I__5294\ : Span4Mux_v
    port map (
            O => \N__26674\,
            I => \N__26671\
        );

    \I__5293\ : Odrv4
    port map (
            O => \N__26671\,
            I => \b2v_inst11.dutycycle_RNITBKN1Z0Z_7\
        );

    \I__5292\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26664\
        );

    \I__5291\ : InMux
    port map (
            O => \N__26667\,
            I => \N__26661\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__26664\,
            I => \N_229\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__26661\,
            I => \N_229\
        );

    \I__5288\ : CascadeMux
    port map (
            O => \N__26656\,
            I => \b2v_inst5.count_enZ0_cascade_\
        );

    \I__5287\ : CascadeMux
    port map (
            O => \N__26653\,
            I => \N__26650\
        );

    \I__5286\ : InMux
    port map (
            O => \N__26650\,
            I => \N__26646\
        );

    \I__5285\ : CascadeMux
    port map (
            O => \N__26649\,
            I => \N__26643\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__26646\,
            I => \N__26639\
        );

    \I__5283\ : InMux
    port map (
            O => \N__26643\,
            I => \N__26633\
        );

    \I__5282\ : InMux
    port map (
            O => \N__26642\,
            I => \N__26633\
        );

    \I__5281\ : Span4Mux_h
    port map (
            O => \N__26639\,
            I => \N__26630\
        );

    \I__5280\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26627\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__26633\,
            I => \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__5278\ : Odrv4
    port map (
            O => \N__26630\,
            I => \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__26627\,
            I => \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__5276\ : InMux
    port map (
            O => \N__26620\,
            I => \N__26617\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__26617\,
            I => \N__26614\
        );

    \I__5274\ : Odrv4
    port map (
            O => \N__26614\,
            I => \b2v_inst11.g0_2_1\
        );

    \I__5273\ : InMux
    port map (
            O => \N__26611\,
            I => \N__26607\
        );

    \I__5272\ : InMux
    port map (
            O => \N__26610\,
            I => \N__26603\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__26607\,
            I => \N__26600\
        );

    \I__5270\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26597\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__26603\,
            I => \N__26594\
        );

    \I__5268\ : Odrv4
    port map (
            O => \N__26600\,
            I => \b2v_inst11.pwm_outZ0\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__26597\,
            I => \b2v_inst11.pwm_outZ0\
        );

    \I__5266\ : Odrv4
    port map (
            O => \N__26594\,
            I => \b2v_inst11.pwm_outZ0\
        );

    \I__5265\ : SRMux
    port map (
            O => \N__26587\,
            I => \N__26584\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__26584\,
            I => \N__26581\
        );

    \I__5263\ : Span4Mux_v
    port map (
            O => \N__26581\,
            I => \N__26578\
        );

    \I__5262\ : Odrv4
    port map (
            O => \N__26578\,
            I => \b2v_inst11.pwm_out_1_sqmuxa\
        );

    \I__5261\ : CascadeMux
    port map (
            O => \N__26575\,
            I => \N__26572\
        );

    \I__5260\ : InMux
    port map (
            O => \N__26572\,
            I => \N__26569\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__26569\,
            I => \b2v_inst20.un4_counter_0_and\
        );

    \I__5258\ : CascadeMux
    port map (
            O => \N__26566\,
            I => \b2v_inst11.count_RNIZ0Z_1_cascade_\
        );

    \I__5257\ : InMux
    port map (
            O => \N__26563\,
            I => \N__26560\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__26560\,
            I => \N__26556\
        );

    \I__5255\ : CascadeMux
    port map (
            O => \N__26559\,
            I => \N__26552\
        );

    \I__5254\ : Span12Mux_s8_h
    port map (
            O => \N__26556\,
            I => \N__26549\
        );

    \I__5253\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26546\
        );

    \I__5252\ : InMux
    port map (
            O => \N__26552\,
            I => \N__26543\
        );

    \I__5251\ : Odrv12
    port map (
            O => \N__26549\,
            I => \b2v_inst11.countZ0Z_1\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__26546\,
            I => \b2v_inst11.countZ0Z_1\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__26543\,
            I => \b2v_inst11.countZ0Z_1\
        );

    \I__5248\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26532\
        );

    \I__5247\ : InMux
    port map (
            O => \N__26535\,
            I => \N__26528\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__26532\,
            I => \N__26525\
        );

    \I__5245\ : InMux
    port map (
            O => \N__26531\,
            I => \N__26522\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__26528\,
            I => \N__26519\
        );

    \I__5243\ : Span4Mux_v
    port map (
            O => \N__26525\,
            I => \N__26512\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__26522\,
            I => \N__26512\
        );

    \I__5241\ : Span4Mux_h
    port map (
            O => \N__26519\,
            I => \N__26509\
        );

    \I__5240\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26506\
        );

    \I__5239\ : InMux
    port map (
            O => \N__26517\,
            I => \N__26503\
        );

    \I__5238\ : Odrv4
    port map (
            O => \N__26512\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__5237\ : Odrv4
    port map (
            O => \N__26509\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__26506\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__26503\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__5234\ : CascadeMux
    port map (
            O => \N__26494\,
            I => \b2v_inst11.countZ0Z_1_cascade_\
        );

    \I__5233\ : InMux
    port map (
            O => \N__26491\,
            I => \N__26470\
        );

    \I__5232\ : InMux
    port map (
            O => \N__26490\,
            I => \N__26470\
        );

    \I__5231\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26470\
        );

    \I__5230\ : InMux
    port map (
            O => \N__26488\,
            I => \N__26470\
        );

    \I__5229\ : InMux
    port map (
            O => \N__26487\,
            I => \N__26465\
        );

    \I__5228\ : InMux
    port map (
            O => \N__26486\,
            I => \N__26465\
        );

    \I__5227\ : InMux
    port map (
            O => \N__26485\,
            I => \N__26455\
        );

    \I__5226\ : InMux
    port map (
            O => \N__26484\,
            I => \N__26455\
        );

    \I__5225\ : InMux
    port map (
            O => \N__26483\,
            I => \N__26455\
        );

    \I__5224\ : InMux
    port map (
            O => \N__26482\,
            I => \N__26446\
        );

    \I__5223\ : InMux
    port map (
            O => \N__26481\,
            I => \N__26446\
        );

    \I__5222\ : InMux
    port map (
            O => \N__26480\,
            I => \N__26446\
        );

    \I__5221\ : InMux
    port map (
            O => \N__26479\,
            I => \N__26446\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__26470\,
            I => \N__26441\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__26465\,
            I => \N__26441\
        );

    \I__5218\ : InMux
    port map (
            O => \N__26464\,
            I => \N__26433\
        );

    \I__5217\ : InMux
    port map (
            O => \N__26463\,
            I => \N__26433\
        );

    \I__5216\ : InMux
    port map (
            O => \N__26462\,
            I => \N__26433\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__26455\,
            I => \N__26428\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__26446\,
            I => \N__26428\
        );

    \I__5213\ : Span4Mux_h
    port map (
            O => \N__26441\,
            I => \N__26425\
        );

    \I__5212\ : InMux
    port map (
            O => \N__26440\,
            I => \N__26422\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__26433\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__5210\ : Odrv4
    port map (
            O => \N__26428\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__5209\ : Odrv4
    port map (
            O => \N__26425\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__26422\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__5207\ : InMux
    port map (
            O => \N__26413\,
            I => \N__26410\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__26410\,
            I => \b2v_inst11.count_0_1\
        );

    \I__5205\ : InMux
    port map (
            O => \N__26407\,
            I => \N__26404\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__26404\,
            I => \N__26400\
        );

    \I__5203\ : InMux
    port map (
            O => \N__26403\,
            I => \N__26397\
        );

    \I__5202\ : Span4Mux_h
    port map (
            O => \N__26400\,
            I => \N__26393\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__26397\,
            I => \N__26390\
        );

    \I__5200\ : InMux
    port map (
            O => \N__26396\,
            I => \N__26387\
        );

    \I__5199\ : Odrv4
    port map (
            O => \N__26393\,
            I => \b2v_inst11.countZ0Z_8\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__26390\,
            I => \b2v_inst11.countZ0Z_8\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__26387\,
            I => \b2v_inst11.countZ0Z_8\
        );

    \I__5196\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26374\
        );

    \I__5195\ : InMux
    port map (
            O => \N__26379\,
            I => \N__26374\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__26374\,
            I => \b2v_inst11.un1_count_cry_7_c_RNIOU0EZ0\
        );

    \I__5193\ : InMux
    port map (
            O => \N__26371\,
            I => \N__26368\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__26368\,
            I => \b2v_inst11.count_0_8\
        );

    \I__5191\ : CascadeMux
    port map (
            O => \N__26365\,
            I => \N__26361\
        );

    \I__5190\ : InMux
    port map (
            O => \N__26364\,
            I => \N__26358\
        );

    \I__5189\ : InMux
    port map (
            O => \N__26361\,
            I => \N__26355\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__26358\,
            I => \N__26351\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__26355\,
            I => \N__26348\
        );

    \I__5186\ : CascadeMux
    port map (
            O => \N__26354\,
            I => \N__26345\
        );

    \I__5185\ : Span4Mux_h
    port map (
            O => \N__26351\,
            I => \N__26342\
        );

    \I__5184\ : Span4Mux_s3_h
    port map (
            O => \N__26348\,
            I => \N__26339\
        );

    \I__5183\ : InMux
    port map (
            O => \N__26345\,
            I => \N__26336\
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__26342\,
            I => \b2v_inst11.countZ0Z_9\
        );

    \I__5181\ : Odrv4
    port map (
            O => \N__26339\,
            I => \b2v_inst11.countZ0Z_9\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__26336\,
            I => \b2v_inst11.countZ0Z_9\
        );

    \I__5179\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26323\
        );

    \I__5178\ : InMux
    port map (
            O => \N__26328\,
            I => \N__26323\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__26323\,
            I => \b2v_inst11.un1_count_cry_8_c_RNIP02EZ0\
        );

    \I__5176\ : InMux
    port map (
            O => \N__26320\,
            I => \N__26317\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__26317\,
            I => \b2v_inst11.count_0_9\
        );

    \I__5174\ : InMux
    port map (
            O => \N__26314\,
            I => \N__26311\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__26311\,
            I => \b2v_inst5.curr_state_3_0\
        );

    \I__5172\ : CascadeMux
    port map (
            O => \N__26308\,
            I => \N__26302\
        );

    \I__5171\ : InMux
    port map (
            O => \N__26307\,
            I => \N__26298\
        );

    \I__5170\ : InMux
    port map (
            O => \N__26306\,
            I => \N__26289\
        );

    \I__5169\ : InMux
    port map (
            O => \N__26305\,
            I => \N__26289\
        );

    \I__5168\ : InMux
    port map (
            O => \N__26302\,
            I => \N__26289\
        );

    \I__5167\ : InMux
    port map (
            O => \N__26301\,
            I => \N__26289\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__26298\,
            I => \b2v_inst5.curr_stateZ0Z_0\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__26289\,
            I => \b2v_inst5.curr_stateZ0Z_0\
        );

    \I__5164\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26279\
        );

    \I__5163\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26274\
        );

    \I__5162\ : InMux
    port map (
            O => \N__26282\,
            I => \N__26274\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__26279\,
            I => \G_2727\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__26274\,
            I => \G_2727\
        );

    \I__5159\ : CascadeMux
    port map (
            O => \N__26269\,
            I => \b2v_inst5.curr_stateZ0Z_0_cascade_\
        );

    \I__5158\ : InMux
    port map (
            O => \N__26266\,
            I => \N__26263\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__26263\,
            I => \b2v_inst5.m4_0\
        );

    \I__5156\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26257\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__26257\,
            I => \N__26254\
        );

    \I__5154\ : Span4Mux_h
    port map (
            O => \N__26254\,
            I => \N__26250\
        );

    \I__5153\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26247\
        );

    \I__5152\ : Span4Mux_v
    port map (
            O => \N__26250\,
            I => \N__26244\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__26247\,
            I => \N__26241\
        );

    \I__5150\ : Odrv4
    port map (
            O => \N__26244\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1\
        );

    \I__5149\ : Odrv12
    port map (
            O => \N__26241\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1\
        );

    \I__5148\ : InMux
    port map (
            O => \N__26236\,
            I => \N__26225\
        );

    \I__5147\ : InMux
    port map (
            O => \N__26235\,
            I => \N__26225\
        );

    \I__5146\ : InMux
    port map (
            O => \N__26234\,
            I => \N__26220\
        );

    \I__5145\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26216\
        );

    \I__5144\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26207\
        );

    \I__5143\ : CascadeMux
    port map (
            O => \N__26231\,
            I => \N__26204\
        );

    \I__5142\ : CascadeMux
    port map (
            O => \N__26230\,
            I => \N__26200\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__26225\,
            I => \N__26196\
        );

    \I__5140\ : CascadeMux
    port map (
            O => \N__26224\,
            I => \N__26193\
        );

    \I__5139\ : InMux
    port map (
            O => \N__26223\,
            I => \N__26190\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__26220\,
            I => \N__26184\
        );

    \I__5137\ : InMux
    port map (
            O => \N__26219\,
            I => \N__26181\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__26216\,
            I => \N__26175\
        );

    \I__5135\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26168\
        );

    \I__5134\ : InMux
    port map (
            O => \N__26214\,
            I => \N__26168\
        );

    \I__5133\ : InMux
    port map (
            O => \N__26213\,
            I => \N__26168\
        );

    \I__5132\ : InMux
    port map (
            O => \N__26212\,
            I => \N__26163\
        );

    \I__5131\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26163\
        );

    \I__5130\ : InMux
    port map (
            O => \N__26210\,
            I => \N__26160\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__26207\,
            I => \N__26157\
        );

    \I__5128\ : InMux
    port map (
            O => \N__26204\,
            I => \N__26148\
        );

    \I__5127\ : InMux
    port map (
            O => \N__26203\,
            I => \N__26148\
        );

    \I__5126\ : InMux
    port map (
            O => \N__26200\,
            I => \N__26148\
        );

    \I__5125\ : InMux
    port map (
            O => \N__26199\,
            I => \N__26148\
        );

    \I__5124\ : Span4Mux_v
    port map (
            O => \N__26196\,
            I => \N__26145\
        );

    \I__5123\ : InMux
    port map (
            O => \N__26193\,
            I => \N__26142\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__26190\,
            I => \N__26139\
        );

    \I__5121\ : InMux
    port map (
            O => \N__26189\,
            I => \N__26134\
        );

    \I__5120\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26134\
        );

    \I__5119\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26131\
        );

    \I__5118\ : Span4Mux_h
    port map (
            O => \N__26184\,
            I => \N__26126\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__26181\,
            I => \N__26126\
        );

    \I__5116\ : InMux
    port map (
            O => \N__26180\,
            I => \N__26119\
        );

    \I__5115\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26119\
        );

    \I__5114\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26119\
        );

    \I__5113\ : Span4Mux_h
    port map (
            O => \N__26175\,
            I => \N__26112\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__26168\,
            I => \N__26112\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__26163\,
            I => \N__26112\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__26160\,
            I => \N__26105\
        );

    \I__5109\ : Span4Mux_v
    port map (
            O => \N__26157\,
            I => \N__26105\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__26148\,
            I => \N__26105\
        );

    \I__5107\ : Odrv4
    port map (
            O => \N__26145\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__26142\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__5105\ : Odrv12
    port map (
            O => \N__26139\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__26134\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__26131\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__5102\ : Odrv4
    port map (
            O => \N__26126\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__26119\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__5100\ : Odrv4
    port map (
            O => \N__26112\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__5099\ : Odrv4
    port map (
            O => \N__26105\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__5098\ : InMux
    port map (
            O => \N__26086\,
            I => \N__26080\
        );

    \I__5097\ : InMux
    port map (
            O => \N__26085\,
            I => \N__26080\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__26080\,
            I => \b2v_inst11.un1_count_cry_2_c_RNIJKRDZ0\
        );

    \I__5095\ : InMux
    port map (
            O => \N__26077\,
            I => \N__26074\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__26074\,
            I => \b2v_inst11.count_0_3\
        );

    \I__5093\ : InMux
    port map (
            O => \N__26071\,
            I => \N__26067\
        );

    \I__5092\ : CascadeMux
    port map (
            O => \N__26070\,
            I => \N__26063\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__26067\,
            I => \N__26060\
        );

    \I__5090\ : InMux
    port map (
            O => \N__26066\,
            I => \N__26057\
        );

    \I__5089\ : InMux
    port map (
            O => \N__26063\,
            I => \N__26054\
        );

    \I__5088\ : Odrv4
    port map (
            O => \N__26060\,
            I => \b2v_inst11.countZ0Z_13\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__26057\,
            I => \b2v_inst11.countZ0Z_13\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__26054\,
            I => \b2v_inst11.countZ0Z_13\
        );

    \I__5085\ : CascadeMux
    port map (
            O => \N__26047\,
            I => \N__26044\
        );

    \I__5084\ : InMux
    port map (
            O => \N__26044\,
            I => \N__26038\
        );

    \I__5083\ : InMux
    port map (
            O => \N__26043\,
            I => \N__26038\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__26038\,
            I => \b2v_inst11.un1_count_cry_12_c_RNI48TZ0Z6\
        );

    \I__5081\ : InMux
    port map (
            O => \N__26035\,
            I => \N__26032\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__26032\,
            I => \b2v_inst11.count_0_13\
        );

    \I__5079\ : InMux
    port map (
            O => \N__26029\,
            I => \N__26026\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__26026\,
            I => \N__26022\
        );

    \I__5077\ : CascadeMux
    port map (
            O => \N__26025\,
            I => \N__26018\
        );

    \I__5076\ : Span4Mux_v
    port map (
            O => \N__26022\,
            I => \N__26015\
        );

    \I__5075\ : InMux
    port map (
            O => \N__26021\,
            I => \N__26012\
        );

    \I__5074\ : InMux
    port map (
            O => \N__26018\,
            I => \N__26009\
        );

    \I__5073\ : Odrv4
    port map (
            O => \N__26015\,
            I => \b2v_inst11.countZ0Z_4\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__26012\,
            I => \b2v_inst11.countZ0Z_4\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__26009\,
            I => \b2v_inst11.countZ0Z_4\
        );

    \I__5070\ : InMux
    port map (
            O => \N__26002\,
            I => \N__25996\
        );

    \I__5069\ : InMux
    port map (
            O => \N__26001\,
            I => \N__25996\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__25996\,
            I => \b2v_inst11.un1_count_cry_3_c_RNIKMSDZ0\
        );

    \I__5067\ : InMux
    port map (
            O => \N__25993\,
            I => \N__25990\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__25990\,
            I => \b2v_inst11.count_0_4\
        );

    \I__5065\ : InMux
    port map (
            O => \N__25987\,
            I => \N__25984\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__25984\,
            I => \N__25980\
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__25983\,
            I => \N__25976\
        );

    \I__5062\ : Span4Mux_v
    port map (
            O => \N__25980\,
            I => \N__25973\
        );

    \I__5061\ : InMux
    port map (
            O => \N__25979\,
            I => \N__25970\
        );

    \I__5060\ : InMux
    port map (
            O => \N__25976\,
            I => \N__25967\
        );

    \I__5059\ : Odrv4
    port map (
            O => \N__25973\,
            I => \b2v_inst11.countZ0Z_5\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__25970\,
            I => \b2v_inst11.countZ0Z_5\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__25967\,
            I => \b2v_inst11.countZ0Z_5\
        );

    \I__5056\ : InMux
    port map (
            O => \N__25960\,
            I => \N__25954\
        );

    \I__5055\ : InMux
    port map (
            O => \N__25959\,
            I => \N__25954\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__25954\,
            I => \b2v_inst11.un1_count_cry_4_c_RNILOTDZ0\
        );

    \I__5053\ : InMux
    port map (
            O => \N__25951\,
            I => \N__25948\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__25948\,
            I => \b2v_inst11.count_0_5\
        );

    \I__5051\ : InMux
    port map (
            O => \N__25945\,
            I => \N__25942\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__25942\,
            I => \N__25939\
        );

    \I__5049\ : Span4Mux_v
    port map (
            O => \N__25939\,
            I => \N__25936\
        );

    \I__5048\ : Odrv4
    port map (
            O => \N__25936\,
            I => \b2v_inst11.count_0_0\
        );

    \I__5047\ : InMux
    port map (
            O => \N__25933\,
            I => \N__25930\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__25930\,
            I => \N__25927\
        );

    \I__5045\ : Odrv4
    port map (
            O => \N__25927\,
            I => \b2v_inst11.count_RNI_2_0\
        );

    \I__5044\ : CascadeMux
    port map (
            O => \N__25924\,
            I => \b2v_inst11.countZ0Z_0_cascade_\
        );

    \I__5043\ : CascadeMux
    port map (
            O => \N__25921\,
            I => \N__25916\
        );

    \I__5042\ : InMux
    port map (
            O => \N__25920\,
            I => \N__25913\
        );

    \I__5041\ : InMux
    port map (
            O => \N__25919\,
            I => \N__25910\
        );

    \I__5040\ : InMux
    port map (
            O => \N__25916\,
            I => \N__25907\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__25913\,
            I => \N__25904\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__25910\,
            I => \N__25899\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__25907\,
            I => \N__25899\
        );

    \I__5036\ : Odrv4
    port map (
            O => \N__25904\,
            I => \b2v_inst11.countZ0Z_2\
        );

    \I__5035\ : Odrv4
    port map (
            O => \N__25899\,
            I => \b2v_inst11.countZ0Z_2\
        );

    \I__5034\ : InMux
    port map (
            O => \N__25894\,
            I => \N__25890\
        );

    \I__5033\ : CascadeMux
    port map (
            O => \N__25893\,
            I => \N__25886\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__25890\,
            I => \N__25883\
        );

    \I__5031\ : InMux
    port map (
            O => \N__25889\,
            I => \N__25880\
        );

    \I__5030\ : InMux
    port map (
            O => \N__25886\,
            I => \N__25877\
        );

    \I__5029\ : Odrv4
    port map (
            O => \N__25883\,
            I => \b2v_inst11.countZ0Z_7\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__25880\,
            I => \b2v_inst11.countZ0Z_7\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__25877\,
            I => \b2v_inst11.countZ0Z_7\
        );

    \I__5026\ : InMux
    port map (
            O => \N__25870\,
            I => \N__25867\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__25867\,
            I => \N__25863\
        );

    \I__5024\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25859\
        );

    \I__5023\ : Span12Mux_s11_v
    port map (
            O => \N__25863\,
            I => \N__25856\
        );

    \I__5022\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25853\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__25859\,
            I => \b2v_inst11.countZ0Z_15\
        );

    \I__5020\ : Odrv12
    port map (
            O => \N__25856\,
            I => \b2v_inst11.countZ0Z_15\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__25853\,
            I => \b2v_inst11.countZ0Z_15\
        );

    \I__5018\ : InMux
    port map (
            O => \N__25846\,
            I => \N__25843\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__25843\,
            I => \N__25839\
        );

    \I__5016\ : InMux
    port map (
            O => \N__25842\,
            I => \N__25836\
        );

    \I__5015\ : Span4Mux_v
    port map (
            O => \N__25839\,
            I => \N__25832\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__25836\,
            I => \N__25829\
        );

    \I__5013\ : InMux
    port map (
            O => \N__25835\,
            I => \N__25826\
        );

    \I__5012\ : Odrv4
    port map (
            O => \N__25832\,
            I => \b2v_inst11.countZ0Z_11\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__25829\,
            I => \b2v_inst11.countZ0Z_11\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__25826\,
            I => \b2v_inst11.countZ0Z_11\
        );

    \I__5009\ : InMux
    port map (
            O => \N__25819\,
            I => \N__25816\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__25816\,
            I => \N__25811\
        );

    \I__5007\ : InMux
    port map (
            O => \N__25815\,
            I => \N__25808\
        );

    \I__5006\ : CascadeMux
    port map (
            O => \N__25814\,
            I => \N__25805\
        );

    \I__5005\ : Span4Mux_v
    port map (
            O => \N__25811\,
            I => \N__25802\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__25808\,
            I => \N__25799\
        );

    \I__5003\ : InMux
    port map (
            O => \N__25805\,
            I => \N__25796\
        );

    \I__5002\ : Odrv4
    port map (
            O => \N__25802\,
            I => \b2v_inst11.countZ0Z_10\
        );

    \I__5001\ : Odrv4
    port map (
            O => \N__25799\,
            I => \b2v_inst11.countZ0Z_10\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__25796\,
            I => \b2v_inst11.countZ0Z_10\
        );

    \I__4999\ : InMux
    port map (
            O => \N__25789\,
            I => \N__25784\
        );

    \I__4998\ : CascadeMux
    port map (
            O => \N__25788\,
            I => \N__25781\
        );

    \I__4997\ : InMux
    port map (
            O => \N__25787\,
            I => \N__25778\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__25784\,
            I => \N__25775\
        );

    \I__4995\ : InMux
    port map (
            O => \N__25781\,
            I => \N__25772\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__25778\,
            I => \b2v_inst11.countZ0Z_12\
        );

    \I__4993\ : Odrv4
    port map (
            O => \N__25775\,
            I => \b2v_inst11.countZ0Z_12\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__25772\,
            I => \b2v_inst11.countZ0Z_12\
        );

    \I__4991\ : InMux
    port map (
            O => \N__25765\,
            I => \N__25762\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__25762\,
            I => \b2v_inst11.un79_clk_100khzlt6\
        );

    \I__4989\ : CascadeMux
    port map (
            O => \N__25759\,
            I => \N__25754\
        );

    \I__4988\ : InMux
    port map (
            O => \N__25758\,
            I => \N__25751\
        );

    \I__4987\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25748\
        );

    \I__4986\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25745\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__25751\,
            I => \b2v_inst11.countZ0Z_6\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__25748\,
            I => \b2v_inst11.countZ0Z_6\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__25745\,
            I => \b2v_inst11.countZ0Z_6\
        );

    \I__4982\ : CascadeMux
    port map (
            O => \N__25738\,
            I => \b2v_inst11.un79_clk_100khzlto15_5_cascade_\
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__25735\,
            I => \N__25732\
        );

    \I__4980\ : InMux
    port map (
            O => \N__25732\,
            I => \N__25727\
        );

    \I__4979\ : InMux
    port map (
            O => \N__25731\,
            I => \N__25724\
        );

    \I__4978\ : InMux
    port map (
            O => \N__25730\,
            I => \N__25721\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__25727\,
            I => \N__25718\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__25724\,
            I => \b2v_inst11.countZ0Z_14\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__25721\,
            I => \b2v_inst11.countZ0Z_14\
        );

    \I__4974\ : Odrv4
    port map (
            O => \N__25718\,
            I => \b2v_inst11.countZ0Z_14\
        );

    \I__4973\ : CascadeMux
    port map (
            O => \N__25711\,
            I => \b2v_inst11.un79_clk_100khzlto15_7_cascade_\
        );

    \I__4972\ : InMux
    port map (
            O => \N__25708\,
            I => \N__25705\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__25705\,
            I => \b2v_inst11.un79_clk_100khzlto15_4\
        );

    \I__4970\ : CascadeMux
    port map (
            O => \N__25702\,
            I => \N__25697\
        );

    \I__4969\ : InMux
    port map (
            O => \N__25701\,
            I => \N__25693\
        );

    \I__4968\ : InMux
    port map (
            O => \N__25700\,
            I => \N__25686\
        );

    \I__4967\ : InMux
    port map (
            O => \N__25697\,
            I => \N__25686\
        );

    \I__4966\ : InMux
    port map (
            O => \N__25696\,
            I => \N__25686\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__25693\,
            I => \N__25683\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__25686\,
            I => \N__25680\
        );

    \I__4963\ : Span4Mux_v
    port map (
            O => \N__25683\,
            I => \N__25676\
        );

    \I__4962\ : Span4Mux_h
    port map (
            O => \N__25680\,
            I => \N__25673\
        );

    \I__4961\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25670\
        );

    \I__4960\ : Odrv4
    port map (
            O => \N__25676\,
            I => \b2v_inst11.count_RNIZ0Z_13\
        );

    \I__4959\ : Odrv4
    port map (
            O => \N__25673\,
            I => \b2v_inst11.count_RNIZ0Z_13\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__25670\,
            I => \b2v_inst11.count_RNIZ0Z_13\
        );

    \I__4957\ : InMux
    port map (
            O => \N__25663\,
            I => \N__25657\
        );

    \I__4956\ : InMux
    port map (
            O => \N__25662\,
            I => \N__25657\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__25657\,
            I => \N__25649\
        );

    \I__4954\ : InMux
    port map (
            O => \N__25656\,
            I => \N__25646\
        );

    \I__4953\ : InMux
    port map (
            O => \N__25655\,
            I => \N__25637\
        );

    \I__4952\ : InMux
    port map (
            O => \N__25654\,
            I => \N__25637\
        );

    \I__4951\ : InMux
    port map (
            O => \N__25653\,
            I => \N__25637\
        );

    \I__4950\ : InMux
    port map (
            O => \N__25652\,
            I => \N__25637\
        );

    \I__4949\ : Span4Mux_v
    port map (
            O => \N__25649\,
            I => \N__25634\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__25646\,
            I => \b2v_inst11.curr_stateZ0Z_0\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__25637\,
            I => \b2v_inst11.curr_stateZ0Z_0\
        );

    \I__4946\ : Odrv4
    port map (
            O => \N__25634\,
            I => \b2v_inst11.curr_stateZ0Z_0\
        );

    \I__4945\ : CascadeMux
    port map (
            O => \N__25627\,
            I => \b2v_inst11.count_RNIZ0Z_13_cascade_\
        );

    \I__4944\ : InMux
    port map (
            O => \N__25624\,
            I => \N__25621\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__25621\,
            I => \N__25617\
        );

    \I__4942\ : CascadeMux
    port map (
            O => \N__25620\,
            I => \N__25613\
        );

    \I__4941\ : Span4Mux_v
    port map (
            O => \N__25617\,
            I => \N__25610\
        );

    \I__4940\ : InMux
    port map (
            O => \N__25616\,
            I => \N__25607\
        );

    \I__4939\ : InMux
    port map (
            O => \N__25613\,
            I => \N__25604\
        );

    \I__4938\ : Odrv4
    port map (
            O => \N__25610\,
            I => \b2v_inst11.countZ0Z_3\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__25607\,
            I => \b2v_inst11.countZ0Z_3\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__25604\,
            I => \b2v_inst11.countZ0Z_3\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__25597\,
            I => \N__25591\
        );

    \I__4934\ : CascadeMux
    port map (
            O => \N__25596\,
            I => \N__25586\
        );

    \I__4933\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25583\
        );

    \I__4932\ : InMux
    port map (
            O => \N__25594\,
            I => \N__25578\
        );

    \I__4931\ : InMux
    port map (
            O => \N__25591\,
            I => \N__25578\
        );

    \I__4930\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25575\
        );

    \I__4929\ : InMux
    port map (
            O => \N__25589\,
            I => \N__25572\
        );

    \I__4928\ : InMux
    port map (
            O => \N__25586\,
            I => \N__25567\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__25583\,
            I => \N__25562\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__25578\,
            I => \N__25562\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__25575\,
            I => \N__25559\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__25572\,
            I => \N__25556\
        );

    \I__4923\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25553\
        );

    \I__4922\ : CascadeMux
    port map (
            O => \N__25570\,
            I => \N__25545\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__25567\,
            I => \N__25540\
        );

    \I__4920\ : Span4Mux_h
    port map (
            O => \N__25562\,
            I => \N__25540\
        );

    \I__4919\ : Span12Mux_s5_h
    port map (
            O => \N__25559\,
            I => \N__25537\
        );

    \I__4918\ : Span4Mux_v
    port map (
            O => \N__25556\,
            I => \N__25534\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__25553\,
            I => \N__25531\
        );

    \I__4916\ : InMux
    port map (
            O => \N__25552\,
            I => \N__25528\
        );

    \I__4915\ : InMux
    port map (
            O => \N__25551\,
            I => \N__25525\
        );

    \I__4914\ : InMux
    port map (
            O => \N__25550\,
            I => \N__25520\
        );

    \I__4913\ : InMux
    port map (
            O => \N__25549\,
            I => \N__25520\
        );

    \I__4912\ : InMux
    port map (
            O => \N__25548\,
            I => \N__25517\
        );

    \I__4911\ : InMux
    port map (
            O => \N__25545\,
            I => \N__25514\
        );

    \I__4910\ : Span4Mux_v
    port map (
            O => \N__25540\,
            I => \N__25511\
        );

    \I__4909\ : Odrv12
    port map (
            O => \N__25537\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__4908\ : Odrv4
    port map (
            O => \N__25534\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__4907\ : Odrv4
    port map (
            O => \N__25531\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__25528\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__25525\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__25520\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__25517\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__25514\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__4901\ : Odrv4
    port map (
            O => \N__25511\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__4900\ : InMux
    port map (
            O => \N__25492\,
            I => \N__25489\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__25489\,
            I => \b2v_inst11.mult1_un159_sum_cry_2_s\
        );

    \I__4898\ : CascadeMux
    port map (
            O => \N__25486\,
            I => \N__25483\
        );

    \I__4897\ : InMux
    port map (
            O => \N__25483\,
            I => \N__25480\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__25480\,
            I => \b2v_inst11.mult1_un159_sum_cry_3_s\
        );

    \I__4895\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25474\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__25474\,
            I => \b2v_inst11.mult1_un159_sum_cry_4_s\
        );

    \I__4893\ : CascadeMux
    port map (
            O => \N__25471\,
            I => \N__25468\
        );

    \I__4892\ : InMux
    port map (
            O => \N__25468\,
            I => \N__25457\
        );

    \I__4891\ : InMux
    port map (
            O => \N__25467\,
            I => \N__25457\
        );

    \I__4890\ : InMux
    port map (
            O => \N__25466\,
            I => \N__25457\
        );

    \I__4889\ : InMux
    port map (
            O => \N__25465\,
            I => \N__25454\
        );

    \I__4888\ : InMux
    port map (
            O => \N__25464\,
            I => \N__25451\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__25457\,
            I => \b2v_inst11.mult1_un159_sum_s_7\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__25454\,
            I => \b2v_inst11.mult1_un159_sum_s_7\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__25451\,
            I => \b2v_inst11.mult1_un159_sum_s_7\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__25444\,
            I => \N__25440\
        );

    \I__4883\ : InMux
    port map (
            O => \N__25443\,
            I => \N__25432\
        );

    \I__4882\ : InMux
    port map (
            O => \N__25440\,
            I => \N__25432\
        );

    \I__4881\ : InMux
    port map (
            O => \N__25439\,
            I => \N__25432\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__25432\,
            I => \G_2890\
        );

    \I__4879\ : CascadeMux
    port map (
            O => \N__25429\,
            I => \N__25426\
        );

    \I__4878\ : InMux
    port map (
            O => \N__25426\,
            I => \N__25423\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__25423\,
            I => \N__25420\
        );

    \I__4876\ : Odrv4
    port map (
            O => \N__25420\,
            I => \b2v_inst11.mult1_un159_sum_cry_5_s\
        );

    \I__4875\ : InMux
    port map (
            O => \N__25417\,
            I => \N__25414\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__25414\,
            I => \b2v_inst11.mult1_un166_sum_axb_6\
        );

    \I__4873\ : InMux
    port map (
            O => \N__25411\,
            I => \b2v_inst11.mult1_un166_sum_cry_5\
        );

    \I__4872\ : InMux
    port map (
            O => \N__25408\,
            I => \N__25405\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__25405\,
            I => \N__25402\
        );

    \I__4870\ : Span4Mux_v
    port map (
            O => \N__25402\,
            I => \N__25399\
        );

    \I__4869\ : Odrv4
    port map (
            O => \N__25399\,
            I => \b2v_inst11.un85_clk_100khz_0\
        );

    \I__4868\ : InMux
    port map (
            O => \N__25396\,
            I => \N__25393\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__25393\,
            I => \N__25386\
        );

    \I__4866\ : CascadeMux
    port map (
            O => \N__25392\,
            I => \N__25380\
        );

    \I__4865\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25376\
        );

    \I__4864\ : InMux
    port map (
            O => \N__25390\,
            I => \N__25371\
        );

    \I__4863\ : InMux
    port map (
            O => \N__25389\,
            I => \N__25371\
        );

    \I__4862\ : Span4Mux_v
    port map (
            O => \N__25386\,
            I => \N__25368\
        );

    \I__4861\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25365\
        );

    \I__4860\ : InMux
    port map (
            O => \N__25384\,
            I => \N__25361\
        );

    \I__4859\ : InMux
    port map (
            O => \N__25383\,
            I => \N__25355\
        );

    \I__4858\ : InMux
    port map (
            O => \N__25380\,
            I => \N__25355\
        );

    \I__4857\ : InMux
    port map (
            O => \N__25379\,
            I => \N__25352\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__25376\,
            I => \N__25347\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__25371\,
            I => \N__25347\
        );

    \I__4854\ : Span4Mux_h
    port map (
            O => \N__25368\,
            I => \N__25341\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__25365\,
            I => \N__25341\
        );

    \I__4852\ : InMux
    port map (
            O => \N__25364\,
            I => \N__25338\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__25361\,
            I => \N__25334\
        );

    \I__4850\ : CascadeMux
    port map (
            O => \N__25360\,
            I => \N__25330\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__25355\,
            I => \N__25327\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__25352\,
            I => \N__25322\
        );

    \I__4847\ : Span4Mux_v
    port map (
            O => \N__25347\,
            I => \N__25322\
        );

    \I__4846\ : InMux
    port map (
            O => \N__25346\,
            I => \N__25319\
        );

    \I__4845\ : Span4Mux_v
    port map (
            O => \N__25341\,
            I => \N__25315\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__25338\,
            I => \N__25312\
        );

    \I__4843\ : CascadeMux
    port map (
            O => \N__25337\,
            I => \N__25309\
        );

    \I__4842\ : Span4Mux_v
    port map (
            O => \N__25334\,
            I => \N__25305\
        );

    \I__4841\ : InMux
    port map (
            O => \N__25333\,
            I => \N__25300\
        );

    \I__4840\ : InMux
    port map (
            O => \N__25330\,
            I => \N__25300\
        );

    \I__4839\ : Span4Mux_h
    port map (
            O => \N__25327\,
            I => \N__25293\
        );

    \I__4838\ : Span4Mux_v
    port map (
            O => \N__25322\,
            I => \N__25293\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__25319\,
            I => \N__25293\
        );

    \I__4836\ : InMux
    port map (
            O => \N__25318\,
            I => \N__25290\
        );

    \I__4835\ : Span4Mux_v
    port map (
            O => \N__25315\,
            I => \N__25285\
        );

    \I__4834\ : Span4Mux_s3_v
    port map (
            O => \N__25312\,
            I => \N__25285\
        );

    \I__4833\ : InMux
    port map (
            O => \N__25309\,
            I => \N__25282\
        );

    \I__4832\ : InMux
    port map (
            O => \N__25308\,
            I => \N__25279\
        );

    \I__4831\ : Span4Mux_v
    port map (
            O => \N__25305\,
            I => \N__25274\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__25300\,
            I => \N__25274\
        );

    \I__4829\ : Span4Mux_s3_v
    port map (
            O => \N__25293\,
            I => \N__25271\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__25290\,
            I => \N__25268\
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__25285\,
            I => \b2v_inst11.dutycycle\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__25282\,
            I => \b2v_inst11.dutycycle\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__25279\,
            I => \b2v_inst11.dutycycle\
        );

    \I__4824\ : Odrv4
    port map (
            O => \N__25274\,
            I => \b2v_inst11.dutycycle\
        );

    \I__4823\ : Odrv4
    port map (
            O => \N__25271\,
            I => \b2v_inst11.dutycycle\
        );

    \I__4822\ : Odrv4
    port map (
            O => \N__25268\,
            I => \b2v_inst11.dutycycle\
        );

    \I__4821\ : CascadeMux
    port map (
            O => \N__25255\,
            I => \N__25252\
        );

    \I__4820\ : InMux
    port map (
            O => \N__25252\,
            I => \N__25249\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__25249\,
            I => \b2v_inst11.mult1_un159_sum_i\
        );

    \I__4818\ : InMux
    port map (
            O => \N__25246\,
            I => \b2v_inst36.un2_count_1_cry_13\
        );

    \I__4817\ : InMux
    port map (
            O => \N__25243\,
            I => \b2v_inst36.un2_count_1_cry_14\
        );

    \I__4816\ : InMux
    port map (
            O => \N__25240\,
            I => \N__25237\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__25237\,
            I => \b2v_inst36.count_1_12\
        );

    \I__4814\ : CascadeMux
    port map (
            O => \N__25234\,
            I => \b2v_inst36.count_en_cascade_\
        );

    \I__4813\ : InMux
    port map (
            O => \N__25231\,
            I => \N__25225\
        );

    \I__4812\ : InMux
    port map (
            O => \N__25230\,
            I => \N__25225\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__25225\,
            I => \b2v_inst36.count_rst_2\
        );

    \I__4810\ : InMux
    port map (
            O => \N__25222\,
            I => \N__25218\
        );

    \I__4809\ : InMux
    port map (
            O => \N__25221\,
            I => \N__25215\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__25218\,
            I => \b2v_inst36.count_rst_0\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__25215\,
            I => \b2v_inst36.count_rst_0\
        );

    \I__4806\ : InMux
    port map (
            O => \N__25210\,
            I => \N__25207\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__25207\,
            I => \N__25204\
        );

    \I__4804\ : Odrv4
    port map (
            O => \N__25204\,
            I => \b2v_inst36.count_1_14\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__25201\,
            I => \N__25198\
        );

    \I__4802\ : InMux
    port map (
            O => \N__25198\,
            I => \N__25192\
        );

    \I__4801\ : InMux
    port map (
            O => \N__25197\,
            I => \N__25192\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__25192\,
            I => \b2v_inst36.count_rst\
        );

    \I__4799\ : InMux
    port map (
            O => \N__25189\,
            I => \N__25186\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__25186\,
            I => \b2v_inst36.count_1_15\
        );

    \I__4797\ : InMux
    port map (
            O => \N__25183\,
            I => \b2v_inst36.un2_count_1_cry_5\
        );

    \I__4796\ : InMux
    port map (
            O => \N__25180\,
            I => \N__25176\
        );

    \I__4795\ : CascadeMux
    port map (
            O => \N__25179\,
            I => \N__25173\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__25176\,
            I => \N__25169\
        );

    \I__4793\ : InMux
    port map (
            O => \N__25173\,
            I => \N__25166\
        );

    \I__4792\ : InMux
    port map (
            O => \N__25172\,
            I => \N__25163\
        );

    \I__4791\ : Odrv4
    port map (
            O => \N__25169\,
            I => \b2v_inst36.countZ0Z_7\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__25166\,
            I => \b2v_inst36.countZ0Z_7\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__25163\,
            I => \b2v_inst36.countZ0Z_7\
        );

    \I__4788\ : InMux
    port map (
            O => \N__25156\,
            I => \N__25153\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__25153\,
            I => \N__25149\
        );

    \I__4786\ : InMux
    port map (
            O => \N__25152\,
            I => \N__25146\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__25149\,
            I => \b2v_inst36.un2_count_1_cry_6_THRU_CO\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__25146\,
            I => \b2v_inst36.un2_count_1_cry_6_THRU_CO\
        );

    \I__4783\ : InMux
    port map (
            O => \N__25141\,
            I => \b2v_inst36.un2_count_1_cry_6\
        );

    \I__4782\ : CascadeMux
    port map (
            O => \N__25138\,
            I => \N__25134\
        );

    \I__4781\ : InMux
    port map (
            O => \N__25137\,
            I => \N__25131\
        );

    \I__4780\ : InMux
    port map (
            O => \N__25134\,
            I => \N__25128\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__25131\,
            I => \b2v_inst36.un2_count_1_cry_7_THRU_CO\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__25128\,
            I => \b2v_inst36.un2_count_1_cry_7_THRU_CO\
        );

    \I__4777\ : InMux
    port map (
            O => \N__25123\,
            I => \b2v_inst36.un2_count_1_cry_7\
        );

    \I__4776\ : InMux
    port map (
            O => \N__25120\,
            I => \bfn_9_2_0_\
        );

    \I__4775\ : InMux
    port map (
            O => \N__25117\,
            I => \N__25111\
        );

    \I__4774\ : InMux
    port map (
            O => \N__25116\,
            I => \N__25111\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__25111\,
            I => \b2v_inst36.un2_count_1_cry_9_THRU_CO\
        );

    \I__4772\ : InMux
    port map (
            O => \N__25108\,
            I => \b2v_inst36.un2_count_1_cry_9\
        );

    \I__4771\ : InMux
    port map (
            O => \N__25105\,
            I => \b2v_inst36.un2_count_1_cry_10\
        );

    \I__4770\ : InMux
    port map (
            O => \N__25102\,
            I => \b2v_inst36.un2_count_1_cry_11\
        );

    \I__4769\ : InMux
    port map (
            O => \N__25099\,
            I => \b2v_inst36.un2_count_1_cry_12\
        );

    \I__4768\ : IoInMux
    port map (
            O => \N__25096\,
            I => \N__25093\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__25093\,
            I => \N__25090\
        );

    \I__4766\ : IoSpan4Mux
    port map (
            O => \N__25090\,
            I => \N__25087\
        );

    \I__4765\ : Span4Mux_s3_h
    port map (
            O => \N__25087\,
            I => \N__25082\
        );

    \I__4764\ : InMux
    port map (
            O => \N__25086\,
            I => \N__25079\
        );

    \I__4763\ : CascadeMux
    port map (
            O => \N__25085\,
            I => \N__25074\
        );

    \I__4762\ : Span4Mux_v
    port map (
            O => \N__25082\,
            I => \N__25068\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__25079\,
            I => \N__25068\
        );

    \I__4760\ : InMux
    port map (
            O => \N__25078\,
            I => \N__25056\
        );

    \I__4759\ : InMux
    port map (
            O => \N__25077\,
            I => \N__25056\
        );

    \I__4758\ : InMux
    port map (
            O => \N__25074\,
            I => \N__25056\
        );

    \I__4757\ : InMux
    port map (
            O => \N__25073\,
            I => \N__25056\
        );

    \I__4756\ : Span4Mux_v
    port map (
            O => \N__25068\,
            I => \N__25052\
        );

    \I__4755\ : InMux
    port map (
            O => \N__25067\,
            I => \N__25047\
        );

    \I__4754\ : InMux
    port map (
            O => \N__25066\,
            I => \N__25047\
        );

    \I__4753\ : InMux
    port map (
            O => \N__25065\,
            I => \N__25044\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__25056\,
            I => \N__25041\
        );

    \I__4751\ : InMux
    port map (
            O => \N__25055\,
            I => \N__25038\
        );

    \I__4750\ : Span4Mux_s0_v
    port map (
            O => \N__25052\,
            I => \N__25033\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__25047\,
            I => \N__25033\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__25044\,
            I => \N__25030\
        );

    \I__4747\ : Span4Mux_h
    port map (
            O => \N__25041\,
            I => \N__25027\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__25038\,
            I => \N__25022\
        );

    \I__4745\ : Span4Mux_h
    port map (
            O => \N__25033\,
            I => \N__25022\
        );

    \I__4744\ : Span4Mux_h
    port map (
            O => \N__25030\,
            I => \N__25019\
        );

    \I__4743\ : Span4Mux_v
    port map (
            O => \N__25027\,
            I => \N__25016\
        );

    \I__4742\ : Span4Mux_v
    port map (
            O => \N__25022\,
            I => \N__25013\
        );

    \I__4741\ : Odrv4
    port map (
            O => \N__25019\,
            I => \SYNTHESIZED_WIRE_49_i_0_o3_0\
        );

    \I__4740\ : Odrv4
    port map (
            O => \N__25016\,
            I => \SYNTHESIZED_WIRE_49_i_0_o3_0\
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__25013\,
            I => \SYNTHESIZED_WIRE_49_i_0_o3_0\
        );

    \I__4738\ : InMux
    port map (
            O => \N__25006\,
            I => \N__25003\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__25003\,
            I => \N__25000\
        );

    \I__4736\ : Span4Mux_v
    port map (
            O => \N__25000\,
            I => \N__24997\
        );

    \I__4735\ : Odrv4
    port map (
            O => \N__24997\,
            I => \VPP_OK_c\
        );

    \I__4734\ : IoInMux
    port map (
            O => \N__24994\,
            I => \N__24991\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__24991\,
            I => \N__24988\
        );

    \I__4732\ : IoSpan4Mux
    port map (
            O => \N__24988\,
            I => \N__24985\
        );

    \I__4731\ : Odrv4
    port map (
            O => \N__24985\,
            I => \VDDQ_EN_c\
        );

    \I__4730\ : InMux
    port map (
            O => \N__24982\,
            I => \N__24979\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__24979\,
            I => \VCCIO_OK_c\
        );

    \I__4728\ : InMux
    port map (
            O => \N__24976\,
            I => \N__24973\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__24973\,
            I => \V5S_OK_c\
        );

    \I__4726\ : CascadeMux
    port map (
            O => \N__24970\,
            I => \N__24967\
        );

    \I__4725\ : InMux
    port map (
            O => \N__24967\,
            I => \N__24964\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__24964\,
            I => \b2v_inst31.un8_outputZ0Z_0\
        );

    \I__4723\ : InMux
    port map (
            O => \N__24961\,
            I => \N__24958\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__24958\,
            I => \V33S_OK_c\
        );

    \I__4721\ : IoInMux
    port map (
            O => \N__24955\,
            I => \N__24951\
        );

    \I__4720\ : IoInMux
    port map (
            O => \N__24954\,
            I => \N__24948\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__24951\,
            I => \N__24943\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__24948\,
            I => \N__24943\
        );

    \I__4717\ : IoSpan4Mux
    port map (
            O => \N__24943\,
            I => \N__24940\
        );

    \I__4716\ : Span4Mux_s1_h
    port map (
            O => \N__24940\,
            I => \N__24937\
        );

    \I__4715\ : Span4Mux_h
    port map (
            O => \N__24937\,
            I => \N__24934\
        );

    \I__4714\ : Odrv4
    port map (
            O => \N__24934\,
            I => \VCCIN_EN_c\
        );

    \I__4713\ : InMux
    port map (
            O => \N__24931\,
            I => \b2v_inst36.un2_count_1_cry_1\
        );

    \I__4712\ : InMux
    port map (
            O => \N__24928\,
            I => \b2v_inst36.un2_count_1_cry_2\
        );

    \I__4711\ : InMux
    port map (
            O => \N__24925\,
            I => \b2v_inst36.un2_count_1_cry_3\
        );

    \I__4710\ : CascadeMux
    port map (
            O => \N__24922\,
            I => \N__24919\
        );

    \I__4709\ : InMux
    port map (
            O => \N__24919\,
            I => \N__24912\
        );

    \I__4708\ : InMux
    port map (
            O => \N__24918\,
            I => \N__24912\
        );

    \I__4707\ : InMux
    port map (
            O => \N__24917\,
            I => \N__24909\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__24912\,
            I => \b2v_inst36.countZ0Z_5\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__24909\,
            I => \b2v_inst36.countZ0Z_5\
        );

    \I__4704\ : InMux
    port map (
            O => \N__24904\,
            I => \N__24898\
        );

    \I__4703\ : InMux
    port map (
            O => \N__24903\,
            I => \N__24898\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__24898\,
            I => \b2v_inst36.un2_count_1_cry_4_THRU_CO\
        );

    \I__4701\ : InMux
    port map (
            O => \N__24895\,
            I => \b2v_inst36.un2_count_1_cry_4\
        );

    \I__4700\ : InMux
    port map (
            O => \N__24892\,
            I => \N__24889\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__24889\,
            I => \b2v_inst11.un1_clk_100khz_26_and_i_o2_1\
        );

    \I__4698\ : InMux
    port map (
            O => \N__24886\,
            I => \N__24883\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__24883\,
            I => \N__24880\
        );

    \I__4696\ : Odrv12
    port map (
            O => \N__24880\,
            I => \b2v_inst11.dutycycle_RNINJ641_0Z0Z_5\
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__24877\,
            I => \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_cascade_\
        );

    \I__4694\ : InMux
    port map (
            O => \N__24874\,
            I => \N__24871\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__24871\,
            I => \b2v_inst11.N_183\
        );

    \I__4692\ : InMux
    port map (
            O => \N__24868\,
            I => \N__24864\
        );

    \I__4691\ : InMux
    port map (
            O => \N__24867\,
            I => \N__24861\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__24864\,
            I => \N__24858\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__24861\,
            I => \N__24855\
        );

    \I__4688\ : Span12Mux_s4_h
    port map (
            O => \N__24858\,
            I => \N__24851\
        );

    \I__4687\ : Span4Mux_h
    port map (
            O => \N__24855\,
            I => \N__24848\
        );

    \I__4686\ : InMux
    port map (
            O => \N__24854\,
            I => \N__24845\
        );

    \I__4685\ : Odrv12
    port map (
            O => \N__24851\,
            I => \b2v_inst11.func_state_RNI_3Z0Z_1\
        );

    \I__4684\ : Odrv4
    port map (
            O => \N__24848\,
            I => \b2v_inst11.func_state_RNI_3Z0Z_1\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__24845\,
            I => \b2v_inst11.func_state_RNI_3Z0Z_1\
        );

    \I__4682\ : CascadeMux
    port map (
            O => \N__24838\,
            I => \b2v_inst11.N_183_cascade_\
        );

    \I__4681\ : InMux
    port map (
            O => \N__24835\,
            I => \N__24832\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__24832\,
            I => \N__24828\
        );

    \I__4679\ : InMux
    port map (
            O => \N__24831\,
            I => \N__24825\
        );

    \I__4678\ : Odrv4
    port map (
            O => \N__24828\,
            I => \b2v_inst11.N_114_f0_1\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__24825\,
            I => \b2v_inst11.N_114_f0_1\
        );

    \I__4676\ : InMux
    port map (
            O => \N__24820\,
            I => \N__24813\
        );

    \I__4675\ : InMux
    port map (
            O => \N__24819\,
            I => \N__24809\
        );

    \I__4674\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24802\
        );

    \I__4673\ : InMux
    port map (
            O => \N__24817\,
            I => \N__24802\
        );

    \I__4672\ : CascadeMux
    port map (
            O => \N__24816\,
            I => \N__24799\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__24813\,
            I => \N__24796\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__24812\,
            I => \N__24792\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24789\
        );

    \I__4668\ : CascadeMux
    port map (
            O => \N__24808\,
            I => \N__24786\
        );

    \I__4667\ : CascadeMux
    port map (
            O => \N__24807\,
            I => \N__24783\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__24802\,
            I => \N__24776\
        );

    \I__4665\ : InMux
    port map (
            O => \N__24799\,
            I => \N__24773\
        );

    \I__4664\ : Span4Mux_v
    port map (
            O => \N__24796\,
            I => \N__24770\
        );

    \I__4663\ : InMux
    port map (
            O => \N__24795\,
            I => \N__24767\
        );

    \I__4662\ : InMux
    port map (
            O => \N__24792\,
            I => \N__24764\
        );

    \I__4661\ : Span12Mux_s10_v
    port map (
            O => \N__24789\,
            I => \N__24761\
        );

    \I__4660\ : InMux
    port map (
            O => \N__24786\,
            I => \N__24754\
        );

    \I__4659\ : InMux
    port map (
            O => \N__24783\,
            I => \N__24754\
        );

    \I__4658\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24754\
        );

    \I__4657\ : InMux
    port map (
            O => \N__24781\,
            I => \N__24749\
        );

    \I__4656\ : InMux
    port map (
            O => \N__24780\,
            I => \N__24749\
        );

    \I__4655\ : InMux
    port map (
            O => \N__24779\,
            I => \N__24746\
        );

    \I__4654\ : Span4Mux_h
    port map (
            O => \N__24776\,
            I => \N__24741\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__24773\,
            I => \N__24741\
        );

    \I__4652\ : Odrv4
    port map (
            O => \N__24770\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__24767\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__24764\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__4649\ : Odrv12
    port map (
            O => \N__24761\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__24754\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__24749\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__24746\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__4645\ : Odrv4
    port map (
            O => \N__24741\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__4644\ : InMux
    port map (
            O => \N__24724\,
            I => \N__24717\
        );

    \I__4643\ : InMux
    port map (
            O => \N__24723\,
            I => \N__24717\
        );

    \I__4642\ : InMux
    port map (
            O => \N__24722\,
            I => \N__24713\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__24717\,
            I => \N__24710\
        );

    \I__4640\ : InMux
    port map (
            O => \N__24716\,
            I => \N__24707\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__24713\,
            I => \N__24702\
        );

    \I__4638\ : Span4Mux_s1_v
    port map (
            O => \N__24710\,
            I => \N__24702\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__24707\,
            I => \b2v_inst11.N_379\
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__24702\,
            I => \b2v_inst11.N_379\
        );

    \I__4635\ : CascadeMux
    port map (
            O => \N__24697\,
            I => \b2v_inst6.curr_state_RNI8OKQ2Z0Z_0_cascade_\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__24694\,
            I => \N__24691\
        );

    \I__4633\ : InMux
    port map (
            O => \N__24691\,
            I => \N__24684\
        );

    \I__4632\ : InMux
    port map (
            O => \N__24690\,
            I => \N__24684\
        );

    \I__4631\ : CascadeMux
    port map (
            O => \N__24689\,
            I => \N__24681\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__24684\,
            I => \N__24678\
        );

    \I__4629\ : InMux
    port map (
            O => \N__24681\,
            I => \N__24672\
        );

    \I__4628\ : Span4Mux_s1_v
    port map (
            O => \N__24678\,
            I => \N__24669\
        );

    \I__4627\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24664\
        );

    \I__4626\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24664\
        );

    \I__4625\ : InMux
    port map (
            O => \N__24675\,
            I => \N__24661\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__24672\,
            I => \b2v_inst11.un1_clk_100khz_52_and_i_a2Z0Z_1\
        );

    \I__4623\ : Odrv4
    port map (
            O => \N__24669\,
            I => \b2v_inst11.un1_clk_100khz_52_and_i_a2Z0Z_1\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__24664\,
            I => \b2v_inst11.un1_clk_100khz_52_and_i_a2Z0Z_1\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__24661\,
            I => \b2v_inst11.un1_clk_100khz_52_and_i_a2Z0Z_1\
        );

    \I__4620\ : InMux
    port map (
            O => \N__24652\,
            I => \N__24648\
        );

    \I__4619\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24645\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__24648\,
            I => \N__24642\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__24645\,
            I => \N__24639\
        );

    \I__4616\ : Span4Mux_h
    port map (
            O => \N__24642\,
            I => \N__24636\
        );

    \I__4615\ : Span4Mux_h
    port map (
            O => \N__24639\,
            I => \N__24633\
        );

    \I__4614\ : Odrv4
    port map (
            O => \N__24636\,
            I => \b2v_inst11.func_state_RNIDINH9Z0Z_0\
        );

    \I__4613\ : Odrv4
    port map (
            O => \N__24633\,
            I => \b2v_inst11.func_state_RNIDINH9Z0Z_0\
        );

    \I__4612\ : CascadeMux
    port map (
            O => \N__24628\,
            I => \N__24625\
        );

    \I__4611\ : InMux
    port map (
            O => \N__24625\,
            I => \N__24621\
        );

    \I__4610\ : InMux
    port map (
            O => \N__24624\,
            I => \N__24618\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__24621\,
            I => \N__24615\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__24618\,
            I => \b2v_inst11.func_stateZ0Z_1\
        );

    \I__4607\ : Odrv4
    port map (
            O => \N__24615\,
            I => \b2v_inst11.func_stateZ0Z_1\
        );

    \I__4606\ : InMux
    port map (
            O => \N__24610\,
            I => \N__24607\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__24607\,
            I => \b2v_inst6.curr_state_RNI8OKQ2Z0Z_0\
        );

    \I__4604\ : CascadeMux
    port map (
            O => \N__24604\,
            I => \N__24601\
        );

    \I__4603\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24595\
        );

    \I__4602\ : InMux
    port map (
            O => \N__24600\,
            I => \N__24595\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__24595\,
            I => \b2v_inst6.delayed_vccin_vccinaux_ok_0\
        );

    \I__4600\ : CascadeMux
    port map (
            O => \N__24592\,
            I => \b2v_inst11.func_state_cascade_\
        );

    \I__4599\ : CascadeMux
    port map (
            O => \N__24589\,
            I => \b2v_inst11.N_303_cascade_\
        );

    \I__4598\ : InMux
    port map (
            O => \N__24586\,
            I => \N__24583\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__24583\,
            I => \b2v_inst11.dutycycle_eena_1\
        );

    \I__4596\ : CascadeMux
    port map (
            O => \N__24580\,
            I => \N__24576\
        );

    \I__4595\ : InMux
    port map (
            O => \N__24579\,
            I => \N__24573\
        );

    \I__4594\ : InMux
    port map (
            O => \N__24576\,
            I => \N__24570\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__24573\,
            I => \N__24567\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__24570\,
            I => \N__24564\
        );

    \I__4591\ : Span4Mux_h
    port map (
            O => \N__24567\,
            I => \N__24559\
        );

    \I__4590\ : Span4Mux_h
    port map (
            O => \N__24564\,
            I => \N__24559\
        );

    \I__4589\ : Odrv4
    port map (
            O => \N__24559\,
            I => \b2v_inst11.N_70\
        );

    \I__4588\ : CascadeMux
    port map (
            O => \N__24556\,
            I => \b2v_inst11.dutycycle_eena_1_cascade_\
        );

    \I__4587\ : InMux
    port map (
            O => \N__24553\,
            I => \N__24547\
        );

    \I__4586\ : InMux
    port map (
            O => \N__24552\,
            I => \N__24547\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__24547\,
            I => \b2v_inst11.dutycycleZ1Z_2\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__24544\,
            I => \N__24541\
        );

    \I__4583\ : InMux
    port map (
            O => \N__24541\,
            I => \N__24538\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__24538\,
            I => \N__24534\
        );

    \I__4581\ : InMux
    port map (
            O => \N__24537\,
            I => \N__24531\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__24534\,
            I => \b2v_inst11.dutycycle_eena_0\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__24531\,
            I => \b2v_inst11.dutycycle_eena_0\
        );

    \I__4578\ : InMux
    port map (
            O => \N__24526\,
            I => \N__24522\
        );

    \I__4577\ : InMux
    port map (
            O => \N__24525\,
            I => \N__24519\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__24522\,
            I => \N__24516\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__24519\,
            I => \N__24513\
        );

    \I__4574\ : Span4Mux_v
    port map (
            O => \N__24516\,
            I => \N__24508\
        );

    \I__4573\ : Span4Mux_h
    port map (
            O => \N__24513\,
            I => \N__24505\
        );

    \I__4572\ : InMux
    port map (
            O => \N__24512\,
            I => \N__24500\
        );

    \I__4571\ : InMux
    port map (
            O => \N__24511\,
            I => \N__24500\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__24508\,
            I => \b2v_inst11.N_169\
        );

    \I__4569\ : Odrv4
    port map (
            O => \N__24505\,
            I => \b2v_inst11.N_169\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__24500\,
            I => \b2v_inst11.N_169\
        );

    \I__4567\ : InMux
    port map (
            O => \N__24493\,
            I => \N__24490\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__24490\,
            I => \b2v_inst11.N_375\
        );

    \I__4565\ : CascadeMux
    port map (
            O => \N__24487\,
            I => \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_sxZ0_cascade_\
        );

    \I__4564\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24478\
        );

    \I__4563\ : InMux
    port map (
            O => \N__24483\,
            I => \N__24473\
        );

    \I__4562\ : InMux
    port map (
            O => \N__24482\,
            I => \N__24473\
        );

    \I__4561\ : CascadeMux
    port map (
            O => \N__24481\,
            I => \N__24470\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__24478\,
            I => \N__24465\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__24473\,
            I => \N__24461\
        );

    \I__4558\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24456\
        );

    \I__4557\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24456\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__24468\,
            I => \N__24452\
        );

    \I__4555\ : Span4Mux_h
    port map (
            O => \N__24465\,
            I => \N__24449\
        );

    \I__4554\ : InMux
    port map (
            O => \N__24464\,
            I => \N__24446\
        );

    \I__4553\ : Sp12to4
    port map (
            O => \N__24461\,
            I => \N__24441\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__24456\,
            I => \N__24441\
        );

    \I__4551\ : InMux
    port map (
            O => \N__24455\,
            I => \N__24436\
        );

    \I__4550\ : InMux
    port map (
            O => \N__24452\,
            I => \N__24436\
        );

    \I__4549\ : Odrv4
    port map (
            O => \N__24449\,
            I => \SYNTHESIZED_WIRE_47keep_fast\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__24446\,
            I => \SYNTHESIZED_WIRE_47keep_fast\
        );

    \I__4547\ : Odrv12
    port map (
            O => \N__24441\,
            I => \SYNTHESIZED_WIRE_47keep_fast\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__24436\,
            I => \SYNTHESIZED_WIRE_47keep_fast\
        );

    \I__4545\ : InMux
    port map (
            O => \N__24427\,
            I => \N__24424\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__24424\,
            I => \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_1\
        );

    \I__4543\ : InMux
    port map (
            O => \N__24421\,
            I => \N__24418\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__24418\,
            I => \N__24415\
        );

    \I__4541\ : Odrv12
    port map (
            O => \N__24415\,
            I => \b2v_inst11.m15_e_3\
        );

    \I__4540\ : InMux
    port map (
            O => \N__24412\,
            I => \N__24409\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__24409\,
            I => \b2v_inst11.un1_dutycycle_inv_4_0\
        );

    \I__4538\ : InMux
    port map (
            O => \N__24406\,
            I => \N__24403\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__24403\,
            I => \N__24400\
        );

    \I__4536\ : Odrv4
    port map (
            O => \N__24400\,
            I => \b2v_inst11.g0_9_1\
        );

    \I__4535\ : CascadeMux
    port map (
            O => \N__24397\,
            I => \b2v_inst11.g1_0_1_cascade_\
        );

    \I__4534\ : InMux
    port map (
            O => \N__24394\,
            I => \N__24390\
        );

    \I__4533\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24387\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__24390\,
            I => \b2v_inst11.un1_dutycycle_164_0\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__24387\,
            I => \b2v_inst11.un1_dutycycle_164_0\
        );

    \I__4530\ : CascadeMux
    port map (
            O => \N__24382\,
            I => \N__24379\
        );

    \I__4529\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24375\
        );

    \I__4528\ : CascadeMux
    port map (
            O => \N__24378\,
            I => \N__24372\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__24375\,
            I => \N__24369\
        );

    \I__4526\ : InMux
    port map (
            O => \N__24372\,
            I => \N__24366\
        );

    \I__4525\ : Span4Mux_v
    port map (
            O => \N__24369\,
            I => \N__24361\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__24366\,
            I => \N__24358\
        );

    \I__4523\ : InMux
    port map (
            O => \N__24365\,
            I => \N__24353\
        );

    \I__4522\ : InMux
    port map (
            O => \N__24364\,
            I => \N__24353\
        );

    \I__4521\ : Span4Mux_h
    port map (
            O => \N__24361\,
            I => \N__24348\
        );

    \I__4520\ : Span4Mux_s2_v
    port map (
            O => \N__24358\,
            I => \N__24348\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__24353\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_5\
        );

    \I__4518\ : Odrv4
    port map (
            O => \N__24348\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_5\
        );

    \I__4517\ : CascadeMux
    port map (
            O => \N__24343\,
            I => \N__24340\
        );

    \I__4516\ : InMux
    port map (
            O => \N__24340\,
            I => \N__24337\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__24337\,
            I => \N__24334\
        );

    \I__4514\ : Span12Mux_s5_v
    port map (
            O => \N__24334\,
            I => \N__24331\
        );

    \I__4513\ : Odrv12
    port map (
            O => \N__24331\,
            I => \b2v_inst11.mult1_un152_sum_i\
        );

    \I__4512\ : InMux
    port map (
            O => \N__24328\,
            I => \N__24325\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__24325\,
            I => \N__24321\
        );

    \I__4510\ : InMux
    port map (
            O => \N__24324\,
            I => \N__24318\
        );

    \I__4509\ : Span4Mux_h
    port map (
            O => \N__24321\,
            I => \N__24308\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__24318\,
            I => \N__24308\
        );

    \I__4507\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24305\
        );

    \I__4506\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24302\
        );

    \I__4505\ : InMux
    port map (
            O => \N__24315\,
            I => \N__24298\
        );

    \I__4504\ : InMux
    port map (
            O => \N__24314\,
            I => \N__24295\
        );

    \I__4503\ : InMux
    port map (
            O => \N__24313\,
            I => \N__24292\
        );

    \I__4502\ : Span4Mux_h
    port map (
            O => \N__24308\,
            I => \N__24286\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__24305\,
            I => \N__24286\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__24302\,
            I => \N__24283\
        );

    \I__4499\ : InMux
    port map (
            O => \N__24301\,
            I => \N__24280\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__24298\,
            I => \N__24274\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__24295\,
            I => \N__24269\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__24292\,
            I => \N__24269\
        );

    \I__4495\ : InMux
    port map (
            O => \N__24291\,
            I => \N__24266\
        );

    \I__4494\ : Span4Mux_v
    port map (
            O => \N__24286\,
            I => \N__24259\
        );

    \I__4493\ : Span4Mux_h
    port map (
            O => \N__24283\,
            I => \N__24259\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__24280\,
            I => \N__24259\
        );

    \I__4491\ : InMux
    port map (
            O => \N__24279\,
            I => \N__24252\
        );

    \I__4490\ : InMux
    port map (
            O => \N__24278\,
            I => \N__24252\
        );

    \I__4489\ : InMux
    port map (
            O => \N__24277\,
            I => \N__24252\
        );

    \I__4488\ : Span4Mux_v
    port map (
            O => \N__24274\,
            I => \N__24247\
        );

    \I__4487\ : Span4Mux_h
    port map (
            O => \N__24269\,
            I => \N__24247\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__24266\,
            I => \b2v_inst11.N_3013_i\
        );

    \I__4485\ : Odrv4
    port map (
            O => \N__24259\,
            I => \b2v_inst11.N_3013_i\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__24252\,
            I => \b2v_inst11.N_3013_i\
        );

    \I__4483\ : Odrv4
    port map (
            O => \N__24247\,
            I => \b2v_inst11.N_3013_i\
        );

    \I__4482\ : SRMux
    port map (
            O => \N__24238\,
            I => \N__24233\
        );

    \I__4481\ : SRMux
    port map (
            O => \N__24237\,
            I => \N__24228\
        );

    \I__4480\ : SRMux
    port map (
            O => \N__24236\,
            I => \N__24224\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__24233\,
            I => \N__24221\
        );

    \I__4478\ : SRMux
    port map (
            O => \N__24232\,
            I => \N__24218\
        );

    \I__4477\ : SRMux
    port map (
            O => \N__24231\,
            I => \N__24215\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__24228\,
            I => \N__24211\
        );

    \I__4475\ : SRMux
    port map (
            O => \N__24227\,
            I => \N__24207\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__24224\,
            I => \N__24204\
        );

    \I__4473\ : Span4Mux_v
    port map (
            O => \N__24221\,
            I => \N__24197\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__24218\,
            I => \N__24197\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__24215\,
            I => \N__24197\
        );

    \I__4470\ : SRMux
    port map (
            O => \N__24214\,
            I => \N__24194\
        );

    \I__4469\ : Span4Mux_h
    port map (
            O => \N__24211\,
            I => \N__24191\
        );

    \I__4468\ : SRMux
    port map (
            O => \N__24210\,
            I => \N__24188\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__24207\,
            I => \N__24184\
        );

    \I__4466\ : Span4Mux_v
    port map (
            O => \N__24204\,
            I => \N__24179\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__24197\,
            I => \N__24179\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__24194\,
            I => \N__24176\
        );

    \I__4463\ : Sp12to4
    port map (
            O => \N__24191\,
            I => \N__24171\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__24188\,
            I => \N__24171\
        );

    \I__4461\ : SRMux
    port map (
            O => \N__24187\,
            I => \N__24168\
        );

    \I__4460\ : Span4Mux_h
    port map (
            O => \N__24184\,
            I => \N__24165\
        );

    \I__4459\ : Span4Mux_h
    port map (
            O => \N__24179\,
            I => \N__24157\
        );

    \I__4458\ : Span4Mux_v
    port map (
            O => \N__24176\,
            I => \N__24154\
        );

    \I__4457\ : Span12Mux_s6_v
    port map (
            O => \N__24171\,
            I => \N__24151\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__24168\,
            I => \N__24148\
        );

    \I__4455\ : Span4Mux_v
    port map (
            O => \N__24165\,
            I => \N__24145\
        );

    \I__4454\ : SRMux
    port map (
            O => \N__24164\,
            I => \N__24142\
        );

    \I__4453\ : SRMux
    port map (
            O => \N__24163\,
            I => \N__24139\
        );

    \I__4452\ : SRMux
    port map (
            O => \N__24162\,
            I => \N__24136\
        );

    \I__4451\ : SRMux
    port map (
            O => \N__24161\,
            I => \N__24133\
        );

    \I__4450\ : SRMux
    port map (
            O => \N__24160\,
            I => \N__24130\
        );

    \I__4449\ : Odrv4
    port map (
            O => \N__24157\,
            I => \b2v_inst11.N_221_iZ0\
        );

    \I__4448\ : Odrv4
    port map (
            O => \N__24154\,
            I => \b2v_inst11.N_221_iZ0\
        );

    \I__4447\ : Odrv12
    port map (
            O => \N__24151\,
            I => \b2v_inst11.N_221_iZ0\
        );

    \I__4446\ : Odrv12
    port map (
            O => \N__24148\,
            I => \b2v_inst11.N_221_iZ0\
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__24145\,
            I => \b2v_inst11.N_221_iZ0\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__24142\,
            I => \b2v_inst11.N_221_iZ0\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__24139\,
            I => \b2v_inst11.N_221_iZ0\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__24136\,
            I => \b2v_inst11.N_221_iZ0\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__24133\,
            I => \b2v_inst11.N_221_iZ0\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__24130\,
            I => \b2v_inst11.N_221_iZ0\
        );

    \I__4439\ : InMux
    port map (
            O => \N__24109\,
            I => \N__24106\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__24106\,
            I => \N__24103\
        );

    \I__4437\ : Span4Mux_v
    port map (
            O => \N__24103\,
            I => \N__24100\
        );

    \I__4436\ : Odrv4
    port map (
            O => \N__24100\,
            I => \b2v_inst11.g0_1_1\
        );

    \I__4435\ : CascadeMux
    port map (
            O => \N__24097\,
            I => \N__24093\
        );

    \I__4434\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24089\
        );

    \I__4433\ : InMux
    port map (
            O => \N__24093\,
            I => \N__24086\
        );

    \I__4432\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24083\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__24089\,
            I => \N__24079\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__24086\,
            I => \N__24076\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__24083\,
            I => \N__24073\
        );

    \I__4428\ : InMux
    port map (
            O => \N__24082\,
            I => \N__24070\
        );

    \I__4427\ : Span4Mux_s2_v
    port map (
            O => \N__24079\,
            I => \N__24067\
        );

    \I__4426\ : Span4Mux_s2_v
    port map (
            O => \N__24076\,
            I => \N__24062\
        );

    \I__4425\ : Span4Mux_s2_v
    port map (
            O => \N__24073\,
            I => \N__24062\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__24070\,
            I => \N__24059\
        );

    \I__4423\ : Span4Mux_v
    port map (
            O => \N__24067\,
            I => \N__24055\
        );

    \I__4422\ : Span4Mux_v
    port map (
            O => \N__24062\,
            I => \N__24052\
        );

    \I__4421\ : Span4Mux_s3_v
    port map (
            O => \N__24059\,
            I => \N__24049\
        );

    \I__4420\ : InMux
    port map (
            O => \N__24058\,
            I => \N__24046\
        );

    \I__4419\ : Odrv4
    port map (
            O => \N__24055\,
            I => \b2v_inst11.N_182\
        );

    \I__4418\ : Odrv4
    port map (
            O => \N__24052\,
            I => \b2v_inst11.N_182\
        );

    \I__4417\ : Odrv4
    port map (
            O => \N__24049\,
            I => \b2v_inst11.N_182\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__24046\,
            I => \b2v_inst11.N_182\
        );

    \I__4415\ : CascadeMux
    port map (
            O => \N__24037\,
            I => \N__24034\
        );

    \I__4414\ : InMux
    port map (
            O => \N__24034\,
            I => \N__24031\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__24031\,
            I => \b2v_inst11.func_state_RNIT4D71_0Z0Z_1\
        );

    \I__4412\ : InMux
    port map (
            O => \N__24028\,
            I => \N__24022\
        );

    \I__4411\ : InMux
    port map (
            O => \N__24027\,
            I => \N__24022\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__24022\,
            I => \b2v_inst11.dutycycle_0_5\
        );

    \I__4409\ : InMux
    port map (
            O => \N__24019\,
            I => \N__24013\
        );

    \I__4408\ : InMux
    port map (
            O => \N__24018\,
            I => \N__24013\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__24013\,
            I => \N__24010\
        );

    \I__4406\ : Span4Mux_h
    port map (
            O => \N__24010\,
            I => \N__24007\
        );

    \I__4405\ : Odrv4
    port map (
            O => \N__24007\,
            I => \b2v_inst11.g1_4_0\
        );

    \I__4404\ : CascadeMux
    port map (
            O => \N__24004\,
            I => \b2v_inst11.func_state_RNIT4D71_0Z0Z_1_cascade_\
        );

    \I__4403\ : CascadeMux
    port map (
            O => \N__24001\,
            I => \dutycycle_RNIIOE3D_0_5_cascade_\
        );

    \I__4402\ : CascadeMux
    port map (
            O => \N__23998\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_5_cascade_\
        );

    \I__4401\ : CascadeMux
    port map (
            O => \N__23995\,
            I => \b2v_inst11.un1_dutycycle_53_axb_3_1_cascade_\
        );

    \I__4400\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23989\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__23989\,
            I => \N__23986\
        );

    \I__4398\ : Span4Mux_h
    port map (
            O => \N__23986\,
            I => \N__23983\
        );

    \I__4397\ : Span4Mux_v
    port map (
            O => \N__23983\,
            I => \N__23980\
        );

    \I__4396\ : Odrv4
    port map (
            O => \N__23980\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_2\
        );

    \I__4395\ : InMux
    port map (
            O => \N__23977\,
            I => \N__23974\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__23974\,
            I => \b2v_inst11.un1_i3_mux_1\
        );

    \I__4393\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23968\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__23968\,
            I => \N__23965\
        );

    \I__4391\ : Span4Mux_h
    port map (
            O => \N__23965\,
            I => \N__23962\
        );

    \I__4390\ : Odrv4
    port map (
            O => \N__23962\,
            I => \b2v_inst11.g0_6_2\
        );

    \I__4389\ : CascadeMux
    port map (
            O => \N__23959\,
            I => \b2v_inst5.curr_stateZ0Z_1_cascade_\
        );

    \I__4388\ : CascadeMux
    port map (
            O => \N__23956\,
            I => \curr_state_RNI5VS71_0_1_cascade_\
        );

    \I__4387\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23950\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__23950\,
            I => \N__23946\
        );

    \I__4385\ : InMux
    port map (
            O => \N__23949\,
            I => \N__23943\
        );

    \I__4384\ : Span4Mux_s2_v
    port map (
            O => \N__23946\,
            I => \N__23938\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__23943\,
            I => \N__23938\
        );

    \I__4382\ : Span4Mux_v
    port map (
            O => \N__23938\,
            I => \N__23935\
        );

    \I__4381\ : Odrv4
    port map (
            O => \N__23935\,
            I => \b2v_inst11.mult1_un145_sum\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__23932\,
            I => \RSMRSTn_RNI8DFE_cascade_\
        );

    \I__4379\ : InMux
    port map (
            O => \N__23929\,
            I => \N__23926\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__23926\,
            I => \b2v_inst11.count_0_11\
        );

    \I__4377\ : InMux
    port map (
            O => \N__23923\,
            I => \N__23917\
        );

    \I__4376\ : InMux
    port map (
            O => \N__23922\,
            I => \N__23917\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__23917\,
            I => \N__23914\
        );

    \I__4374\ : Odrv4
    port map (
            O => \N__23914\,
            I => \b2v_inst11.un1_count_cry_1_c_RNIIIQDZ0\
        );

    \I__4373\ : InMux
    port map (
            O => \N__23911\,
            I => \N__23908\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__23908\,
            I => \b2v_inst11.count_0_2\
        );

    \I__4371\ : InMux
    port map (
            O => \N__23905\,
            I => \N__23901\
        );

    \I__4370\ : InMux
    port map (
            O => \N__23904\,
            I => \N__23898\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__23901\,
            I => \b2v_inst11.un1_count_cry_11_c_RNI36SZ0Z6\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__23898\,
            I => \b2v_inst11.un1_count_cry_11_c_RNI36SZ0Z6\
        );

    \I__4367\ : InMux
    port map (
            O => \N__23893\,
            I => \N__23890\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__23890\,
            I => \b2v_inst11.count_0_12\
        );

    \I__4365\ : CascadeMux
    port map (
            O => \N__23887\,
            I => \G_2727_cascade_\
        );

    \I__4364\ : InMux
    port map (
            O => \N__23884\,
            I => \N__23881\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__23881\,
            I => \b2v_inst5.curr_state_2_1\
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__23878\,
            I => \N_229_cascade_\
        );

    \I__4361\ : InMux
    port map (
            O => \N__23875\,
            I => \N__23863\
        );

    \I__4360\ : InMux
    port map (
            O => \N__23874\,
            I => \N__23863\
        );

    \I__4359\ : InMux
    port map (
            O => \N__23873\,
            I => \N__23863\
        );

    \I__4358\ : InMux
    port map (
            O => \N__23872\,
            I => \N__23863\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__23863\,
            I => \b2v_inst5.curr_stateZ0Z_1\
        );

    \I__4356\ : InMux
    port map (
            O => \N__23860\,
            I => \b2v_inst11.un1_count_cry_10\
        );

    \I__4355\ : InMux
    port map (
            O => \N__23857\,
            I => \b2v_inst11.un1_count_cry_11\
        );

    \I__4354\ : InMux
    port map (
            O => \N__23854\,
            I => \b2v_inst11.un1_count_cry_12\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__23851\,
            I => \N__23848\
        );

    \I__4352\ : InMux
    port map (
            O => \N__23848\,
            I => \N__23842\
        );

    \I__4351\ : InMux
    port map (
            O => \N__23847\,
            I => \N__23842\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__23842\,
            I => \N__23839\
        );

    \I__4349\ : Odrv4
    port map (
            O => \N__23839\,
            I => \b2v_inst11.un1_count_cry_13_c_RNI5AUZ0Z6\
        );

    \I__4348\ : InMux
    port map (
            O => \N__23836\,
            I => \b2v_inst11.un1_count_cry_13\
        );

    \I__4347\ : InMux
    port map (
            O => \N__23833\,
            I => \b2v_inst11.un1_count_cry_14\
        );

    \I__4346\ : CascadeMux
    port map (
            O => \N__23830\,
            I => \N__23827\
        );

    \I__4345\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23821\
        );

    \I__4344\ : InMux
    port map (
            O => \N__23826\,
            I => \N__23821\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__23821\,
            I => \N__23818\
        );

    \I__4342\ : Odrv4
    port map (
            O => \N__23818\,
            I => \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6\
        );

    \I__4341\ : CascadeMux
    port map (
            O => \N__23815\,
            I => \N__23811\
        );

    \I__4340\ : InMux
    port map (
            O => \N__23814\,
            I => \N__23806\
        );

    \I__4339\ : InMux
    port map (
            O => \N__23811\,
            I => \N__23806\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__23806\,
            I => \b2v_inst11.un1_count_cry_9_c_RNIQ23EZ0\
        );

    \I__4337\ : InMux
    port map (
            O => \N__23803\,
            I => \N__23800\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__23800\,
            I => \b2v_inst11.count_0_10\
        );

    \I__4335\ : InMux
    port map (
            O => \N__23797\,
            I => \N__23791\
        );

    \I__4334\ : InMux
    port map (
            O => \N__23796\,
            I => \N__23791\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__23791\,
            I => \b2v_inst11.un1_count_cry_10_c_RNI24RZ0Z6\
        );

    \I__4332\ : InMux
    port map (
            O => \N__23788\,
            I => \b2v_inst11.un1_count_cry_1\
        );

    \I__4331\ : InMux
    port map (
            O => \N__23785\,
            I => \b2v_inst11.un1_count_cry_2\
        );

    \I__4330\ : InMux
    port map (
            O => \N__23782\,
            I => \b2v_inst11.un1_count_cry_3\
        );

    \I__4329\ : InMux
    port map (
            O => \N__23779\,
            I => \b2v_inst11.un1_count_cry_4\
        );

    \I__4328\ : InMux
    port map (
            O => \N__23776\,
            I => \N__23770\
        );

    \I__4327\ : InMux
    port map (
            O => \N__23775\,
            I => \N__23770\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__23770\,
            I => \b2v_inst11.un1_count_cry_5_c_RNIMQUDZ0\
        );

    \I__4325\ : InMux
    port map (
            O => \N__23767\,
            I => \b2v_inst11.un1_count_cry_5\
        );

    \I__4324\ : InMux
    port map (
            O => \N__23764\,
            I => \N__23758\
        );

    \I__4323\ : InMux
    port map (
            O => \N__23763\,
            I => \N__23758\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__23758\,
            I => \b2v_inst11.un1_count_cry_6_c_RNINSVDZ0\
        );

    \I__4321\ : InMux
    port map (
            O => \N__23755\,
            I => \b2v_inst11.un1_count_cry_6\
        );

    \I__4320\ : InMux
    port map (
            O => \N__23752\,
            I => \b2v_inst11.un1_count_cry_7\
        );

    \I__4319\ : InMux
    port map (
            O => \N__23749\,
            I => \bfn_8_7_0_\
        );

    \I__4318\ : InMux
    port map (
            O => \N__23746\,
            I => \b2v_inst11.un1_count_cry_9\
        );

    \I__4317\ : InMux
    port map (
            O => \N__23743\,
            I => \N__23740\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__23740\,
            I => \b2v_inst11.count_0_14\
        );

    \I__4315\ : InMux
    port map (
            O => \N__23737\,
            I => \N__23734\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__23734\,
            I => \b2v_inst11.count_0_6\
        );

    \I__4313\ : InMux
    port map (
            O => \N__23731\,
            I => \N__23728\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__23728\,
            I => \b2v_inst11.count_0_15\
        );

    \I__4311\ : InMux
    port map (
            O => \N__23725\,
            I => \N__23722\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__23722\,
            I => \b2v_inst11.count_0_7\
        );

    \I__4309\ : CascadeMux
    port map (
            O => \N__23719\,
            I => \N__23715\
        );

    \I__4308\ : InMux
    port map (
            O => \N__23718\,
            I => \N__23710\
        );

    \I__4307\ : InMux
    port map (
            O => \N__23715\,
            I => \N__23702\
        );

    \I__4306\ : InMux
    port map (
            O => \N__23714\,
            I => \N__23702\
        );

    \I__4305\ : InMux
    port map (
            O => \N__23713\,
            I => \N__23702\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__23710\,
            I => \N__23699\
        );

    \I__4303\ : InMux
    port map (
            O => \N__23709\,
            I => \N__23696\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__23702\,
            I => \b2v_inst11.mult1_un145_sum_s_8\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__23699\,
            I => \b2v_inst11.mult1_un145_sum_s_8\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__23696\,
            I => \b2v_inst11.mult1_un145_sum_s_8\
        );

    \I__4299\ : CascadeMux
    port map (
            O => \N__23689\,
            I => \N__23685\
        );

    \I__4298\ : InMux
    port map (
            O => \N__23688\,
            I => \N__23677\
        );

    \I__4297\ : InMux
    port map (
            O => \N__23685\,
            I => \N__23677\
        );

    \I__4296\ : InMux
    port map (
            O => \N__23684\,
            I => \N__23677\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__23677\,
            I => \b2v_inst11.mult1_un145_sum_i_0_8\
        );

    \I__4294\ : InMux
    port map (
            O => \N__23674\,
            I => \b2v_inst11.mult1_un159_sum_cry_1\
        );

    \I__4293\ : InMux
    port map (
            O => \N__23671\,
            I => \N__23668\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__23668\,
            I => \b2v_inst11.mult1_un152_sum_cry_3_s\
        );

    \I__4291\ : InMux
    port map (
            O => \N__23665\,
            I => \b2v_inst11.mult1_un159_sum_cry_2\
        );

    \I__4290\ : CascadeMux
    port map (
            O => \N__23662\,
            I => \N__23659\
        );

    \I__4289\ : InMux
    port map (
            O => \N__23659\,
            I => \N__23656\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__23656\,
            I => \b2v_inst11.mult1_un152_sum_cry_4_s\
        );

    \I__4287\ : InMux
    port map (
            O => \N__23653\,
            I => \b2v_inst11.mult1_un159_sum_cry_3\
        );

    \I__4286\ : InMux
    port map (
            O => \N__23650\,
            I => \N__23647\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__23647\,
            I => \b2v_inst11.mult1_un152_sum_cry_5_s\
        );

    \I__4284\ : InMux
    port map (
            O => \N__23644\,
            I => \b2v_inst11.mult1_un159_sum_cry_4\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__23641\,
            I => \N__23638\
        );

    \I__4282\ : InMux
    port map (
            O => \N__23638\,
            I => \N__23635\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__23635\,
            I => \b2v_inst11.mult1_un152_sum_cry_6_s\
        );

    \I__4280\ : InMux
    port map (
            O => \N__23632\,
            I => \b2v_inst11.mult1_un159_sum_cry_5\
        );

    \I__4279\ : InMux
    port map (
            O => \N__23629\,
            I => \N__23626\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__23626\,
            I => \b2v_inst11.mult1_un159_sum_axb_7\
        );

    \I__4277\ : InMux
    port map (
            O => \N__23623\,
            I => \b2v_inst11.mult1_un159_sum_cry_6\
        );

    \I__4276\ : CascadeMux
    port map (
            O => \N__23620\,
            I => \N__23616\
        );

    \I__4275\ : InMux
    port map (
            O => \N__23619\,
            I => \N__23610\
        );

    \I__4274\ : InMux
    port map (
            O => \N__23616\,
            I => \N__23603\
        );

    \I__4273\ : InMux
    port map (
            O => \N__23615\,
            I => \N__23603\
        );

    \I__4272\ : InMux
    port map (
            O => \N__23614\,
            I => \N__23603\
        );

    \I__4271\ : InMux
    port map (
            O => \N__23613\,
            I => \N__23600\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__23610\,
            I => \b2v_inst11.mult1_un152_sum_s_8\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__23603\,
            I => \b2v_inst11.mult1_un152_sum_s_8\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__23600\,
            I => \b2v_inst11.mult1_un152_sum_s_8\
        );

    \I__4267\ : CascadeMux
    port map (
            O => \N__23593\,
            I => \N__23589\
        );

    \I__4266\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23581\
        );

    \I__4265\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23581\
        );

    \I__4264\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23581\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__23581\,
            I => \b2v_inst11.mult1_un152_sum_i_0_8\
        );

    \I__4262\ : CascadeMux
    port map (
            O => \N__23578\,
            I => \b2v_inst36.countZ0Z_10_cascade_\
        );

    \I__4261\ : InMux
    port map (
            O => \N__23575\,
            I => \N__23572\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__23572\,
            I => \b2v_inst36.count_1_10\
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__23569\,
            I => \N__23566\
        );

    \I__4258\ : InMux
    port map (
            O => \N__23566\,
            I => \N__23563\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__23563\,
            I => \N__23560\
        );

    \I__4256\ : Odrv4
    port map (
            O => \N__23560\,
            I => \b2v_inst11.mult1_un145_sum_i\
        );

    \I__4255\ : InMux
    port map (
            O => \N__23557\,
            I => \b2v_inst11.mult1_un152_sum_cry_2\
        );

    \I__4254\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23551\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__23551\,
            I => \b2v_inst11.mult1_un145_sum_cry_3_s\
        );

    \I__4252\ : InMux
    port map (
            O => \N__23548\,
            I => \b2v_inst11.mult1_un152_sum_cry_3\
        );

    \I__4251\ : CascadeMux
    port map (
            O => \N__23545\,
            I => \N__23542\
        );

    \I__4250\ : InMux
    port map (
            O => \N__23542\,
            I => \N__23539\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__23539\,
            I => \b2v_inst11.mult1_un145_sum_cry_4_s\
        );

    \I__4248\ : InMux
    port map (
            O => \N__23536\,
            I => \b2v_inst11.mult1_un152_sum_cry_4\
        );

    \I__4247\ : InMux
    port map (
            O => \N__23533\,
            I => \N__23530\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__23530\,
            I => \b2v_inst11.mult1_un145_sum_cry_5_s\
        );

    \I__4245\ : InMux
    port map (
            O => \N__23527\,
            I => \b2v_inst11.mult1_un152_sum_cry_5\
        );

    \I__4244\ : CascadeMux
    port map (
            O => \N__23524\,
            I => \N__23521\
        );

    \I__4243\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23518\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__23518\,
            I => \N__23515\
        );

    \I__4241\ : Odrv4
    port map (
            O => \N__23515\,
            I => \b2v_inst11.mult1_un145_sum_cry_6_s\
        );

    \I__4240\ : InMux
    port map (
            O => \N__23512\,
            I => \b2v_inst11.mult1_un152_sum_cry_6\
        );

    \I__4239\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23506\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__23506\,
            I => \b2v_inst11.mult1_un152_sum_axb_8\
        );

    \I__4237\ : InMux
    port map (
            O => \N__23503\,
            I => \b2v_inst11.mult1_un152_sum_cry_7\
        );

    \I__4236\ : CascadeMux
    port map (
            O => \N__23500\,
            I => \b2v_inst36.count_rst_9_cascade_\
        );

    \I__4235\ : CascadeMux
    port map (
            O => \N__23497\,
            I => \b2v_inst36.countZ0Z_5_cascade_\
        );

    \I__4234\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23491\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__23491\,
            I => \b2v_inst36.count_1_5\
        );

    \I__4232\ : InMux
    port map (
            O => \N__23488\,
            I => \N__23485\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__23485\,
            I => \b2v_inst36.count_rst_7\
        );

    \I__4230\ : CascadeMux
    port map (
            O => \N__23482\,
            I => \b2v_inst36.count_rst_6_cascade_\
        );

    \I__4229\ : CascadeMux
    port map (
            O => \N__23479\,
            I => \b2v_inst36.countZ0Z_8_cascade_\
        );

    \I__4228\ : InMux
    port map (
            O => \N__23476\,
            I => \N__23473\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__23473\,
            I => \b2v_inst36.count_1_8\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__23470\,
            I => \b2v_inst36.count_rst_4_cascade_\
        );

    \I__4225\ : InMux
    port map (
            O => \N__23467\,
            I => \N__23463\
        );

    \I__4224\ : InMux
    port map (
            O => \N__23466\,
            I => \N__23460\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__23463\,
            I => \b2v_inst11.func_state_RNI_0Z0Z_0\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__23460\,
            I => \b2v_inst11.func_state_RNI_0Z0Z_0\
        );

    \I__4221\ : InMux
    port map (
            O => \N__23455\,
            I => \N__23452\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__23452\,
            I => \b2v_inst11.g1_1\
        );

    \I__4219\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23443\
        );

    \I__4218\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23443\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__23443\,
            I => \b2v_inst11.func_state_RNI673P9Z0Z_0\
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__23440\,
            I => \N__23436\
        );

    \I__4215\ : InMux
    port map (
            O => \N__23439\,
            I => \N__23431\
        );

    \I__4214\ : InMux
    port map (
            O => \N__23436\,
            I => \N__23431\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__23431\,
            I => \b2v_inst11.func_stateZ1Z_0\
        );

    \I__4212\ : CascadeMux
    port map (
            O => \N__23428\,
            I => \N__23424\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__23427\,
            I => \N__23419\
        );

    \I__4210\ : InMux
    port map (
            O => \N__23424\,
            I => \N__23416\
        );

    \I__4209\ : InMux
    port map (
            O => \N__23423\,
            I => \N__23409\
        );

    \I__4208\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23409\
        );

    \I__4207\ : InMux
    port map (
            O => \N__23419\,
            I => \N__23406\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__23416\,
            I => \N__23403\
        );

    \I__4205\ : InMux
    port map (
            O => \N__23415\,
            I => \N__23398\
        );

    \I__4204\ : InMux
    port map (
            O => \N__23414\,
            I => \N__23398\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__23409\,
            I => \N__23395\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__23406\,
            I => \b2v_inst11.count_off_RNIZ0Z_9\
        );

    \I__4201\ : Odrv4
    port map (
            O => \N__23403\,
            I => \b2v_inst11.count_off_RNIZ0Z_9\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__23398\,
            I => \b2v_inst11.count_off_RNIZ0Z_9\
        );

    \I__4199\ : Odrv4
    port map (
            O => \N__23395\,
            I => \b2v_inst11.count_off_RNIZ0Z_9\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__23386\,
            I => \b2v_inst11.N_335_cascade_\
        );

    \I__4197\ : CascadeMux
    port map (
            O => \N__23383\,
            I => \N__23379\
        );

    \I__4196\ : CascadeMux
    port map (
            O => \N__23382\,
            I => \N__23371\
        );

    \I__4195\ : InMux
    port map (
            O => \N__23379\,
            I => \N__23368\
        );

    \I__4194\ : InMux
    port map (
            O => \N__23378\,
            I => \N__23365\
        );

    \I__4193\ : InMux
    port map (
            O => \N__23377\,
            I => \N__23360\
        );

    \I__4192\ : InMux
    port map (
            O => \N__23376\,
            I => \N__23360\
        );

    \I__4191\ : InMux
    port map (
            O => \N__23375\,
            I => \N__23355\
        );

    \I__4190\ : InMux
    port map (
            O => \N__23374\,
            I => \N__23355\
        );

    \I__4189\ : InMux
    port map (
            O => \N__23371\,
            I => \N__23352\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__23368\,
            I => \N__23347\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__23365\,
            I => \N__23347\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__23360\,
            I => \N__23344\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__23355\,
            I => \N__23333\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__23352\,
            I => \N__23333\
        );

    \I__4183\ : Span4Mux_s2_v
    port map (
            O => \N__23347\,
            I => \N__23333\
        );

    \I__4182\ : Span4Mux_s2_v
    port map (
            O => \N__23344\,
            I => \N__23330\
        );

    \I__4181\ : InMux
    port map (
            O => \N__23343\,
            I => \N__23327\
        );

    \I__4180\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23320\
        );

    \I__4179\ : InMux
    port map (
            O => \N__23341\,
            I => \N__23320\
        );

    \I__4178\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23320\
        );

    \I__4177\ : Span4Mux_h
    port map (
            O => \N__23333\,
            I => \N__23317\
        );

    \I__4176\ : Odrv4
    port map (
            O => \N__23330\,
            I => \b2v_inst11.count_off_RNIQ1RAS1Z0Z_9\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__23327\,
            I => \b2v_inst11.count_off_RNIQ1RAS1Z0Z_9\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__23320\,
            I => \b2v_inst11.count_off_RNIQ1RAS1Z0Z_9\
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__23317\,
            I => \b2v_inst11.count_off_RNIQ1RAS1Z0Z_9\
        );

    \I__4172\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23305\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__23305\,
            I => \b2v_inst11.func_state_1_ss0_i_0_o2_0\
        );

    \I__4170\ : CascadeMux
    port map (
            O => \N__23302\,
            I => \b2v_inst36.count_rst_11_cascade_\
        );

    \I__4169\ : CascadeMux
    port map (
            O => \N__23299\,
            I => \b2v_inst36.countZ0Z_7_cascade_\
        );

    \I__4168\ : InMux
    port map (
            O => \N__23296\,
            I => \N__23293\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__23293\,
            I => \b2v_inst36.count_1_7\
        );

    \I__4166\ : InMux
    port map (
            O => \N__23290\,
            I => \N__23287\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__23287\,
            I => \N__23281\
        );

    \I__4164\ : CascadeMux
    port map (
            O => \N__23286\,
            I => \N__23278\
        );

    \I__4163\ : CascadeMux
    port map (
            O => \N__23285\,
            I => \N__23275\
        );

    \I__4162\ : InMux
    port map (
            O => \N__23284\,
            I => \N__23272\
        );

    \I__4161\ : Span4Mux_h
    port map (
            O => \N__23281\,
            I => \N__23269\
        );

    \I__4160\ : InMux
    port map (
            O => \N__23278\,
            I => \N__23264\
        );

    \I__4159\ : InMux
    port map (
            O => \N__23275\,
            I => \N__23264\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__23272\,
            I => \N__23261\
        );

    \I__4157\ : Odrv4
    port map (
            O => \N__23269\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__23264\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\
        );

    \I__4155\ : Odrv12
    port map (
            O => \N__23261\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\
        );

    \I__4154\ : CascadeMux
    port map (
            O => \N__23254\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1_cascade_\
        );

    \I__4153\ : InMux
    port map (
            O => \N__23251\,
            I => \N__23248\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__23248\,
            I => \N__23245\
        );

    \I__4151\ : Odrv12
    port map (
            O => \N__23245\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_sx\
        );

    \I__4150\ : InMux
    port map (
            O => \N__23242\,
            I => \N__23239\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__23239\,
            I => \N__23235\
        );

    \I__4148\ : InMux
    port map (
            O => \N__23238\,
            I => \N__23232\
        );

    \I__4147\ : Sp12to4
    port map (
            O => \N__23235\,
            I => \N__23226\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__23232\,
            I => \N__23226\
        );

    \I__4145\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23223\
        );

    \I__4144\ : Span12Mux_s3_v
    port map (
            O => \N__23226\,
            I => \N__23220\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__23223\,
            I => \N__23217\
        );

    \I__4142\ : Odrv12
    port map (
            O => \N__23220\,
            I => \b2v_inst11.func_state_RNI_0Z0Z_1\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__23217\,
            I => \b2v_inst11.func_state_RNI_0Z0Z_1\
        );

    \I__4140\ : InMux
    port map (
            O => \N__23212\,
            I => \N__23209\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__23209\,
            I => \b2v_inst11.func_state_1_m0_0_0_1\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__23206\,
            I => \N__23201\
        );

    \I__4137\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23196\
        );

    \I__4136\ : InMux
    port map (
            O => \N__23204\,
            I => \N__23196\
        );

    \I__4135\ : InMux
    port map (
            O => \N__23201\,
            I => \N__23193\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__23196\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_0\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__23193\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_0\
        );

    \I__4132\ : InMux
    port map (
            O => \N__23188\,
            I => \N__23185\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__23185\,
            I => \N__23180\
        );

    \I__4130\ : CascadeMux
    port map (
            O => \N__23184\,
            I => \N__23177\
        );

    \I__4129\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23171\
        );

    \I__4128\ : Span4Mux_s2_v
    port map (
            O => \N__23180\,
            I => \N__23168\
        );

    \I__4127\ : InMux
    port map (
            O => \N__23177\,
            I => \N__23165\
        );

    \I__4126\ : InMux
    port map (
            O => \N__23176\,
            I => \N__23162\
        );

    \I__4125\ : InMux
    port map (
            O => \N__23175\,
            I => \N__23157\
        );

    \I__4124\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23157\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__23171\,
            I => \N__23154\
        );

    \I__4122\ : Odrv4
    port map (
            O => \N__23168\,
            I => \b2v_inst11.N_360\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__23165\,
            I => \b2v_inst11.N_360\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__23162\,
            I => \b2v_inst11.N_360\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__23157\,
            I => \b2v_inst11.N_360\
        );

    \I__4118\ : Odrv4
    port map (
            O => \N__23154\,
            I => \b2v_inst11.N_360\
        );

    \I__4117\ : InMux
    port map (
            O => \N__23143\,
            I => \N__23140\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__23140\,
            I => \N__23137\
        );

    \I__4115\ : Odrv12
    port map (
            O => \N__23137\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__23134\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_0_cascade_\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__23131\,
            I => \N__23128\
        );

    \I__4112\ : InMux
    port map (
            O => \N__23128\,
            I => \N__23122\
        );

    \I__4111\ : InMux
    port map (
            O => \N__23127\,
            I => \N__23122\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__23122\,
            I => \N__23118\
        );

    \I__4109\ : InMux
    port map (
            O => \N__23121\,
            I => \N__23115\
        );

    \I__4108\ : Span4Mux_v
    port map (
            O => \N__23118\,
            I => \N__23103\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__23115\,
            I => \N__23103\
        );

    \I__4106\ : InMux
    port map (
            O => \N__23114\,
            I => \N__23100\
        );

    \I__4105\ : InMux
    port map (
            O => \N__23113\,
            I => \N__23093\
        );

    \I__4104\ : InMux
    port map (
            O => \N__23112\,
            I => \N__23093\
        );

    \I__4103\ : InMux
    port map (
            O => \N__23111\,
            I => \N__23093\
        );

    \I__4102\ : InMux
    port map (
            O => \N__23110\,
            I => \N__23090\
        );

    \I__4101\ : InMux
    port map (
            O => \N__23109\,
            I => \N__23087\
        );

    \I__4100\ : InMux
    port map (
            O => \N__23108\,
            I => \N__23084\
        );

    \I__4099\ : Span4Mux_h
    port map (
            O => \N__23103\,
            I => \N__23077\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__23100\,
            I => \N__23077\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__23093\,
            I => \N__23077\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__23090\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__23087\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__23084\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__4093\ : Odrv4
    port map (
            O => \N__23077\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__4092\ : CascadeMux
    port map (
            O => \N__23068\,
            I => \b2v_inst11.func_stateZ0Z_0_cascade_\
        );

    \I__4091\ : CascadeMux
    port map (
            O => \N__23065\,
            I => \b2v_inst11.N_3013_i_cascade_\
        );

    \I__4090\ : InMux
    port map (
            O => \N__23062\,
            I => \N__23059\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__23059\,
            I => \b2v_inst11.N_330\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__23056\,
            I => \N__23050\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__23055\,
            I => \N__23047\
        );

    \I__4086\ : InMux
    port map (
            O => \N__23054\,
            I => \N__23044\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__23053\,
            I => \N__23040\
        );

    \I__4084\ : InMux
    port map (
            O => \N__23050\,
            I => \N__23037\
        );

    \I__4083\ : InMux
    port map (
            O => \N__23047\,
            I => \N__23034\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__23044\,
            I => \N__23031\
        );

    \I__4081\ : InMux
    port map (
            O => \N__23043\,
            I => \N__23028\
        );

    \I__4080\ : InMux
    port map (
            O => \N__23040\,
            I => \N__23025\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__23037\,
            I => \N__23020\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__23034\,
            I => \N__23020\
        );

    \I__4077\ : Span4Mux_v
    port map (
            O => \N__23031\,
            I => \N__23017\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__23028\,
            I => \N__23014\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__23025\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__4074\ : Odrv4
    port map (
            O => \N__23020\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__23017\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__4072\ : Odrv12
    port map (
            O => \N__23014\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__4071\ : CascadeMux
    port map (
            O => \N__23005\,
            I => \b2v_inst11.dutycycle_1_0_0_cascade_\
        );

    \I__4070\ : InMux
    port map (
            O => \N__23002\,
            I => \N__22999\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__22999\,
            I => \N__22996\
        );

    \I__4068\ : Span4Mux_h
    port map (
            O => \N__22996\,
            I => \N__22993\
        );

    \I__4067\ : Odrv4
    port map (
            O => \N__22993\,
            I => \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIZ0\
        );

    \I__4066\ : InMux
    port map (
            O => \N__22990\,
            I => \N__22987\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__22987\,
            I => \b2v_inst11.g1\
        );

    \I__4064\ : InMux
    port map (
            O => \N__22984\,
            I => \N__22978\
        );

    \I__4063\ : InMux
    port map (
            O => \N__22983\,
            I => \N__22978\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__22978\,
            I => \b2v_inst11.dutycycle_0_6\
        );

    \I__4061\ : CascadeMux
    port map (
            O => \N__22975\,
            I => \b2v_inst11.g1_cascade_\
        );

    \I__4060\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22968\
        );

    \I__4059\ : InMux
    port map (
            O => \N__22971\,
            I => \N__22965\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__22968\,
            I => \b2v_inst11.g1_0\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__22965\,
            I => \b2v_inst11.g1_0\
        );

    \I__4056\ : InMux
    port map (
            O => \N__22960\,
            I => \N__22957\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__22957\,
            I => \N__22954\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__22954\,
            I => \b2v_inst11.dutycycle_eena\
        );

    \I__4053\ : InMux
    port map (
            O => \N__22951\,
            I => \N__22948\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__22948\,
            I => \b2v_inst11.dutycycle_1_0_0\
        );

    \I__4051\ : CascadeMux
    port map (
            O => \N__22945\,
            I => \b2v_inst11.dutycycle_eena_cascade_\
        );

    \I__4050\ : InMux
    port map (
            O => \N__22942\,
            I => \N__22936\
        );

    \I__4049\ : InMux
    port map (
            O => \N__22941\,
            I => \N__22936\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__22936\,
            I => \b2v_inst11.dutycycleZ1Z_0\
        );

    \I__4047\ : CascadeMux
    port map (
            O => \N__22933\,
            I => \N__22930\
        );

    \I__4046\ : InMux
    port map (
            O => \N__22930\,
            I => \N__22924\
        );

    \I__4045\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22924\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__22924\,
            I => \N__22921\
        );

    \I__4043\ : Span4Mux_s2_h
    port map (
            O => \N__22921\,
            I => \N__22918\
        );

    \I__4042\ : Span4Mux_h
    port map (
            O => \N__22918\,
            I => \N__22915\
        );

    \I__4041\ : Odrv4
    port map (
            O => \N__22915\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3\
        );

    \I__4040\ : InMux
    port map (
            O => \N__22912\,
            I => \N__22909\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__22909\,
            I => \b2v_inst11.un1_clk_100khz_2_i_o3_out\
        );

    \I__4038\ : InMux
    port map (
            O => \N__22906\,
            I => \N__22903\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__22903\,
            I => \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8\
        );

    \I__4036\ : InMux
    port map (
            O => \N__22900\,
            I => \N__22897\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__22897\,
            I => \b2v_inst11.dutycycle_1_0_1\
        );

    \I__4034\ : InMux
    port map (
            O => \N__22894\,
            I => \N__22888\
        );

    \I__4033\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22888\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__22888\,
            I => \b2v_inst11.dutycycleZ1Z_1\
        );

    \I__4031\ : CascadeMux
    port map (
            O => \N__22885\,
            I => \b2v_inst11.dutycycle_1_0_1_cascade_\
        );

    \I__4030\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22879\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__22879\,
            I => \N__22876\
        );

    \I__4028\ : Span4Mux_s3_v
    port map (
            O => \N__22876\,
            I => \N__22872\
        );

    \I__4027\ : InMux
    port map (
            O => \N__22875\,
            I => \N__22869\
        );

    \I__4026\ : Span4Mux_h
    port map (
            O => \N__22872\,
            I => \N__22866\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__22869\,
            I => \N__22863\
        );

    \I__4024\ : Span4Mux_h
    port map (
            O => \N__22866\,
            I => \N__22860\
        );

    \I__4023\ : Span4Mux_h
    port map (
            O => \N__22863\,
            I => \N__22857\
        );

    \I__4022\ : Odrv4
    port map (
            O => \N__22860\,
            I => \b2v_inst11.func_state_RNI_1Z0Z_0\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__22857\,
            I => \b2v_inst11.func_state_RNI_1Z0Z_0\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__22852\,
            I => \b2v_inst11.func_state_RNI_0Z0Z_1_cascade_\
        );

    \I__4019\ : CascadeMux
    port map (
            O => \N__22849\,
            I => \b2v_inst11.un1_func_state25_4_i_a2_1_cascade_\
        );

    \I__4018\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22843\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__22843\,
            I => \N__22840\
        );

    \I__4016\ : Span4Mux_s2_h
    port map (
            O => \N__22840\,
            I => \N__22837\
        );

    \I__4015\ : Span4Mux_h
    port map (
            O => \N__22837\,
            I => \N__22834\
        );

    \I__4014\ : Odrv4
    port map (
            O => \N__22834\,
            I => \b2v_inst11.N_321\
        );

    \I__4013\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22828\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__22828\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_3\
        );

    \I__4011\ : InMux
    port map (
            O => \N__22825\,
            I => \N__22819\
        );

    \I__4010\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22819\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__22819\,
            I => \N__22816\
        );

    \I__4008\ : Odrv4
    port map (
            O => \N__22816\,
            I => \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__22813\,
            I => \N__22810\
        );

    \I__4006\ : InMux
    port map (
            O => \N__22810\,
            I => \N__22804\
        );

    \I__4005\ : InMux
    port map (
            O => \N__22809\,
            I => \N__22804\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__22804\,
            I => \b2v_inst11.dutycycle_e_1_3\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__22801\,
            I => \N__22797\
        );

    \I__4002\ : InMux
    port map (
            O => \N__22800\,
            I => \N__22792\
        );

    \I__4001\ : InMux
    port map (
            O => \N__22797\,
            I => \N__22792\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__22792\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__22789\,
            I => \b2v_inst11.dutycycleZ0Z_6_cascade_\
        );

    \I__3998\ : InMux
    port map (
            O => \N__22786\,
            I => \N__22780\
        );

    \I__3997\ : InMux
    port map (
            O => \N__22785\,
            I => \N__22768\
        );

    \I__3996\ : InMux
    port map (
            O => \N__22784\,
            I => \N__22765\
        );

    \I__3995\ : CascadeMux
    port map (
            O => \N__22783\,
            I => \N__22758\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__22780\,
            I => \N__22755\
        );

    \I__3993\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22750\
        );

    \I__3992\ : InMux
    port map (
            O => \N__22778\,
            I => \N__22750\
        );

    \I__3991\ : InMux
    port map (
            O => \N__22777\,
            I => \N__22743\
        );

    \I__3990\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22743\
        );

    \I__3989\ : InMux
    port map (
            O => \N__22775\,
            I => \N__22743\
        );

    \I__3988\ : InMux
    port map (
            O => \N__22774\,
            I => \N__22738\
        );

    \I__3987\ : InMux
    port map (
            O => \N__22773\,
            I => \N__22738\
        );

    \I__3986\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22735\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__22771\,
            I => \N__22730\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__22768\,
            I => \N__22722\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__22765\,
            I => \N__22719\
        );

    \I__3982\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22716\
        );

    \I__3981\ : InMux
    port map (
            O => \N__22763\,
            I => \N__22711\
        );

    \I__3980\ : InMux
    port map (
            O => \N__22762\,
            I => \N__22711\
        );

    \I__3979\ : InMux
    port map (
            O => \N__22761\,
            I => \N__22708\
        );

    \I__3978\ : InMux
    port map (
            O => \N__22758\,
            I => \N__22705\
        );

    \I__3977\ : Span4Mux_h
    port map (
            O => \N__22755\,
            I => \N__22702\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__22750\,
            I => \N__22699\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__22743\,
            I => \N__22692\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__22738\,
            I => \N__22692\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__22735\,
            I => \N__22692\
        );

    \I__3972\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22681\
        );

    \I__3971\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22681\
        );

    \I__3970\ : InMux
    port map (
            O => \N__22730\,
            I => \N__22681\
        );

    \I__3969\ : InMux
    port map (
            O => \N__22729\,
            I => \N__22681\
        );

    \I__3968\ : InMux
    port map (
            O => \N__22728\,
            I => \N__22681\
        );

    \I__3967\ : InMux
    port map (
            O => \N__22727\,
            I => \N__22674\
        );

    \I__3966\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22674\
        );

    \I__3965\ : InMux
    port map (
            O => \N__22725\,
            I => \N__22674\
        );

    \I__3964\ : Span4Mux_h
    port map (
            O => \N__22722\,
            I => \N__22669\
        );

    \I__3963\ : Span4Mux_h
    port map (
            O => \N__22719\,
            I => \N__22669\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__22716\,
            I => \N__22664\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__22711\,
            I => \N__22664\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__22708\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__22705\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3958\ : Odrv4
    port map (
            O => \N__22702\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__22699\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3956\ : Odrv4
    port map (
            O => \N__22692\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__22681\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__22674\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__22669\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3952\ : Odrv12
    port map (
            O => \N__22664\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__3951\ : InMux
    port map (
            O => \N__22645\,
            I => \N__22642\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__22642\,
            I => \N__22639\
        );

    \I__3949\ : Odrv4
    port map (
            O => \N__22639\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_3\
        );

    \I__3948\ : CascadeMux
    port map (
            O => \N__22636\,
            I => \b2v_inst11.func_state_RNINJ641_0Z0Z_1_cascade_\
        );

    \I__3947\ : CascadeMux
    port map (
            O => \N__22633\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1_cascade_\
        );

    \I__3946\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22627\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__22627\,
            I => \b2v_inst11.g0_2_3\
        );

    \I__3944\ : InMux
    port map (
            O => \N__22624\,
            I => \N__22621\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__22621\,
            I => \N__22618\
        );

    \I__3942\ : Odrv4
    port map (
            O => \N__22618\,
            I => \b2v_inst11.g0_2_2\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__22615\,
            I => \N__22612\
        );

    \I__3940\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22609\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__22609\,
            I => \N__22606\
        );

    \I__3938\ : Odrv4
    port map (
            O => \N__22606\,
            I => \b2v_inst11.g0_1_1_0\
        );

    \I__3937\ : CascadeMux
    port map (
            O => \N__22603\,
            I => \N__22600\
        );

    \I__3936\ : InMux
    port map (
            O => \N__22600\,
            I => \N__22597\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__22597\,
            I => \N__22594\
        );

    \I__3934\ : Span4Mux_s3_v
    port map (
            O => \N__22594\,
            I => \N__22589\
        );

    \I__3933\ : InMux
    port map (
            O => \N__22593\,
            I => \N__22581\
        );

    \I__3932\ : InMux
    port map (
            O => \N__22592\,
            I => \N__22578\
        );

    \I__3931\ : Span4Mux_h
    port map (
            O => \N__22589\,
            I => \N__22574\
        );

    \I__3930\ : InMux
    port map (
            O => \N__22588\,
            I => \N__22567\
        );

    \I__3929\ : InMux
    port map (
            O => \N__22587\,
            I => \N__22567\
        );

    \I__3928\ : InMux
    port map (
            O => \N__22586\,
            I => \N__22567\
        );

    \I__3927\ : InMux
    port map (
            O => \N__22585\,
            I => \N__22562\
        );

    \I__3926\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22562\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__22581\,
            I => \N__22557\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__22578\,
            I => \N__22557\
        );

    \I__3923\ : CascadeMux
    port map (
            O => \N__22577\,
            I => \N__22554\
        );

    \I__3922\ : Span4Mux_v
    port map (
            O => \N__22574\,
            I => \N__22550\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__22567\,
            I => \N__22547\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__22562\,
            I => \N__22542\
        );

    \I__3919\ : Span4Mux_h
    port map (
            O => \N__22557\,
            I => \N__22542\
        );

    \I__3918\ : InMux
    port map (
            O => \N__22554\,
            I => \N__22537\
        );

    \I__3917\ : InMux
    port map (
            O => \N__22553\,
            I => \N__22537\
        );

    \I__3916\ : Odrv4
    port map (
            O => \N__22550\,
            I => \b2v_inst11.func_state_RNIJU083Z0Z_0\
        );

    \I__3915\ : Odrv12
    port map (
            O => \N__22547\,
            I => \b2v_inst11.func_state_RNIJU083Z0Z_0\
        );

    \I__3914\ : Odrv4
    port map (
            O => \N__22542\,
            I => \b2v_inst11.func_state_RNIJU083Z0Z_0\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__22537\,
            I => \b2v_inst11.func_state_RNIJU083Z0Z_0\
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__22528\,
            I => \b2v_inst11.un1_clk_100khz_43_and_i_o2_0_0_1_cascade_\
        );

    \I__3911\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22522\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__22522\,
            I => \N__22519\
        );

    \I__3909\ : Span4Mux_h
    port map (
            O => \N__22519\,
            I => \N__22516\
        );

    \I__3908\ : Odrv4
    port map (
            O => \N__22516\,
            I => \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJTZ0Z69\
        );

    \I__3907\ : InMux
    port map (
            O => \N__22513\,
            I => \N__22510\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__22510\,
            I => \b2v_inst11.dutycycle_RNI4I3C2Z0Z_10\
        );

    \I__3905\ : CascadeMux
    port map (
            O => \N__22507\,
            I => \b2v_inst11.dutycycle_RNI4I3C2Z0Z_10_cascade_\
        );

    \I__3904\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22501\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__22501\,
            I => \b2v_inst11.dutycycle_RNIAI7C4Z0Z_10\
        );

    \I__3902\ : CascadeMux
    port map (
            O => \N__22498\,
            I => \N__22494\
        );

    \I__3901\ : InMux
    port map (
            O => \N__22497\,
            I => \N__22486\
        );

    \I__3900\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22486\
        );

    \I__3899\ : InMux
    port map (
            O => \N__22493\,
            I => \N__22486\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__22486\,
            I => \b2v_inst11.dutycycleZ1Z_10\
        );

    \I__3897\ : CascadeMux
    port map (
            O => \N__22483\,
            I => \N__22480\
        );

    \I__3896\ : InMux
    port map (
            O => \N__22480\,
            I => \N__22477\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__22477\,
            I => \N__22474\
        );

    \I__3894\ : Span4Mux_h
    port map (
            O => \N__22474\,
            I => \N__22471\
        );

    \I__3893\ : Odrv4
    port map (
            O => \N__22471\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_5\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__22468\,
            I => \b2v_inst11.d_i3_mux_cascade_\
        );

    \I__3891\ : InMux
    port map (
            O => \N__22465\,
            I => \N__22462\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__22462\,
            I => \N__22459\
        );

    \I__3889\ : Span4Mux_h
    port map (
            O => \N__22459\,
            I => \N__22456\
        );

    \I__3888\ : Odrv4
    port map (
            O => \N__22456\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_5\
        );

    \I__3887\ : CascadeMux
    port map (
            O => \N__22453\,
            I => \N__22450\
        );

    \I__3886\ : InMux
    port map (
            O => \N__22450\,
            I => \N__22447\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__22447\,
            I => \N__22443\
        );

    \I__3884\ : InMux
    port map (
            O => \N__22446\,
            I => \N__22440\
        );

    \I__3883\ : Span4Mux_h
    port map (
            O => \N__22443\,
            I => \N__22437\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__22440\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_3\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__22437\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_3\
        );

    \I__3880\ : InMux
    port map (
            O => \N__22432\,
            I => \N__22429\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__22429\,
            I => \b2v_inst11.curr_state_0_0\
        );

    \I__3878\ : InMux
    port map (
            O => \N__22426\,
            I => \N__22423\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__22423\,
            I => \b2v_inst11.curr_state_3_0\
        );

    \I__3876\ : CascadeMux
    port map (
            O => \N__22420\,
            I => \b2v_inst11.curr_stateZ0Z_0_cascade_\
        );

    \I__3875\ : CascadeMux
    port map (
            O => \N__22417\,
            I => \b2v_inst11.count_0_sqmuxa_i_cascade_\
        );

    \I__3874\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22411\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__22411\,
            I => \N__22408\
        );

    \I__3872\ : Span4Mux_v
    port map (
            O => \N__22408\,
            I => \N__22405\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__22405\,
            I => \b2v_inst11.N_349\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__22402\,
            I => \N__22397\
        );

    \I__3869\ : InMux
    port map (
            O => \N__22401\,
            I => \N__22393\
        );

    \I__3868\ : InMux
    port map (
            O => \N__22400\,
            I => \N__22386\
        );

    \I__3867\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22386\
        );

    \I__3866\ : InMux
    port map (
            O => \N__22396\,
            I => \N__22386\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__22393\,
            I => \N__22383\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__22386\,
            I => \N__22380\
        );

    \I__3863\ : Span4Mux_h
    port map (
            O => \N__22383\,
            I => \N__22377\
        );

    \I__3862\ : Span4Mux_v
    port map (
            O => \N__22380\,
            I => \N__22374\
        );

    \I__3861\ : Span4Mux_h
    port map (
            O => \N__22377\,
            I => \N__22371\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__22374\,
            I => \b2v_inst11.un1_clk_100khz_32_and_i_o2_0_0_1\
        );

    \I__3859\ : Odrv4
    port map (
            O => \N__22371\,
            I => \b2v_inst11.un1_clk_100khz_32_and_i_o2_0_0_1\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__22366\,
            I => \b2v_inst11.dutycycle_RNIAI7C4Z0Z_10_cascade_\
        );

    \I__3857\ : CascadeMux
    port map (
            O => \N__22363\,
            I => \N__22356\
        );

    \I__3856\ : CascadeMux
    port map (
            O => \N__22362\,
            I => \N__22351\
        );

    \I__3855\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22342\
        );

    \I__3854\ : InMux
    port map (
            O => \N__22360\,
            I => \N__22337\
        );

    \I__3853\ : InMux
    port map (
            O => \N__22359\,
            I => \N__22337\
        );

    \I__3852\ : InMux
    port map (
            O => \N__22356\,
            I => \N__22334\
        );

    \I__3851\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22331\
        );

    \I__3850\ : InMux
    port map (
            O => \N__22354\,
            I => \N__22324\
        );

    \I__3849\ : InMux
    port map (
            O => \N__22351\,
            I => \N__22324\
        );

    \I__3848\ : InMux
    port map (
            O => \N__22350\,
            I => \N__22324\
        );

    \I__3847\ : InMux
    port map (
            O => \N__22349\,
            I => \N__22321\
        );

    \I__3846\ : InMux
    port map (
            O => \N__22348\,
            I => \N__22318\
        );

    \I__3845\ : InMux
    port map (
            O => \N__22347\,
            I => \N__22311\
        );

    \I__3844\ : InMux
    port map (
            O => \N__22346\,
            I => \N__22311\
        );

    \I__3843\ : InMux
    port map (
            O => \N__22345\,
            I => \N__22311\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__22342\,
            I => \N__22305\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__22337\,
            I => \N__22302\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__22334\,
            I => \N__22295\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__22331\,
            I => \N__22295\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__22324\,
            I => \N__22295\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__22321\,
            I => \N__22288\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__22318\,
            I => \N__22288\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__22311\,
            I => \N__22288\
        );

    \I__3834\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22284\
        );

    \I__3833\ : InMux
    port map (
            O => \N__22309\,
            I => \N__22279\
        );

    \I__3832\ : InMux
    port map (
            O => \N__22308\,
            I => \N__22279\
        );

    \I__3831\ : Span4Mux_h
    port map (
            O => \N__22305\,
            I => \N__22276\
        );

    \I__3830\ : Span4Mux_h
    port map (
            O => \N__22302\,
            I => \N__22269\
        );

    \I__3829\ : Span4Mux_v
    port map (
            O => \N__22295\,
            I => \N__22269\
        );

    \I__3828\ : Span4Mux_v
    port map (
            O => \N__22288\,
            I => \N__22269\
        );

    \I__3827\ : InMux
    port map (
            O => \N__22287\,
            I => \N__22266\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__22284\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__22279\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__3824\ : Odrv4
    port map (
            O => \N__22276\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__3823\ : Odrv4
    port map (
            O => \N__22269\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__22266\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__3821\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22250\
        );

    \I__3820\ : InMux
    port map (
            O => \N__22254\,
            I => \N__22245\
        );

    \I__3819\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22245\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__22250\,
            I => \N__22233\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__22245\,
            I => \N__22233\
        );

    \I__3816\ : InMux
    port map (
            O => \N__22244\,
            I => \N__22228\
        );

    \I__3815\ : InMux
    port map (
            O => \N__22243\,
            I => \N__22228\
        );

    \I__3814\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22224\
        );

    \I__3813\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22221\
        );

    \I__3812\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22216\
        );

    \I__3811\ : InMux
    port map (
            O => \N__22239\,
            I => \N__22216\
        );

    \I__3810\ : InMux
    port map (
            O => \N__22238\,
            I => \N__22213\
        );

    \I__3809\ : Span4Mux_v
    port map (
            O => \N__22233\,
            I => \N__22210\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__22228\,
            I => \N__22207\
        );

    \I__3807\ : InMux
    port map (
            O => \N__22227\,
            I => \N__22204\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__22224\,
            I => \N__22199\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__22221\,
            I => \N__22199\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__22216\,
            I => \N__22194\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__22213\,
            I => \N__22194\
        );

    \I__3802\ : Span4Mux_v
    port map (
            O => \N__22210\,
            I => \N__22191\
        );

    \I__3801\ : Span4Mux_v
    port map (
            O => \N__22207\,
            I => \N__22188\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__22204\,
            I => \N__22181\
        );

    \I__3799\ : Span4Mux_v
    port map (
            O => \N__22199\,
            I => \N__22181\
        );

    \I__3798\ : Span4Mux_h
    port map (
            O => \N__22194\,
            I => \N__22181\
        );

    \I__3797\ : Odrv4
    port map (
            O => \N__22191\,
            I => \b2v_inst11.N_418\
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__22188\,
            I => \b2v_inst11.N_418\
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__22181\,
            I => \b2v_inst11.N_418\
        );

    \I__3794\ : CascadeMux
    port map (
            O => \N__22174\,
            I => \N__22171\
        );

    \I__3793\ : InMux
    port map (
            O => \N__22171\,
            I => \N__22168\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__22168\,
            I => \b2v_inst11.mult1_un61_sum_i_8\
        );

    \I__3791\ : InMux
    port map (
            O => \N__22165\,
            I => \N__22162\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__22162\,
            I => \b2v_inst11.N_5661_i\
        );

    \I__3789\ : InMux
    port map (
            O => \N__22159\,
            I => \bfn_7_7_0_\
        );

    \I__3788\ : InMux
    port map (
            O => \N__22156\,
            I => \N__22153\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__22153\,
            I => \N__22150\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__22150\,
            I => \b2v_inst36.curr_state_RNI8TT2Z0Z_0\
        );

    \I__3785\ : CascadeMux
    port map (
            O => \N__22147\,
            I => \b2v_inst11.pwm_out_en_cascade_\
        );

    \I__3784\ : IoInMux
    port map (
            O => \N__22144\,
            I => \N__22141\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__22141\,
            I => \N__22138\
        );

    \I__3782\ : Span4Mux_s0_v
    port map (
            O => \N__22138\,
            I => \N__22135\
        );

    \I__3781\ : Span4Mux_v
    port map (
            O => \N__22135\,
            I => \N__22132\
        );

    \I__3780\ : Span4Mux_v
    port map (
            O => \N__22132\,
            I => \N__22129\
        );

    \I__3779\ : Odrv4
    port map (
            O => \N__22129\,
            I => \PWRBTN_LED_c\
        );

    \I__3778\ : InMux
    port map (
            O => \N__22126\,
            I => \N__22123\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__22123\,
            I => \b2v_inst11.pwm_out_1_sqmuxa_0\
        );

    \I__3776\ : InMux
    port map (
            O => \N__22120\,
            I => \N__22117\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__22117\,
            I => \b2v_inst11.N_5653_i\
        );

    \I__3774\ : CascadeMux
    port map (
            O => \N__22114\,
            I => \N__22111\
        );

    \I__3773\ : InMux
    port map (
            O => \N__22111\,
            I => \N__22108\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__22108\,
            I => \b2v_inst11.un85_clk_100khz_8\
        );

    \I__3771\ : InMux
    port map (
            O => \N__22105\,
            I => \N__22102\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__22102\,
            I => \b2v_inst11.N_5654_i\
        );

    \I__3769\ : InMux
    port map (
            O => \N__22099\,
            I => \N__22096\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__22096\,
            I => \N__22093\
        );

    \I__3767\ : Span4Mux_v
    port map (
            O => \N__22093\,
            I => \N__22090\
        );

    \I__3766\ : Odrv4
    port map (
            O => \N__22090\,
            I => \b2v_inst11.un85_clk_100khz_9\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__22087\,
            I => \N__22084\
        );

    \I__3764\ : InMux
    port map (
            O => \N__22084\,
            I => \N__22081\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__22081\,
            I => \b2v_inst11.N_5655_i\
        );

    \I__3762\ : CascadeMux
    port map (
            O => \N__22078\,
            I => \N__22075\
        );

    \I__3761\ : InMux
    port map (
            O => \N__22075\,
            I => \N__22072\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__22072\,
            I => \b2v_inst11.un85_clk_100khz_10\
        );

    \I__3759\ : InMux
    port map (
            O => \N__22069\,
            I => \N__22066\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__22066\,
            I => \b2v_inst11.N_5656_i\
        );

    \I__3757\ : InMux
    port map (
            O => \N__22063\,
            I => \N__22060\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__22060\,
            I => \N__22057\
        );

    \I__3755\ : Span4Mux_v
    port map (
            O => \N__22057\,
            I => \N__22054\
        );

    \I__3754\ : Odrv4
    port map (
            O => \N__22054\,
            I => \b2v_inst11.un85_clk_100khz_11\
        );

    \I__3753\ : CascadeMux
    port map (
            O => \N__22051\,
            I => \N__22048\
        );

    \I__3752\ : InMux
    port map (
            O => \N__22048\,
            I => \N__22045\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__22045\,
            I => \b2v_inst11.N_5657_i\
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__22042\,
            I => \N__22039\
        );

    \I__3749\ : InMux
    port map (
            O => \N__22039\,
            I => \N__22036\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__22036\,
            I => \N__22033\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__22033\,
            I => \b2v_inst11.un85_clk_100khz_12\
        );

    \I__3746\ : InMux
    port map (
            O => \N__22030\,
            I => \N__22027\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__22027\,
            I => \b2v_inst11.N_5658_i\
        );

    \I__3744\ : InMux
    port map (
            O => \N__22024\,
            I => \N__22021\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__22021\,
            I => \b2v_inst11.un85_clk_100khz_13\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__22018\,
            I => \N__22015\
        );

    \I__3741\ : InMux
    port map (
            O => \N__22015\,
            I => \N__22012\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__22012\,
            I => \b2v_inst11.N_5659_i\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__22009\,
            I => \N__22006\
        );

    \I__3738\ : InMux
    port map (
            O => \N__22006\,
            I => \N__22003\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__22003\,
            I => \b2v_inst11.un85_clk_100khz_14\
        );

    \I__3736\ : InMux
    port map (
            O => \N__22000\,
            I => \N__21997\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__21997\,
            I => \b2v_inst11.N_5660_i\
        );

    \I__3734\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21991\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__21991\,
            I => \b2v_inst11.mult1_un131_sum_i\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__21988\,
            I => \N__21985\
        );

    \I__3731\ : InMux
    port map (
            O => \N__21985\,
            I => \N__21982\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__21982\,
            I => \N__21979\
        );

    \I__3729\ : Span4Mux_h
    port map (
            O => \N__21979\,
            I => \N__21976\
        );

    \I__3728\ : Odrv4
    port map (
            O => \N__21976\,
            I => \b2v_inst11.un1_count_cry_0_i\
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__21973\,
            I => \N__21970\
        );

    \I__3726\ : InMux
    port map (
            O => \N__21970\,
            I => \N__21967\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__21967\,
            I => \b2v_inst11.un85_clk_100khz_1\
        );

    \I__3724\ : InMux
    port map (
            O => \N__21964\,
            I => \N__21961\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__21961\,
            I => \b2v_inst11.N_5647_i\
        );

    \I__3722\ : InMux
    port map (
            O => \N__21958\,
            I => \N__21955\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__21955\,
            I => \b2v_inst11.un85_clk_100khz_2\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__21952\,
            I => \N__21949\
        );

    \I__3719\ : InMux
    port map (
            O => \N__21949\,
            I => \N__21946\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__21946\,
            I => \b2v_inst11.N_5648_i\
        );

    \I__3717\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21940\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__21940\,
            I => \b2v_inst11.un85_clk_100khz_3\
        );

    \I__3715\ : CascadeMux
    port map (
            O => \N__21937\,
            I => \N__21934\
        );

    \I__3714\ : InMux
    port map (
            O => \N__21934\,
            I => \N__21931\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__21931\,
            I => \N__21928\
        );

    \I__3712\ : Odrv12
    port map (
            O => \N__21928\,
            I => \b2v_inst11.N_5649_i\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__21925\,
            I => \N__21922\
        );

    \I__3710\ : InMux
    port map (
            O => \N__21922\,
            I => \N__21919\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__21919\,
            I => \N__21916\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__21916\,
            I => \b2v_inst11.un85_clk_100khz_4\
        );

    \I__3707\ : InMux
    port map (
            O => \N__21913\,
            I => \N__21910\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__21910\,
            I => \b2v_inst11.N_5650_i\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__21907\,
            I => \N__21904\
        );

    \I__3704\ : InMux
    port map (
            O => \N__21904\,
            I => \N__21901\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__21901\,
            I => \b2v_inst11.un85_clk_100khz_5\
        );

    \I__3702\ : InMux
    port map (
            O => \N__21898\,
            I => \N__21895\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__21895\,
            I => \b2v_inst11.N_5651_i\
        );

    \I__3700\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21889\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__21889\,
            I => \b2v_inst11.un85_clk_100khz_6\
        );

    \I__3698\ : CascadeMux
    port map (
            O => \N__21886\,
            I => \N__21883\
        );

    \I__3697\ : InMux
    port map (
            O => \N__21883\,
            I => \N__21880\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__21880\,
            I => \b2v_inst11.N_5652_i\
        );

    \I__3695\ : CascadeMux
    port map (
            O => \N__21877\,
            I => \N__21874\
        );

    \I__3694\ : InMux
    port map (
            O => \N__21874\,
            I => \N__21871\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__21871\,
            I => \b2v_inst11.un85_clk_100khz_7\
        );

    \I__3692\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21865\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__21865\,
            I => \b2v_inst11.mult1_un138_sum_axb_8\
        );

    \I__3690\ : InMux
    port map (
            O => \N__21862\,
            I => \b2v_inst11.mult1_un138_sum_cry_7\
        );

    \I__3689\ : CascadeMux
    port map (
            O => \N__21859\,
            I => \N__21856\
        );

    \I__3688\ : InMux
    port map (
            O => \N__21856\,
            I => \N__21846\
        );

    \I__3687\ : InMux
    port map (
            O => \N__21855\,
            I => \N__21846\
        );

    \I__3686\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21846\
        );

    \I__3685\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21843\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__21846\,
            I => \b2v_inst11.mult1_un138_sum_s_8\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__21843\,
            I => \b2v_inst11.mult1_un138_sum_s_8\
        );

    \I__3682\ : CascadeMux
    port map (
            O => \N__21838\,
            I => \b2v_inst11.mult1_un138_sum_s_8_cascade_\
        );

    \I__3681\ : InMux
    port map (
            O => \N__21835\,
            I => \N__21832\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__21832\,
            I => \N__21828\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__21831\,
            I => \N__21825\
        );

    \I__3678\ : Span4Mux_v
    port map (
            O => \N__21828\,
            I => \N__21819\
        );

    \I__3677\ : InMux
    port map (
            O => \N__21825\,
            I => \N__21812\
        );

    \I__3676\ : InMux
    port map (
            O => \N__21824\,
            I => \N__21812\
        );

    \I__3675\ : InMux
    port map (
            O => \N__21823\,
            I => \N__21812\
        );

    \I__3674\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21809\
        );

    \I__3673\ : Odrv4
    port map (
            O => \N__21819\,
            I => \b2v_inst11.mult1_un82_sum_s_8\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__21812\,
            I => \b2v_inst11.mult1_un82_sum_s_8\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__21809\,
            I => \b2v_inst11.mult1_un82_sum_s_8\
        );

    \I__3670\ : CascadeMux
    port map (
            O => \N__21802\,
            I => \N__21798\
        );

    \I__3669\ : InMux
    port map (
            O => \N__21801\,
            I => \N__21793\
        );

    \I__3668\ : InMux
    port map (
            O => \N__21798\,
            I => \N__21788\
        );

    \I__3667\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21788\
        );

    \I__3666\ : InMux
    port map (
            O => \N__21796\,
            I => \N__21785\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__21793\,
            I => \b2v_inst11.mult1_un131_sum_s_8\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__21788\,
            I => \b2v_inst11.mult1_un131_sum_s_8\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__21785\,
            I => \b2v_inst11.mult1_un131_sum_s_8\
        );

    \I__3662\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21775\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__21775\,
            I => \N__21771\
        );

    \I__3660\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21768\
        );

    \I__3659\ : Span4Mux_s2_v
    port map (
            O => \N__21771\,
            I => \N__21763\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__21768\,
            I => \N__21763\
        );

    \I__3657\ : Span4Mux_v
    port map (
            O => \N__21763\,
            I => \N__21760\
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__21760\,
            I => \b2v_inst11.mult1_un138_sum\
        );

    \I__3655\ : CascadeMux
    port map (
            O => \N__21757\,
            I => \N__21754\
        );

    \I__3654\ : InMux
    port map (
            O => \N__21754\,
            I => \N__21751\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__21751\,
            I => \N__21748\
        );

    \I__3652\ : Odrv4
    port map (
            O => \N__21748\,
            I => \b2v_inst11.mult1_un138_sum_i\
        );

    \I__3651\ : InMux
    port map (
            O => \N__21745\,
            I => \N__21741\
        );

    \I__3650\ : InMux
    port map (
            O => \N__21744\,
            I => \N__21738\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__21741\,
            I => \N__21735\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__21738\,
            I => \N__21732\
        );

    \I__3647\ : Span4Mux_h
    port map (
            O => \N__21735\,
            I => \N__21729\
        );

    \I__3646\ : Span4Mux_h
    port map (
            O => \N__21732\,
            I => \N__21726\
        );

    \I__3645\ : Odrv4
    port map (
            O => \N__21729\,
            I => \b2v_inst11.mult1_un131_sum\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__21726\,
            I => \b2v_inst11.mult1_un131_sum\
        );

    \I__3643\ : InMux
    port map (
            O => \N__21721\,
            I => \b2v_inst11.mult1_un145_sum_cry_7\
        );

    \I__3642\ : CascadeMux
    port map (
            O => \N__21718\,
            I => \N__21714\
        );

    \I__3641\ : InMux
    port map (
            O => \N__21717\,
            I => \N__21706\
        );

    \I__3640\ : InMux
    port map (
            O => \N__21714\,
            I => \N__21706\
        );

    \I__3639\ : InMux
    port map (
            O => \N__21713\,
            I => \N__21706\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__21706\,
            I => \b2v_inst11.mult1_un138_sum_i_0_8\
        );

    \I__3637\ : InMux
    port map (
            O => \N__21703\,
            I => \N__21700\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__21700\,
            I => \b2v_inst11.mult1_un138_sum_cry_3_s\
        );

    \I__3635\ : InMux
    port map (
            O => \N__21697\,
            I => \b2v_inst11.mult1_un138_sum_cry_2\
        );

    \I__3634\ : CascadeMux
    port map (
            O => \N__21694\,
            I => \N__21691\
        );

    \I__3633\ : InMux
    port map (
            O => \N__21691\,
            I => \N__21688\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__21688\,
            I => \b2v_inst11.mult1_un131_sum_cry_3_s\
        );

    \I__3631\ : CascadeMux
    port map (
            O => \N__21685\,
            I => \N__21682\
        );

    \I__3630\ : InMux
    port map (
            O => \N__21682\,
            I => \N__21679\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__21679\,
            I => \b2v_inst11.mult1_un138_sum_cry_4_s\
        );

    \I__3628\ : InMux
    port map (
            O => \N__21676\,
            I => \b2v_inst11.mult1_un138_sum_cry_3\
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__21673\,
            I => \N__21670\
        );

    \I__3626\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21667\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__21667\,
            I => \N__21664\
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__21664\,
            I => \b2v_inst11.mult1_un131_sum_cry_4_s\
        );

    \I__3623\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21658\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__21658\,
            I => \b2v_inst11.mult1_un138_sum_cry_5_s\
        );

    \I__3621\ : InMux
    port map (
            O => \N__21655\,
            I => \b2v_inst11.mult1_un138_sum_cry_4\
        );

    \I__3620\ : InMux
    port map (
            O => \N__21652\,
            I => \N__21649\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__21649\,
            I => \b2v_inst11.mult1_un131_sum_cry_5_s\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__21646\,
            I => \N__21643\
        );

    \I__3617\ : InMux
    port map (
            O => \N__21643\,
            I => \N__21640\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__21640\,
            I => \b2v_inst11.mult1_un138_sum_cry_6_s\
        );

    \I__3615\ : InMux
    port map (
            O => \N__21637\,
            I => \b2v_inst11.mult1_un138_sum_cry_5\
        );

    \I__3614\ : InMux
    port map (
            O => \N__21634\,
            I => \N__21631\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__21631\,
            I => \b2v_inst11.mult1_un131_sum_cry_6_s\
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__21628\,
            I => \N__21624\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__21627\,
            I => \N__21620\
        );

    \I__3610\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21613\
        );

    \I__3609\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21613\
        );

    \I__3608\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21613\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__21613\,
            I => \b2v_inst11.mult1_un131_sum_i_0_8\
        );

    \I__3606\ : InMux
    port map (
            O => \N__21610\,
            I => \N__21607\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__21607\,
            I => \b2v_inst11.mult1_un145_sum_axb_8\
        );

    \I__3604\ : InMux
    port map (
            O => \N__21604\,
            I => \b2v_inst11.mult1_un138_sum_cry_6\
        );

    \I__3603\ : InMux
    port map (
            O => \N__21601\,
            I => \N__21592\
        );

    \I__3602\ : InMux
    port map (
            O => \N__21600\,
            I => \N__21592\
        );

    \I__3601\ : InMux
    port map (
            O => \N__21599\,
            I => \N__21586\
        );

    \I__3600\ : InMux
    port map (
            O => \N__21598\,
            I => \N__21586\
        );

    \I__3599\ : InMux
    port map (
            O => \N__21597\,
            I => \N__21583\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__21592\,
            I => \N__21580\
        );

    \I__3597\ : InMux
    port map (
            O => \N__21591\,
            I => \N__21577\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__21586\,
            I => \N__21574\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__21583\,
            I => \N__21571\
        );

    \I__3594\ : Span4Mux_h
    port map (
            O => \N__21580\,
            I => \N__21568\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__21577\,
            I => \N__21563\
        );

    \I__3592\ : Span4Mux_v
    port map (
            O => \N__21574\,
            I => \N__21563\
        );

    \I__3591\ : Span4Mux_s3_h
    port map (
            O => \N__21571\,
            I => \N__21560\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__21568\,
            I => \b2v_inst11.func_state_RNI_1Z0Z_1\
        );

    \I__3589\ : Odrv4
    port map (
            O => \N__21563\,
            I => \b2v_inst11.func_state_RNI_1Z0Z_1\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__21560\,
            I => \b2v_inst11.func_state_RNI_1Z0Z_1\
        );

    \I__3587\ : InMux
    port map (
            O => \N__21553\,
            I => \N__21550\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__21550\,
            I => \b2v_inst11.func_state_1_m2s2_i_1\
        );

    \I__3585\ : InMux
    port map (
            O => \N__21547\,
            I => \N__21544\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__21544\,
            I => \b2v_inst11.N_73\
        );

    \I__3583\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21538\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__21538\,
            I => \b2v_inst11.func_state_1_m0_0\
        );

    \I__3581\ : CascadeMux
    port map (
            O => \N__21535\,
            I => \b2v_inst11.N_73_cascade_\
        );

    \I__3580\ : InMux
    port map (
            O => \N__21532\,
            I => \N__21529\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__21529\,
            I => \b2v_inst11.count_off_RNIQCBN4Z0Z_9\
        );

    \I__3578\ : InMux
    port map (
            O => \N__21526\,
            I => \N__21523\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__21523\,
            I => \b2v_inst11.func_state_1_m0_1\
        );

    \I__3576\ : InMux
    port map (
            O => \N__21520\,
            I => \b2v_inst11.mult1_un145_sum_cry_2\
        );

    \I__3575\ : InMux
    port map (
            O => \N__21517\,
            I => \b2v_inst11.mult1_un145_sum_cry_3\
        );

    \I__3574\ : InMux
    port map (
            O => \N__21514\,
            I => \b2v_inst11.mult1_un145_sum_cry_4\
        );

    \I__3573\ : InMux
    port map (
            O => \N__21511\,
            I => \b2v_inst11.mult1_un145_sum_cry_5\
        );

    \I__3572\ : InMux
    port map (
            O => \N__21508\,
            I => \b2v_inst11.mult1_un145_sum_cry_6\
        );

    \I__3571\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21502\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__21502\,
            I => \N__21499\
        );

    \I__3569\ : Span4Mux_h
    port map (
            O => \N__21499\,
            I => \N__21496\
        );

    \I__3568\ : Odrv4
    port map (
            O => \N__21496\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_307_N\
        );

    \I__3567\ : InMux
    port map (
            O => \N__21493\,
            I => \N__21489\
        );

    \I__3566\ : InMux
    port map (
            O => \N__21492\,
            I => \N__21486\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__21489\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_5\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__21486\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_5\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__21481\,
            I => \b2v_inst11.N_4_cascade_\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__21478\,
            I => \b2v_inst11.func_state_RNI_0Z0Z_0_cascade_\
        );

    \I__3561\ : InMux
    port map (
            O => \N__21475\,
            I => \N__21472\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__21472\,
            I => \b2v_inst11.func_state_RNINJ641_0Z0Z_0\
        );

    \I__3559\ : CascadeMux
    port map (
            O => \N__21469\,
            I => \b2v_inst11.func_state_RNINJ641_0Z0Z_0_cascade_\
        );

    \I__3558\ : CascadeMux
    port map (
            O => \N__21466\,
            I => \b2v_inst11.count_off_RNIQCBN4Z0Z_9_cascade_\
        );

    \I__3557\ : InMux
    port map (
            O => \N__21463\,
            I => \N__21460\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__21460\,
            I => \b2v_inst11.N_333\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__21457\,
            I => \N__21454\
        );

    \I__3554\ : InMux
    port map (
            O => \N__21454\,
            I => \N__21448\
        );

    \I__3553\ : InMux
    port map (
            O => \N__21453\,
            I => \N__21448\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__21448\,
            I => \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNPZ0Z5\
        );

    \I__3551\ : InMux
    port map (
            O => \N__21445\,
            I => \b2v_inst11.un1_dutycycle_94_cry_10\
        );

    \I__3550\ : InMux
    port map (
            O => \N__21442\,
            I => \N__21437\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__21441\,
            I => \N__21430\
        );

    \I__3548\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21427\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__21437\,
            I => \N__21424\
        );

    \I__3546\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21421\
        );

    \I__3545\ : InMux
    port map (
            O => \N__21435\,
            I => \N__21418\
        );

    \I__3544\ : InMux
    port map (
            O => \N__21434\,
            I => \N__21410\
        );

    \I__3543\ : InMux
    port map (
            O => \N__21433\,
            I => \N__21410\
        );

    \I__3542\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21406\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__21427\,
            I => \N__21399\
        );

    \I__3540\ : Span4Mux_v
    port map (
            O => \N__21424\,
            I => \N__21399\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__21421\,
            I => \N__21399\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__21418\,
            I => \N__21396\
        );

    \I__3537\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21389\
        );

    \I__3536\ : InMux
    port map (
            O => \N__21416\,
            I => \N__21389\
        );

    \I__3535\ : InMux
    port map (
            O => \N__21415\,
            I => \N__21386\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__21410\,
            I => \N__21383\
        );

    \I__3533\ : InMux
    port map (
            O => \N__21409\,
            I => \N__21380\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__21406\,
            I => \N__21373\
        );

    \I__3531\ : Span4Mux_v
    port map (
            O => \N__21399\,
            I => \N__21373\
        );

    \I__3530\ : Span4Mux_s3_v
    port map (
            O => \N__21396\,
            I => \N__21373\
        );

    \I__3529\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21368\
        );

    \I__3528\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21368\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__21389\,
            I => \b2v_inst11.dutycycleZ0Z_10\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__21386\,
            I => \b2v_inst11.dutycycleZ0Z_10\
        );

    \I__3525\ : Odrv4
    port map (
            O => \N__21383\,
            I => \b2v_inst11.dutycycleZ0Z_10\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__21380\,
            I => \b2v_inst11.dutycycleZ0Z_10\
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__21373\,
            I => \b2v_inst11.dutycycleZ0Z_10\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__21368\,
            I => \b2v_inst11.dutycycleZ0Z_10\
        );

    \I__3521\ : InMux
    port map (
            O => \N__21355\,
            I => \N__21349\
        );

    \I__3520\ : InMux
    port map (
            O => \N__21354\,
            I => \N__21349\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__21349\,
            I => \N__21346\
        );

    \I__3518\ : Span4Mux_h
    port map (
            O => \N__21346\,
            I => \N__21343\
        );

    \I__3517\ : Odrv4
    port map (
            O => \N__21343\,
            I => \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQZ0Z5\
        );

    \I__3516\ : InMux
    port map (
            O => \N__21340\,
            I => \b2v_inst11.un1_dutycycle_94_cry_11\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__21337\,
            I => \N__21332\
        );

    \I__3514\ : InMux
    port map (
            O => \N__21336\,
            I => \N__21329\
        );

    \I__3513\ : InMux
    port map (
            O => \N__21335\,
            I => \N__21326\
        );

    \I__3512\ : InMux
    port map (
            O => \N__21332\,
            I => \N__21321\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__21329\,
            I => \N__21318\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__21326\,
            I => \N__21315\
        );

    \I__3509\ : InMux
    port map (
            O => \N__21325\,
            I => \N__21310\
        );

    \I__3508\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21307\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__21321\,
            I => \N__21303\
        );

    \I__3506\ : Span4Mux_h
    port map (
            O => \N__21318\,
            I => \N__21300\
        );

    \I__3505\ : Span4Mux_v
    port map (
            O => \N__21315\,
            I => \N__21297\
        );

    \I__3504\ : InMux
    port map (
            O => \N__21314\,
            I => \N__21294\
        );

    \I__3503\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21291\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__21310\,
            I => \N__21286\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__21307\,
            I => \N__21286\
        );

    \I__3500\ : InMux
    port map (
            O => \N__21306\,
            I => \N__21283\
        );

    \I__3499\ : Span12Mux_s8_h
    port map (
            O => \N__21303\,
            I => \N__21280\
        );

    \I__3498\ : Odrv4
    port map (
            O => \N__21300\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__3497\ : Odrv4
    port map (
            O => \N__21297\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__21294\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__21291\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__3494\ : Odrv4
    port map (
            O => \N__21286\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__21283\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__3492\ : Odrv12
    port map (
            O => \N__21280\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__3491\ : InMux
    port map (
            O => \N__21265\,
            I => \N__21259\
        );

    \I__3490\ : InMux
    port map (
            O => \N__21264\,
            I => \N__21259\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__21259\,
            I => \N__21256\
        );

    \I__3488\ : Span4Mux_h
    port map (
            O => \N__21256\,
            I => \N__21253\
        );

    \I__3487\ : Odrv4
    port map (
            O => \N__21253\,
            I => \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5\
        );

    \I__3486\ : InMux
    port map (
            O => \N__21250\,
            I => \b2v_inst11.un1_dutycycle_94_cry_12\
        );

    \I__3485\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21241\
        );

    \I__3484\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21235\
        );

    \I__3483\ : InMux
    port map (
            O => \N__21245\,
            I => \N__21235\
        );

    \I__3482\ : InMux
    port map (
            O => \N__21244\,
            I => \N__21232\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__21241\,
            I => \N__21228\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__21240\,
            I => \N__21225\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__21235\,
            I => \N__21220\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__21232\,
            I => \N__21217\
        );

    \I__3477\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21214\
        );

    \I__3476\ : Span4Mux_v
    port map (
            O => \N__21228\,
            I => \N__21211\
        );

    \I__3475\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21206\
        );

    \I__3474\ : InMux
    port map (
            O => \N__21224\,
            I => \N__21206\
        );

    \I__3473\ : InMux
    port map (
            O => \N__21223\,
            I => \N__21203\
        );

    \I__3472\ : Span4Mux_h
    port map (
            O => \N__21220\,
            I => \N__21200\
        );

    \I__3471\ : Odrv12
    port map (
            O => \N__21217\,
            I => \b2v_inst11.dutycycleZ0Z_13\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__21214\,
            I => \b2v_inst11.dutycycleZ0Z_13\
        );

    \I__3469\ : Odrv4
    port map (
            O => \N__21211\,
            I => \b2v_inst11.dutycycleZ0Z_13\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__21206\,
            I => \b2v_inst11.dutycycleZ0Z_13\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__21203\,
            I => \b2v_inst11.dutycycleZ0Z_13\
        );

    \I__3466\ : Odrv4
    port map (
            O => \N__21200\,
            I => \b2v_inst11.dutycycleZ0Z_13\
        );

    \I__3465\ : CascadeMux
    port map (
            O => \N__21187\,
            I => \N__21183\
        );

    \I__3464\ : CascadeMux
    port map (
            O => \N__21186\,
            I => \N__21180\
        );

    \I__3463\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21177\
        );

    \I__3462\ : InMux
    port map (
            O => \N__21180\,
            I => \N__21174\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__21177\,
            I => \N__21169\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__21174\,
            I => \N__21169\
        );

    \I__3459\ : Odrv12
    port map (
            O => \N__21169\,
            I => \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5\
        );

    \I__3458\ : InMux
    port map (
            O => \N__21166\,
            I => \b2v_inst11.un1_dutycycle_94_cry_13\
        );

    \I__3457\ : InMux
    port map (
            O => \N__21163\,
            I => \N__21160\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__21160\,
            I => \N__21157\
        );

    \I__3455\ : Span4Mux_s3_v
    port map (
            O => \N__21157\,
            I => \N__21150\
        );

    \I__3454\ : InMux
    port map (
            O => \N__21156\,
            I => \N__21144\
        );

    \I__3453\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21144\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__21154\,
            I => \N__21141\
        );

    \I__3451\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21137\
        );

    \I__3450\ : Span4Mux_v
    port map (
            O => \N__21150\,
            I => \N__21134\
        );

    \I__3449\ : InMux
    port map (
            O => \N__21149\,
            I => \N__21131\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__21144\,
            I => \N__21128\
        );

    \I__3447\ : InMux
    port map (
            O => \N__21141\,
            I => \N__21123\
        );

    \I__3446\ : InMux
    port map (
            O => \N__21140\,
            I => \N__21123\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__21137\,
            I => \N__21120\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__21134\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__21131\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__3442\ : Odrv4
    port map (
            O => \N__21128\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__21123\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__21120\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__3439\ : InMux
    port map (
            O => \N__21109\,
            I => \b2v_inst11.un1_dutycycle_94_cry_14\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__21106\,
            I => \N__21102\
        );

    \I__3437\ : InMux
    port map (
            O => \N__21105\,
            I => \N__21099\
        );

    \I__3436\ : InMux
    port map (
            O => \N__21102\,
            I => \N__21096\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__21099\,
            I => \N__21091\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__21096\,
            I => \N__21091\
        );

    \I__3433\ : Span12Mux_s5_h
    port map (
            O => \N__21091\,
            I => \N__21088\
        );

    \I__3432\ : Odrv12
    port map (
            O => \N__21088\,
            I => \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5\
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__21085\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_5_cascade_\
        );

    \I__3430\ : InMux
    port map (
            O => \N__21082\,
            I => \N__21079\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__21079\,
            I => \b2v_inst11.N_156\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__21076\,
            I => \b2v_inst11.N_156_cascade_\
        );

    \I__3427\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21070\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__21070\,
            I => \b2v_inst11.N_331\
        );

    \I__3425\ : InMux
    port map (
            O => \N__21067\,
            I => \b2v_inst11.un1_dutycycle_94_cry_2\
        );

    \I__3424\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21058\
        );

    \I__3423\ : InMux
    port map (
            O => \N__21063\,
            I => \N__21058\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__21058\,
            I => \N__21055\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__21055\,
            I => \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09\
        );

    \I__3420\ : InMux
    port map (
            O => \N__21052\,
            I => \b2v_inst11.un1_dutycycle_94_cry_3\
        );

    \I__3419\ : InMux
    port map (
            O => \N__21049\,
            I => \b2v_inst11.un1_dutycycle_94_cry_4\
        );

    \I__3418\ : InMux
    port map (
            O => \N__21046\,
            I => \b2v_inst11.un1_dutycycle_94_cry_5_cZ0\
        );

    \I__3417\ : InMux
    port map (
            O => \N__21043\,
            I => \N__21040\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__21040\,
            I => \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39\
        );

    \I__3415\ : InMux
    port map (
            O => \N__21037\,
            I => \b2v_inst11.un1_dutycycle_94_cry_6_cZ0\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__21034\,
            I => \N__21031\
        );

    \I__3413\ : InMux
    port map (
            O => \N__21031\,
            I => \N__21028\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__21028\,
            I => \N__21025\
        );

    \I__3411\ : Span4Mux_h
    port map (
            O => \N__21025\,
            I => \N__21022\
        );

    \I__3410\ : Odrv4
    port map (
            O => \N__21022\,
            I => \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHPZ0Z49\
        );

    \I__3409\ : InMux
    port map (
            O => \N__21019\,
            I => \bfn_6_14_0_\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__21016\,
            I => \N__21008\
        );

    \I__3407\ : InMux
    port map (
            O => \N__21015\,
            I => \N__21005\
        );

    \I__3406\ : InMux
    port map (
            O => \N__21014\,
            I => \N__21002\
        );

    \I__3405\ : InMux
    port map (
            O => \N__21013\,
            I => \N__20999\
        );

    \I__3404\ : InMux
    port map (
            O => \N__21012\,
            I => \N__20989\
        );

    \I__3403\ : InMux
    port map (
            O => \N__21011\,
            I => \N__20989\
        );

    \I__3402\ : InMux
    port map (
            O => \N__21008\,
            I => \N__20986\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__21005\,
            I => \N__20983\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__21002\,
            I => \N__20980\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__20999\,
            I => \N__20977\
        );

    \I__3398\ : InMux
    port map (
            O => \N__20998\,
            I => \N__20971\
        );

    \I__3397\ : InMux
    port map (
            O => \N__20997\,
            I => \N__20971\
        );

    \I__3396\ : InMux
    port map (
            O => \N__20996\,
            I => \N__20968\
        );

    \I__3395\ : InMux
    port map (
            O => \N__20995\,
            I => \N__20963\
        );

    \I__3394\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20963\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__20989\,
            I => \N__20960\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__20986\,
            I => \N__20949\
        );

    \I__3391\ : Span4Mux_v
    port map (
            O => \N__20983\,
            I => \N__20949\
        );

    \I__3390\ : Span4Mux_h
    port map (
            O => \N__20980\,
            I => \N__20949\
        );

    \I__3389\ : Span4Mux_h
    port map (
            O => \N__20977\,
            I => \N__20946\
        );

    \I__3388\ : InMux
    port map (
            O => \N__20976\,
            I => \N__20943\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__20971\,
            I => \N__20934\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__20968\,
            I => \N__20934\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__20963\,
            I => \N__20934\
        );

    \I__3384\ : Span4Mux_h
    port map (
            O => \N__20960\,
            I => \N__20934\
        );

    \I__3383\ : InMux
    port map (
            O => \N__20959\,
            I => \N__20925\
        );

    \I__3382\ : InMux
    port map (
            O => \N__20958\,
            I => \N__20925\
        );

    \I__3381\ : InMux
    port map (
            O => \N__20957\,
            I => \N__20925\
        );

    \I__3380\ : InMux
    port map (
            O => \N__20956\,
            I => \N__20925\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__20949\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__3378\ : Odrv4
    port map (
            O => \N__20946\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__20943\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__3376\ : Odrv4
    port map (
            O => \N__20934\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__20925\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__20914\,
            I => \N__20911\
        );

    \I__3373\ : InMux
    port map (
            O => \N__20911\,
            I => \N__20905\
        );

    \I__3372\ : InMux
    port map (
            O => \N__20910\,
            I => \N__20905\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__20905\,
            I => \N__20902\
        );

    \I__3370\ : Odrv4
    port map (
            O => \N__20902\,
            I => \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59\
        );

    \I__3369\ : InMux
    port map (
            O => \N__20899\,
            I => \b2v_inst11.un1_dutycycle_94_cry_8_cZ0\
        );

    \I__3368\ : InMux
    port map (
            O => \N__20896\,
            I => \b2v_inst11.un1_dutycycle_94_cry_9_cZ0\
        );

    \I__3367\ : CascadeMux
    port map (
            O => \N__20893\,
            I => \N__20887\
        );

    \I__3366\ : InMux
    port map (
            O => \N__20892\,
            I => \N__20884\
        );

    \I__3365\ : InMux
    port map (
            O => \N__20891\,
            I => \N__20881\
        );

    \I__3364\ : InMux
    port map (
            O => \N__20890\,
            I => \N__20877\
        );

    \I__3363\ : InMux
    port map (
            O => \N__20887\,
            I => \N__20871\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__20884\,
            I => \N__20866\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__20881\,
            I => \N__20866\
        );

    \I__3360\ : InMux
    port map (
            O => \N__20880\,
            I => \N__20863\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__20877\,
            I => \N__20860\
        );

    \I__3358\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20853\
        );

    \I__3357\ : InMux
    port map (
            O => \N__20875\,
            I => \N__20853\
        );

    \I__3356\ : InMux
    port map (
            O => \N__20874\,
            I => \N__20853\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__20871\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__3354\ : Odrv12
    port map (
            O => \N__20866\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__20863\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__3352\ : Odrv4
    port map (
            O => \N__20860\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__20853\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__20842\,
            I => \b2v_inst11.dutycycle_RNI74A23Z0Z_7_cascade_\
        );

    \I__3349\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20836\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__20836\,
            I => \b2v_inst11.dutycycle_e_1_7\
        );

    \I__3347\ : InMux
    port map (
            O => \N__20833\,
            I => \N__20830\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__20830\,
            I => \b2v_inst11.dutycycle_RNI74A23Z0Z_7\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__20827\,
            I => \b2v_inst11.dutycycle_e_1_7_cascade_\
        );

    \I__3344\ : InMux
    port map (
            O => \N__20824\,
            I => \N__20821\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__20821\,
            I => \N__20818\
        );

    \I__3342\ : Span4Mux_h
    port map (
            O => \N__20818\,
            I => \N__20815\
        );

    \I__3341\ : Odrv4
    port map (
            O => \N__20815\,
            I => \b2v_inst11.dutycycle_RNI01TT1Z0Z_7\
        );

    \I__3340\ : CascadeMux
    port map (
            O => \N__20812\,
            I => \b2v_inst11.dutycycle_RNI25OT3Z0Z_7_cascade_\
        );

    \I__3339\ : CascadeMux
    port map (
            O => \N__20809\,
            I => \N__20806\
        );

    \I__3338\ : InMux
    port map (
            O => \N__20806\,
            I => \N__20803\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__20803\,
            I => \b2v_inst11.func_state_RNIGALV4Z0Z_0\
        );

    \I__3336\ : InMux
    port map (
            O => \N__20800\,
            I => \N__20788\
        );

    \I__3335\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20788\
        );

    \I__3334\ : InMux
    port map (
            O => \N__20798\,
            I => \N__20788\
        );

    \I__3333\ : InMux
    port map (
            O => \N__20797\,
            I => \N__20788\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__20788\,
            I => \b2v_inst11.dutycycleZ1Z_7\
        );

    \I__3331\ : InMux
    port map (
            O => \N__20785\,
            I => \N__20782\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__20782\,
            I => \b2v_inst11.dutycycle_RNIGSFQZ0Z_7\
        );

    \I__3329\ : InMux
    port map (
            O => \N__20779\,
            I => \b2v_inst11.un1_dutycycle_94_cry_0_cZ0\
        );

    \I__3328\ : InMux
    port map (
            O => \N__20776\,
            I => \N__20773\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__20773\,
            I => \N__20770\
        );

    \I__3326\ : Span4Mux_h
    port map (
            O => \N__20770\,
            I => \N__20767\
        );

    \I__3325\ : Odrv4
    port map (
            O => \N__20767\,
            I => \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDUZ0Z8\
        );

    \I__3324\ : InMux
    port map (
            O => \N__20764\,
            I => \b2v_inst11.un1_dutycycle_94_cry_1\
        );

    \I__3323\ : CascadeMux
    port map (
            O => \N__20761\,
            I => \b2v_inst11.dutycycleZ0Z_8_cascade_\
        );

    \I__3322\ : CascadeMux
    port map (
            O => \N__20758\,
            I => \b2v_inst11.dutycycle_RNIAI7C4Z0Z_4_cascade_\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__20755\,
            I => \N__20752\
        );

    \I__3320\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20749\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__20749\,
            I => \b2v_inst11.dutycycle_eena_2_0_1\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__20746\,
            I => \b2v_inst11.func_state_RNI3JFN6Z0Z_0_cascade_\
        );

    \I__3317\ : InMux
    port map (
            O => \N__20743\,
            I => \N__20737\
        );

    \I__3316\ : InMux
    port map (
            O => \N__20742\,
            I => \N__20737\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__20737\,
            I => \b2v_inst11.dutycycle_RNI3JFN6Z0Z_4\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__20734\,
            I => \N__20730\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__20733\,
            I => \N__20727\
        );

    \I__3312\ : InMux
    port map (
            O => \N__20730\,
            I => \N__20722\
        );

    \I__3311\ : InMux
    port map (
            O => \N__20727\,
            I => \N__20722\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__20722\,
            I => \b2v_inst11.dutycycleZ1Z_4\
        );

    \I__3309\ : InMux
    port map (
            O => \N__20719\,
            I => \N__20713\
        );

    \I__3308\ : InMux
    port map (
            O => \N__20718\,
            I => \N__20713\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__20713\,
            I => \b2v_inst11.dutycycleZ1Z_9\
        );

    \I__3306\ : InMux
    port map (
            O => \N__20710\,
            I => \N__20707\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__20707\,
            I => \b2v_inst11.func_state_RNI3JFN6Z0Z_0\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__20704\,
            I => \b2v_inst11.dutycycle_RNI0KJ31Z0Z_7_cascade_\
        );

    \I__3303\ : InMux
    port map (
            O => \N__20701\,
            I => \N__20695\
        );

    \I__3302\ : InMux
    port map (
            O => \N__20700\,
            I => \N__20695\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__20695\,
            I => \b2v_inst11.dutycycleZ0Z_14\
        );

    \I__3300\ : InMux
    port map (
            O => \N__20692\,
            I => \N__20688\
        );

    \I__3299\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20685\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__20688\,
            I => \N__20680\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__20685\,
            I => \N__20680\
        );

    \I__3296\ : Odrv4
    port map (
            O => \N__20680\,
            I => \b2v_inst11.dutycycle_en_11\
        );

    \I__3295\ : CascadeMux
    port map (
            O => \N__20677\,
            I => \b2v_inst11.dutycycleZ0Z_13_cascade_\
        );

    \I__3294\ : InMux
    port map (
            O => \N__20674\,
            I => \N__20671\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__20671\,
            I => \b2v_inst11.un2_count_clk_17_0_a2_1_4\
        );

    \I__3292\ : InMux
    port map (
            O => \N__20668\,
            I => \N__20665\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__20665\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_4\
        );

    \I__3290\ : CascadeMux
    port map (
            O => \N__20662\,
            I => \b2v_inst11.un1_dutycycle_53_50_a4_0_cascade_\
        );

    \I__3289\ : InMux
    port map (
            O => \N__20659\,
            I => \N__20655\
        );

    \I__3288\ : InMux
    port map (
            O => \N__20658\,
            I => \N__20652\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__20655\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_10\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__20652\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_10\
        );

    \I__3285\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20644\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__20644\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_7\
        );

    \I__3283\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20638\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__20638\,
            I => \N__20635\
        );

    \I__3281\ : Sp12to4
    port map (
            O => \N__20635\,
            I => \N__20632\
        );

    \I__3280\ : Odrv12
    port map (
            O => \N__20632\,
            I => \VCCST_OK_c\
        );

    \I__3279\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20619\
        );

    \I__3278\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20619\
        );

    \I__3277\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20619\
        );

    \I__3276\ : InMux
    port map (
            O => \N__20626\,
            I => \N__20616\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__20619\,
            I => \N__20613\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__20616\,
            I => \N__20610\
        );

    \I__3273\ : Odrv12
    port map (
            O => \N__20613\,
            I => \VDDQ_OK_c\
        );

    \I__3272\ : Odrv12
    port map (
            O => \N__20610\,
            I => \VDDQ_OK_c\
        );

    \I__3271\ : IoInMux
    port map (
            O => \N__20605\,
            I => \N__20602\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__20602\,
            I => \N__20599\
        );

    \I__3269\ : Odrv12
    port map (
            O => \N__20599\,
            I => \VCCIO_EN_c\
        );

    \I__3268\ : InMux
    port map (
            O => \N__20596\,
            I => \N__20593\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__20593\,
            I => \N__20589\
        );

    \I__3266\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20586\
        );

    \I__3265\ : Odrv4
    port map (
            O => \N__20589\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_3\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__20586\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_3\
        );

    \I__3263\ : CascadeMux
    port map (
            O => \N__20581\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_3_cascade_\
        );

    \I__3262\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20575\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__20575\,
            I => \b2v_inst11.un1_dutycycle_53_axb_7_1\
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__20572\,
            I => \N__20569\
        );

    \I__3259\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20566\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__20566\,
            I => \N__20563\
        );

    \I__3257\ : Odrv4
    port map (
            O => \N__20563\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_9\
        );

    \I__3256\ : InMux
    port map (
            O => \N__20560\,
            I => \N__20557\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__20557\,
            I => \b2v_inst16.curr_state_1_0\
        );

    \I__3254\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20551\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__20551\,
            I => \b2v_inst16.curr_stateZ0Z_0\
        );

    \I__3252\ : CascadeMux
    port map (
            O => \N__20548\,
            I => \N__20545\
        );

    \I__3251\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20537\
        );

    \I__3250\ : InMux
    port map (
            O => \N__20544\,
            I => \N__20526\
        );

    \I__3249\ : InMux
    port map (
            O => \N__20543\,
            I => \N__20526\
        );

    \I__3248\ : InMux
    port map (
            O => \N__20542\,
            I => \N__20526\
        );

    \I__3247\ : InMux
    port map (
            O => \N__20541\,
            I => \N__20526\
        );

    \I__3246\ : InMux
    port map (
            O => \N__20540\,
            I => \N__20526\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__20537\,
            I => \b2v_inst16.curr_stateZ0Z_1\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__20526\,
            I => \b2v_inst16.curr_stateZ0Z_1\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__20521\,
            I => \N__20518\
        );

    \I__3242\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20515\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__20515\,
            I => \N__20512\
        );

    \I__3240\ : Odrv4
    port map (
            O => \N__20512\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_0\
        );

    \I__3239\ : InMux
    port map (
            O => \N__20509\,
            I => \N__20506\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__20506\,
            I => \N__20503\
        );

    \I__3237\ : Span4Mux_h
    port map (
            O => \N__20503\,
            I => \N__20500\
        );

    \I__3236\ : Span4Mux_h
    port map (
            O => \N__20500\,
            I => \N__20497\
        );

    \I__3235\ : Odrv4
    port map (
            O => \N__20497\,
            I => \b2v_inst200.count_RNIC03N_3Z0Z_0\
        );

    \I__3234\ : IoInMux
    port map (
            O => \N__20494\,
            I => \N__20490\
        );

    \I__3233\ : IoInMux
    port map (
            O => \N__20493\,
            I => \N__20487\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__20490\,
            I => \N__20484\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__20487\,
            I => \N__20481\
        );

    \I__3230\ : Span4Mux_s1_h
    port map (
            O => \N__20484\,
            I => \N__20478\
        );

    \I__3229\ : IoSpan4Mux
    port map (
            O => \N__20481\,
            I => \N__20475\
        );

    \I__3228\ : Span4Mux_v
    port map (
            O => \N__20478\,
            I => \N__20470\
        );

    \I__3227\ : Span4Mux_s1_h
    port map (
            O => \N__20475\,
            I => \N__20470\
        );

    \I__3226\ : Span4Mux_h
    port map (
            O => \N__20470\,
            I => \N__20467\
        );

    \I__3225\ : Odrv4
    port map (
            O => \N__20467\,
            I => \V105A_EN_c\
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__20464\,
            I => \N__20461\
        );

    \I__3223\ : InMux
    port map (
            O => \N__20461\,
            I => \N__20458\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__20458\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_5\
        );

    \I__3221\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20452\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__20452\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_10\
        );

    \I__3219\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20446\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__20446\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_5\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__20443\,
            I => \N__20439\
        );

    \I__3216\ : InMux
    port map (
            O => \N__20442\,
            I => \N__20436\
        );

    \I__3215\ : InMux
    port map (
            O => \N__20439\,
            I => \N__20433\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__20436\,
            I => \N__20430\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__20433\,
            I => \N__20427\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__20430\,
            I => \b2v_inst11.mult1_un54_sum\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__20427\,
            I => \b2v_inst11.mult1_un54_sum\
        );

    \I__3210\ : InMux
    port map (
            O => \N__20422\,
            I => \N__20419\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__20419\,
            I => \b2v_inst11.mult1_un54_sum_i\
        );

    \I__3208\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20412\
        );

    \I__3207\ : InMux
    port map (
            O => \N__20415\,
            I => \N__20409\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__20412\,
            I => \N__20406\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__20409\,
            I => \N__20403\
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__20406\,
            I => \b2v_inst11.mult1_un61_sum\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__20403\,
            I => \b2v_inst11.mult1_un61_sum\
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__20398\,
            I => \N__20395\
        );

    \I__3201\ : InMux
    port map (
            O => \N__20395\,
            I => \N__20392\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__20392\,
            I => \b2v_inst11.mult1_un61_sum_i\
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__20389\,
            I => \N__20385\
        );

    \I__3198\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20380\
        );

    \I__3197\ : InMux
    port map (
            O => \N__20385\,
            I => \N__20375\
        );

    \I__3196\ : InMux
    port map (
            O => \N__20384\,
            I => \N__20375\
        );

    \I__3195\ : InMux
    port map (
            O => \N__20383\,
            I => \N__20372\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__20380\,
            I => \b2v_inst11.mult1_un68_sum_s_8\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__20375\,
            I => \b2v_inst11.mult1_un68_sum_s_8\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__20372\,
            I => \b2v_inst11.mult1_un68_sum_s_8\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__20365\,
            I => \b2v_inst16.curr_stateZ0Z_1_cascade_\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__20362\,
            I => \b2v_inst16.curr_state_7_0_cascade_\
        );

    \I__3189\ : InMux
    port map (
            O => \N__20359\,
            I => \N__20353\
        );

    \I__3188\ : InMux
    port map (
            O => \N__20358\,
            I => \N__20353\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__20353\,
            I => \N__20350\
        );

    \I__3186\ : Span4Mux_h
    port map (
            O => \N__20350\,
            I => \N__20347\
        );

    \I__3185\ : Span4Mux_v
    port map (
            O => \N__20347\,
            I => \N__20336\
        );

    \I__3184\ : InMux
    port map (
            O => \N__20346\,
            I => \N__20331\
        );

    \I__3183\ : InMux
    port map (
            O => \N__20345\,
            I => \N__20331\
        );

    \I__3182\ : InMux
    port map (
            O => \N__20344\,
            I => \N__20326\
        );

    \I__3181\ : InMux
    port map (
            O => \N__20343\,
            I => \N__20326\
        );

    \I__3180\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20319\
        );

    \I__3179\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20319\
        );

    \I__3178\ : InMux
    port map (
            O => \N__20340\,
            I => \N__20319\
        );

    \I__3177\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20316\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__20336\,
            I => \b2v_inst16.un13_clk_100khz_i\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__20331\,
            I => \b2v_inst16.un13_clk_100khz_i\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__20326\,
            I => \b2v_inst16.un13_clk_100khz_i\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__20319\,
            I => \b2v_inst16.un13_clk_100khz_i\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__20316\,
            I => \b2v_inst16.un13_clk_100khz_i\
        );

    \I__3171\ : CascadeMux
    port map (
            O => \N__20305\,
            I => \N__20302\
        );

    \I__3170\ : InMux
    port map (
            O => \N__20302\,
            I => \N__20299\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__20299\,
            I => \b2v_inst16.curr_state_0_1\
        );

    \I__3168\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20293\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__20293\,
            I => \b2v_inst16.delayed_vddq_pwrgdZ0\
        );

    \I__3166\ : IoInMux
    port map (
            O => \N__20290\,
            I => \N__20287\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__20287\,
            I => \N__20284\
        );

    \I__3164\ : Span4Mux_s2_h
    port map (
            O => \N__20284\,
            I => \N__20281\
        );

    \I__3163\ : Span4Mux_h
    port map (
            O => \N__20281\,
            I => \N__20278\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__20278\,
            I => b2v_inst16_un2_vpp_en_0_i
        );

    \I__3161\ : InMux
    port map (
            O => \N__20275\,
            I => \N__20268\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__20274\,
            I => \N__20265\
        );

    \I__3159\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20256\
        );

    \I__3158\ : InMux
    port map (
            O => \N__20272\,
            I => \N__20256\
        );

    \I__3157\ : InMux
    port map (
            O => \N__20271\,
            I => \N__20256\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__20268\,
            I => \N__20253\
        );

    \I__3155\ : InMux
    port map (
            O => \N__20265\,
            I => \N__20248\
        );

    \I__3154\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20248\
        );

    \I__3153\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20245\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__20256\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__3151\ : Odrv4
    port map (
            O => \N__20253\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__20248\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__20245\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__3148\ : InMux
    port map (
            O => \N__20236\,
            I => \N__20233\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__20233\,
            I => \N__20229\
        );

    \I__3146\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20226\
        );

    \I__3145\ : Span4Mux_s2_v
    port map (
            O => \N__20229\,
            I => \N__20221\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__20226\,
            I => \N__20221\
        );

    \I__3143\ : Odrv4
    port map (
            O => \N__20221\,
            I => \b2v_inst11.mult1_un124_sum\
        );

    \I__3142\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20215\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__20215\,
            I => \b2v_inst11.mult1_un124_sum_i\
        );

    \I__3140\ : InMux
    port map (
            O => \N__20212\,
            I => \N__20209\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__20209\,
            I => \N__20205\
        );

    \I__3138\ : InMux
    port map (
            O => \N__20208\,
            I => \N__20202\
        );

    \I__3137\ : Span4Mux_h
    port map (
            O => \N__20205\,
            I => \N__20197\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__20202\,
            I => \N__20197\
        );

    \I__3135\ : Span4Mux_v
    port map (
            O => \N__20197\,
            I => \N__20194\
        );

    \I__3134\ : Odrv4
    port map (
            O => \N__20194\,
            I => \b2v_inst11.mult1_un89_sum\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__20191\,
            I => \N__20188\
        );

    \I__3132\ : InMux
    port map (
            O => \N__20188\,
            I => \N__20185\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__20185\,
            I => \N__20182\
        );

    \I__3130\ : Span4Mux_s3_v
    port map (
            O => \N__20182\,
            I => \N__20179\
        );

    \I__3129\ : Odrv4
    port map (
            O => \N__20179\,
            I => \b2v_inst11.mult1_un89_sum_i\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__20176\,
            I => \N__20172\
        );

    \I__3127\ : InMux
    port map (
            O => \N__20175\,
            I => \N__20164\
        );

    \I__3126\ : InMux
    port map (
            O => \N__20172\,
            I => \N__20164\
        );

    \I__3125\ : InMux
    port map (
            O => \N__20171\,
            I => \N__20164\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__20164\,
            I => \b2v_inst11.mult1_un61_sum_i_0_8\
        );

    \I__3123\ : InMux
    port map (
            O => \N__20161\,
            I => \N__20158\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__20158\,
            I => \N__20154\
        );

    \I__3121\ : CascadeMux
    port map (
            O => \N__20157\,
            I => \N__20150\
        );

    \I__3120\ : Span4Mux_v
    port map (
            O => \N__20154\,
            I => \N__20145\
        );

    \I__3119\ : InMux
    port map (
            O => \N__20153\,
            I => \N__20142\
        );

    \I__3118\ : InMux
    port map (
            O => \N__20150\,
            I => \N__20137\
        );

    \I__3117\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20137\
        );

    \I__3116\ : InMux
    port map (
            O => \N__20148\,
            I => \N__20134\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__20145\,
            I => \b2v_inst11.mult1_un110_sum_s_8\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__20142\,
            I => \b2v_inst11.mult1_un110_sum_s_8\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__20137\,
            I => \b2v_inst11.mult1_un110_sum_s_8\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__20134\,
            I => \b2v_inst11.mult1_un110_sum_s_8\
        );

    \I__3111\ : IoInMux
    port map (
            O => \N__20125\,
            I => \N__20122\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__20122\,
            I => \N__20119\
        );

    \I__3109\ : IoSpan4Mux
    port map (
            O => \N__20119\,
            I => \N__20115\
        );

    \I__3108\ : InMux
    port map (
            O => \N__20118\,
            I => \N__20111\
        );

    \I__3107\ : Span4Mux_s1_h
    port map (
            O => \N__20115\,
            I => \N__20108\
        );

    \I__3106\ : InMux
    port map (
            O => \N__20114\,
            I => \N__20105\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__20111\,
            I => \N__20102\
        );

    \I__3104\ : Span4Mux_h
    port map (
            O => \N__20108\,
            I => \N__20097\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__20105\,
            I => \N__20097\
        );

    \I__3102\ : Span4Mux_v
    port map (
            O => \N__20102\,
            I => \N__20093\
        );

    \I__3101\ : Span4Mux_v
    port map (
            O => \N__20097\,
            I => \N__20090\
        );

    \I__3100\ : InMux
    port map (
            O => \N__20096\,
            I => \N__20087\
        );

    \I__3099\ : Odrv4
    port map (
            O => \N__20093\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__20090\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__20087\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3096\ : InMux
    port map (
            O => \N__20080\,
            I => \N__20077\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__20077\,
            I => \N__20073\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__20076\,
            I => \N__20070\
        );

    \I__3093\ : Span4Mux_v
    port map (
            O => \N__20073\,
            I => \N__20065\
        );

    \I__3092\ : InMux
    port map (
            O => \N__20070\,
            I => \N__20060\
        );

    \I__3091\ : InMux
    port map (
            O => \N__20069\,
            I => \N__20060\
        );

    \I__3090\ : InMux
    port map (
            O => \N__20068\,
            I => \N__20057\
        );

    \I__3089\ : Odrv4
    port map (
            O => \N__20065\,
            I => \b2v_inst11.mult1_un75_sum_s_8\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__20060\,
            I => \b2v_inst11.mult1_un75_sum_s_8\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__20057\,
            I => \b2v_inst11.mult1_un75_sum_s_8\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__20050\,
            I => \N__20046\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__20049\,
            I => \N__20042\
        );

    \I__3084\ : InMux
    port map (
            O => \N__20046\,
            I => \N__20039\
        );

    \I__3083\ : InMux
    port map (
            O => \N__20045\,
            I => \N__20034\
        );

    \I__3082\ : InMux
    port map (
            O => \N__20042\,
            I => \N__20031\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__20039\,
            I => \N__20028\
        );

    \I__3080\ : InMux
    port map (
            O => \N__20038\,
            I => \N__20025\
        );

    \I__3079\ : InMux
    port map (
            O => \N__20037\,
            I => \N__20022\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__20034\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__20031\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__3076\ : Odrv4
    port map (
            O => \N__20028\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__20025\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__20022\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__3073\ : InMux
    port map (
            O => \N__20011\,
            I => \N__20008\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__20008\,
            I => \N__20004\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__20007\,
            I => \N__20001\
        );

    \I__3070\ : Span4Mux_v
    port map (
            O => \N__20004\,
            I => \N__19996\
        );

    \I__3069\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19991\
        );

    \I__3068\ : InMux
    port map (
            O => \N__20000\,
            I => \N__19991\
        );

    \I__3067\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19988\
        );

    \I__3066\ : Odrv4
    port map (
            O => \N__19996\,
            I => \b2v_inst11.mult1_un96_sum_s_8\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__19991\,
            I => \b2v_inst11.mult1_un96_sum_s_8\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__19988\,
            I => \b2v_inst11.mult1_un96_sum_s_8\
        );

    \I__3063\ : InMux
    port map (
            O => \N__19981\,
            I => \b2v_inst11.mult1_un131_sum_cry_3\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__19978\,
            I => \N__19975\
        );

    \I__3061\ : InMux
    port map (
            O => \N__19975\,
            I => \N__19972\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__19972\,
            I => \N__19969\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__19969\,
            I => \b2v_inst11.mult1_un124_sum_cry_4_s\
        );

    \I__3058\ : InMux
    port map (
            O => \N__19966\,
            I => \b2v_inst11.mult1_un131_sum_cry_4\
        );

    \I__3057\ : InMux
    port map (
            O => \N__19963\,
            I => \N__19960\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__19960\,
            I => \b2v_inst11.mult1_un124_sum_cry_5_s\
        );

    \I__3055\ : InMux
    port map (
            O => \N__19957\,
            I => \b2v_inst11.mult1_un131_sum_cry_5\
        );

    \I__3054\ : InMux
    port map (
            O => \N__19954\,
            I => \N__19951\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__19951\,
            I => \b2v_inst11.mult1_un131_sum_axb_7_l_fx\
        );

    \I__3052\ : CascadeMux
    port map (
            O => \N__19948\,
            I => \N__19945\
        );

    \I__3051\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19941\
        );

    \I__3050\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19938\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__19941\,
            I => \N__19935\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__19938\,
            I => \b2v_inst11.mult1_un124_sum_cry_6_s\
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__19935\,
            I => \b2v_inst11.mult1_un124_sum_cry_6_s\
        );

    \I__3046\ : InMux
    port map (
            O => \N__19930\,
            I => \b2v_inst11.mult1_un131_sum_cry_6\
        );

    \I__3045\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19924\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__19924\,
            I => \b2v_inst11.mult1_un131_sum_axb_8\
        );

    \I__3043\ : InMux
    port map (
            O => \N__19921\,
            I => \b2v_inst11.mult1_un131_sum_cry_7\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__19918\,
            I => \b2v_inst11.mult1_un131_sum_s_8_cascade_\
        );

    \I__3041\ : InMux
    port map (
            O => \N__19915\,
            I => \N__19911\
        );

    \I__3040\ : InMux
    port map (
            O => \N__19914\,
            I => \N__19908\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__19911\,
            I => \N__19903\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__19908\,
            I => \N__19903\
        );

    \I__3037\ : Span4Mux_v
    port map (
            O => \N__19903\,
            I => \N__19900\
        );

    \I__3036\ : Odrv4
    port map (
            O => \N__19900\,
            I => \b2v_inst11.mult1_un68_sum\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__19897\,
            I => \N__19894\
        );

    \I__3034\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19891\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__19891\,
            I => \N__19888\
        );

    \I__3032\ : Odrv4
    port map (
            O => \N__19888\,
            I => \b2v_inst11.mult1_un68_sum_i\
        );

    \I__3031\ : InMux
    port map (
            O => \N__19885\,
            I => \N__19881\
        );

    \I__3030\ : CascadeMux
    port map (
            O => \N__19884\,
            I => \N__19878\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__19881\,
            I => \N__19873\
        );

    \I__3028\ : InMux
    port map (
            O => \N__19878\,
            I => \N__19868\
        );

    \I__3027\ : InMux
    port map (
            O => \N__19877\,
            I => \N__19868\
        );

    \I__3026\ : InMux
    port map (
            O => \N__19876\,
            I => \N__19865\
        );

    \I__3025\ : Odrv12
    port map (
            O => \N__19873\,
            I => \b2v_inst11.mult1_un117_sum_s_8\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__19868\,
            I => \b2v_inst11.mult1_un117_sum_s_8\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__19865\,
            I => \b2v_inst11.mult1_un117_sum_s_8\
        );

    \I__3022\ : InMux
    port map (
            O => \N__19858\,
            I => \N__19855\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__19855\,
            I => \N__19851\
        );

    \I__3020\ : InMux
    port map (
            O => \N__19854\,
            I => \N__19848\
        );

    \I__3019\ : Span4Mux_s2_v
    port map (
            O => \N__19851\,
            I => \N__19843\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__19848\,
            I => \N__19843\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__19843\,
            I => \b2v_inst11.mult1_un117_sum\
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__19840\,
            I => \N__19837\
        );

    \I__3015\ : InMux
    port map (
            O => \N__19837\,
            I => \N__19834\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__19834\,
            I => \N__19831\
        );

    \I__3013\ : Odrv4
    port map (
            O => \N__19831\,
            I => \b2v_inst11.mult1_un117_sum_i\
        );

    \I__3012\ : InMux
    port map (
            O => \N__19828\,
            I => \N__19825\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__19825\,
            I => \b2v_inst11.mult1_un117_sum_cry_3_s\
        );

    \I__3010\ : InMux
    port map (
            O => \N__19822\,
            I => \b2v_inst11.mult1_un124_sum_cry_3\
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__19819\,
            I => \N__19816\
        );

    \I__3008\ : InMux
    port map (
            O => \N__19816\,
            I => \N__19813\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__19813\,
            I => \b2v_inst11.mult1_un117_sum_cry_4_s\
        );

    \I__3006\ : InMux
    port map (
            O => \N__19810\,
            I => \b2v_inst11.mult1_un124_sum_cry_4\
        );

    \I__3005\ : InMux
    port map (
            O => \N__19807\,
            I => \N__19804\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__19804\,
            I => \b2v_inst11.mult1_un117_sum_cry_5_s\
        );

    \I__3003\ : InMux
    port map (
            O => \N__19801\,
            I => \b2v_inst11.mult1_un124_sum_cry_5\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__19798\,
            I => \N__19794\
        );

    \I__3001\ : InMux
    port map (
            O => \N__19797\,
            I => \N__19786\
        );

    \I__3000\ : InMux
    port map (
            O => \N__19794\,
            I => \N__19786\
        );

    \I__2999\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19786\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__19786\,
            I => \b2v_inst11.mult1_un117_sum_i_0_8\
        );

    \I__2997\ : CascadeMux
    port map (
            O => \N__19783\,
            I => \N__19780\
        );

    \I__2996\ : InMux
    port map (
            O => \N__19780\,
            I => \N__19777\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__19777\,
            I => \b2v_inst11.mult1_un117_sum_cry_6_s\
        );

    \I__2994\ : InMux
    port map (
            O => \N__19774\,
            I => \b2v_inst11.mult1_un124_sum_cry_6\
        );

    \I__2993\ : InMux
    port map (
            O => \N__19771\,
            I => \N__19768\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__19768\,
            I => \b2v_inst11.mult1_un124_sum_axb_8\
        );

    \I__2991\ : InMux
    port map (
            O => \N__19765\,
            I => \b2v_inst11.mult1_un124_sum_cry_7\
        );

    \I__2990\ : CascadeMux
    port map (
            O => \N__19762\,
            I => \N__19758\
        );

    \I__2989\ : InMux
    port map (
            O => \N__19761\,
            I => \N__19750\
        );

    \I__2988\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19750\
        );

    \I__2987\ : InMux
    port map (
            O => \N__19757\,
            I => \N__19750\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__19750\,
            I => \b2v_inst11.mult1_un110_sum_i_0_8\
        );

    \I__2985\ : CascadeMux
    port map (
            O => \N__19747\,
            I => \N__19744\
        );

    \I__2984\ : InMux
    port map (
            O => \N__19744\,
            I => \N__19741\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__19741\,
            I => \b2v_inst11.mult1_un124_sum_i_0_8\
        );

    \I__2982\ : InMux
    port map (
            O => \N__19738\,
            I => \b2v_inst11.mult1_un131_sum_cry_2\
        );

    \I__2981\ : InMux
    port map (
            O => \N__19735\,
            I => \N__19732\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__19732\,
            I => \b2v_inst11.mult1_un131_sum_axb_4_l_fx\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__19729\,
            I => \N__19725\
        );

    \I__2978\ : InMux
    port map (
            O => \N__19728\,
            I => \N__19722\
        );

    \I__2977\ : InMux
    port map (
            O => \N__19725\,
            I => \N__19719\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__19722\,
            I => \b2v_inst11.mult1_un124_sum_cry_3_s\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__19719\,
            I => \b2v_inst11.mult1_un124_sum_cry_3_s\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__19714\,
            I => \N__19711\
        );

    \I__2973\ : InMux
    port map (
            O => \N__19711\,
            I => \N__19708\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__19708\,
            I => \N__19705\
        );

    \I__2971\ : Odrv4
    port map (
            O => \N__19705\,
            I => \b2v_inst11.mult1_un110_sum_i\
        );

    \I__2970\ : InMux
    port map (
            O => \N__19702\,
            I => \b2v_inst11.mult1_un117_sum_cry_2\
        );

    \I__2969\ : InMux
    port map (
            O => \N__19699\,
            I => \N__19696\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__19696\,
            I => \b2v_inst11.mult1_un110_sum_cry_3_s\
        );

    \I__2967\ : InMux
    port map (
            O => \N__19693\,
            I => \b2v_inst11.mult1_un117_sum_cry_3\
        );

    \I__2966\ : CascadeMux
    port map (
            O => \N__19690\,
            I => \N__19687\
        );

    \I__2965\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19684\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__19684\,
            I => \b2v_inst11.mult1_un110_sum_cry_4_s\
        );

    \I__2963\ : InMux
    port map (
            O => \N__19681\,
            I => \b2v_inst11.mult1_un117_sum_cry_4\
        );

    \I__2962\ : InMux
    port map (
            O => \N__19678\,
            I => \N__19675\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__19675\,
            I => \b2v_inst11.mult1_un110_sum_cry_5_s\
        );

    \I__2960\ : InMux
    port map (
            O => \N__19672\,
            I => \b2v_inst11.mult1_un117_sum_cry_5\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__19669\,
            I => \N__19666\
        );

    \I__2958\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19663\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__19663\,
            I => \b2v_inst11.mult1_un110_sum_cry_6_s\
        );

    \I__2956\ : InMux
    port map (
            O => \N__19660\,
            I => \b2v_inst11.mult1_un117_sum_cry_6\
        );

    \I__2955\ : InMux
    port map (
            O => \N__19657\,
            I => \N__19654\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__19654\,
            I => \b2v_inst11.mult1_un117_sum_axb_8\
        );

    \I__2953\ : InMux
    port map (
            O => \N__19651\,
            I => \b2v_inst11.mult1_un117_sum_cry_7\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__19648\,
            I => \b2v_inst11.mult1_un117_sum_s_8_cascade_\
        );

    \I__2951\ : InMux
    port map (
            O => \N__19645\,
            I => \b2v_inst11.mult1_un124_sum_cry_2\
        );

    \I__2950\ : InMux
    port map (
            O => \N__19642\,
            I => \N__19638\
        );

    \I__2949\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19634\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__19638\,
            I => \N__19631\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__19637\,
            I => \N__19628\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__19634\,
            I => \N__19625\
        );

    \I__2945\ : Span4Mux_h
    port map (
            O => \N__19631\,
            I => \N__19622\
        );

    \I__2944\ : InMux
    port map (
            O => \N__19628\,
            I => \N__19619\
        );

    \I__2943\ : Span4Mux_h
    port map (
            O => \N__19625\,
            I => \N__19616\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__19622\,
            I => \b2v_inst11.count_clk_RNI_0Z0Z_1\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__19619\,
            I => \b2v_inst11.count_clk_RNI_0Z0Z_1\
        );

    \I__2940\ : Odrv4
    port map (
            O => \N__19616\,
            I => \b2v_inst11.count_clk_RNI_0Z0Z_1\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__19609\,
            I => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_1_cascade_\
        );

    \I__2938\ : InMux
    port map (
            O => \N__19606\,
            I => \N__19602\
        );

    \I__2937\ : InMux
    port map (
            O => \N__19605\,
            I => \N__19599\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__19602\,
            I => \N__19596\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__19599\,
            I => \N__19593\
        );

    \I__2934\ : Span4Mux_s2_v
    port map (
            O => \N__19596\,
            I => \N__19590\
        );

    \I__2933\ : Span4Mux_h
    port map (
            O => \N__19593\,
            I => \N__19585\
        );

    \I__2932\ : Span4Mux_h
    port map (
            O => \N__19590\,
            I => \N__19585\
        );

    \I__2931\ : Odrv4
    port map (
            O => \N__19585\,
            I => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_0_0\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__19582\,
            I => \N__19576\
        );

    \I__2929\ : CascadeMux
    port map (
            O => \N__19581\,
            I => \N__19558\
        );

    \I__2928\ : InMux
    port map (
            O => \N__19580\,
            I => \N__19555\
        );

    \I__2927\ : InMux
    port map (
            O => \N__19579\,
            I => \N__19542\
        );

    \I__2926\ : InMux
    port map (
            O => \N__19576\,
            I => \N__19542\
        );

    \I__2925\ : InMux
    port map (
            O => \N__19575\,
            I => \N__19542\
        );

    \I__2924\ : InMux
    port map (
            O => \N__19574\,
            I => \N__19542\
        );

    \I__2923\ : InMux
    port map (
            O => \N__19573\,
            I => \N__19542\
        );

    \I__2922\ : InMux
    port map (
            O => \N__19572\,
            I => \N__19542\
        );

    \I__2921\ : InMux
    port map (
            O => \N__19571\,
            I => \N__19532\
        );

    \I__2920\ : InMux
    port map (
            O => \N__19570\,
            I => \N__19532\
        );

    \I__2919\ : InMux
    port map (
            O => \N__19569\,
            I => \N__19532\
        );

    \I__2918\ : InMux
    port map (
            O => \N__19568\,
            I => \N__19532\
        );

    \I__2917\ : InMux
    port map (
            O => \N__19567\,
            I => \N__19523\
        );

    \I__2916\ : InMux
    port map (
            O => \N__19566\,
            I => \N__19523\
        );

    \I__2915\ : InMux
    port map (
            O => \N__19565\,
            I => \N__19523\
        );

    \I__2914\ : InMux
    port map (
            O => \N__19564\,
            I => \N__19523\
        );

    \I__2913\ : CascadeMux
    port map (
            O => \N__19563\,
            I => \N__19520\
        );

    \I__2912\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19508\
        );

    \I__2911\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19508\
        );

    \I__2910\ : InMux
    port map (
            O => \N__19558\,
            I => \N__19508\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__19555\,
            I => \N__19503\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__19542\,
            I => \N__19503\
        );

    \I__2907\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19500\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__19532\,
            I => \N__19497\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__19523\,
            I => \N__19494\
        );

    \I__2904\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19481\
        );

    \I__2903\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19481\
        );

    \I__2902\ : InMux
    port map (
            O => \N__19518\,
            I => \N__19481\
        );

    \I__2901\ : InMux
    port map (
            O => \N__19517\,
            I => \N__19481\
        );

    \I__2900\ : InMux
    port map (
            O => \N__19516\,
            I => \N__19481\
        );

    \I__2899\ : InMux
    port map (
            O => \N__19515\,
            I => \N__19481\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__19508\,
            I => \N__19478\
        );

    \I__2897\ : Span4Mux_s3_v
    port map (
            O => \N__19503\,
            I => \N__19473\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__19500\,
            I => \N__19473\
        );

    \I__2895\ : Span4Mux_v
    port map (
            O => \N__19497\,
            I => \N__19459\
        );

    \I__2894\ : Span4Mux_s1_v
    port map (
            O => \N__19494\,
            I => \N__19459\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__19481\,
            I => \N__19459\
        );

    \I__2892\ : Span4Mux_h
    port map (
            O => \N__19478\,
            I => \N__19454\
        );

    \I__2891\ : Span4Mux_h
    port map (
            O => \N__19473\,
            I => \N__19454\
        );

    \I__2890\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19439\
        );

    \I__2889\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19439\
        );

    \I__2888\ : InMux
    port map (
            O => \N__19470\,
            I => \N__19439\
        );

    \I__2887\ : InMux
    port map (
            O => \N__19469\,
            I => \N__19439\
        );

    \I__2886\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19439\
        );

    \I__2885\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19439\
        );

    \I__2884\ : InMux
    port map (
            O => \N__19466\,
            I => \N__19439\
        );

    \I__2883\ : Odrv4
    port map (
            O => \N__19459\,
            I => \b2v_inst11.N_122\
        );

    \I__2882\ : Odrv4
    port map (
            O => \N__19454\,
            I => \b2v_inst11.N_122\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__19439\,
            I => \b2v_inst11.N_122\
        );

    \I__2880\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19423\
        );

    \I__2879\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19423\
        );

    \I__2878\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19418\
        );

    \I__2877\ : InMux
    port map (
            O => \N__19429\,
            I => \N__19418\
        );

    \I__2876\ : InMux
    port map (
            O => \N__19428\,
            I => \N__19415\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__19423\,
            I => \N__19412\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__19418\,
            I => \N__19407\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__19415\,
            I => \N__19407\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__19412\,
            I => \b2v_inst11.N_357\
        );

    \I__2871\ : Odrv12
    port map (
            O => \N__19407\,
            I => \b2v_inst11.N_357\
        );

    \I__2870\ : InMux
    port map (
            O => \N__19402\,
            I => \N__19399\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__19399\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__19396\,
            I => \N__19393\
        );

    \I__2867\ : InMux
    port map (
            O => \N__19393\,
            I => \N__19390\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__19390\,
            I => \N__19387\
        );

    \I__2865\ : Odrv4
    port map (
            O => \N__19387\,
            I => \b2v_inst11.un1_func_state25_6_0_a2_0\
        );

    \I__2864\ : InMux
    port map (
            O => \N__19384\,
            I => \N__19381\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__19381\,
            I => \N__19378\
        );

    \I__2862\ : Span4Mux_s3_v
    port map (
            O => \N__19378\,
            I => \N__19375\
        );

    \I__2861\ : Odrv4
    port map (
            O => \N__19375\,
            I => \b2v_inst11.N_327\
        );

    \I__2860\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19369\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__19369\,
            I => \N__19366\
        );

    \I__2858\ : Span4Mux_s3_v
    port map (
            O => \N__19366\,
            I => \N__19363\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__19363\,
            I => \b2v_inst11.N_328\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__19360\,
            I => \b2v_inst11.func_state_1_m0_0_0_0_cascade_\
        );

    \I__2855\ : InMux
    port map (
            O => \N__19357\,
            I => \N__19354\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__19354\,
            I => \N__19351\
        );

    \I__2853\ : Odrv12
    port map (
            O => \N__19351\,
            I => \b2v_inst11.N_354\
        );

    \I__2852\ : CascadeMux
    port map (
            O => \N__19348\,
            I => \b2v_inst11.N_354_cascade_\
        );

    \I__2851\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19341\
        );

    \I__2850\ : CascadeMux
    port map (
            O => \N__19344\,
            I => \N__19334\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__19341\,
            I => \N__19329\
        );

    \I__2848\ : InMux
    port map (
            O => \N__19340\,
            I => \N__19323\
        );

    \I__2847\ : InMux
    port map (
            O => \N__19339\,
            I => \N__19323\
        );

    \I__2846\ : InMux
    port map (
            O => \N__19338\,
            I => \N__19320\
        );

    \I__2845\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19313\
        );

    \I__2844\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19313\
        );

    \I__2843\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19308\
        );

    \I__2842\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19308\
        );

    \I__2841\ : Span4Mux_v
    port map (
            O => \N__19329\,
            I => \N__19305\
        );

    \I__2840\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19302\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__19323\,
            I => \N__19297\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__19320\,
            I => \N__19297\
        );

    \I__2837\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19292\
        );

    \I__2836\ : InMux
    port map (
            O => \N__19318\,
            I => \N__19292\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__19313\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_11\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__19308\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_11\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__19305\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_11\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__19302\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_11\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__19297\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_11\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__19292\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_11\
        );

    \I__2829\ : InMux
    port map (
            O => \N__19279\,
            I => \N__19276\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__19276\,
            I => \b2v_inst11.g2_1_1\
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__19273\,
            I => \b2v_inst11.g3_0_1_cascade_\
        );

    \I__2826\ : InMux
    port map (
            O => \N__19270\,
            I => \N__19267\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__19267\,
            I => \b2v_inst11.N_14_0\
        );

    \I__2824\ : InMux
    port map (
            O => \N__19264\,
            I => \N__19261\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__19261\,
            I => \b2v_inst11.dutycycle_RNI_6Z0Z_5\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__19258\,
            I => \b2v_inst11.dutycycle_RNI_6Z0Z_5_cascade_\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__19255\,
            I => \b2v_inst11.G_6_i_0_cascade_\
        );

    \I__2820\ : InMux
    port map (
            O => \N__19252\,
            I => \N__19249\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__19249\,
            I => \b2v_inst11.G_6_i_a4_1_1\
        );

    \I__2818\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19243\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__19243\,
            I => \b2v_inst11.un1_dutycycle_53_7_1\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__19240\,
            I => \N__19236\
        );

    \I__2815\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19231\
        );

    \I__2814\ : InMux
    port map (
            O => \N__19236\,
            I => \N__19231\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__19231\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__2812\ : InMux
    port map (
            O => \N__19228\,
            I => \N__19222\
        );

    \I__2811\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19222\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__19222\,
            I => \b2v_inst11.dutycycle_RNIGKEF3Z0Z_11\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__19219\,
            I => \b2v_inst11.dutycycleZ0Z_7_cascade_\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__19216\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_\
        );

    \I__2807\ : CascadeMux
    port map (
            O => \N__19213\,
            I => \N__19210\
        );

    \I__2806\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19207\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__19207\,
            I => \N__19204\
        );

    \I__2804\ : Odrv12
    port map (
            O => \N__19204\,
            I => \b2v_inst11.un1_dutycycle_53_8_0\
        );

    \I__2803\ : InMux
    port map (
            O => \N__19201\,
            I => \N__19198\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__19198\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_11\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__19195\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_7_cascade_\
        );

    \I__2800\ : CascadeMux
    port map (
            O => \N__19192\,
            I => \N__19189\
        );

    \I__2799\ : InMux
    port map (
            O => \N__19189\,
            I => \N__19186\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__19186\,
            I => \N__19183\
        );

    \I__2797\ : Odrv12
    port map (
            O => \N__19183\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_12\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__19180\,
            I => \b2v_inst11.m18_i_1_0_cascade_\
        );

    \I__2795\ : InMux
    port map (
            O => \N__19177\,
            I => \N__19174\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__19174\,
            I => \N__19171\
        );

    \I__2793\ : Odrv4
    port map (
            O => \N__19171\,
            I => \b2v_inst11.dutycycle_RNI_11Z0Z_9\
        );

    \I__2792\ : InMux
    port map (
            O => \N__19168\,
            I => \N__19165\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__19165\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_7\
        );

    \I__2790\ : InMux
    port map (
            O => \N__19162\,
            I => \N__19159\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__19159\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_7\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__19156\,
            I => \N__19151\
        );

    \I__2787\ : CascadeMux
    port map (
            O => \N__19155\,
            I => \N__19147\
        );

    \I__2786\ : CascadeMux
    port map (
            O => \N__19154\,
            I => \N__19144\
        );

    \I__2785\ : InMux
    port map (
            O => \N__19151\,
            I => \N__19134\
        );

    \I__2784\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19134\
        );

    \I__2783\ : InMux
    port map (
            O => \N__19147\,
            I => \N__19125\
        );

    \I__2782\ : InMux
    port map (
            O => \N__19144\,
            I => \N__19125\
        );

    \I__2781\ : InMux
    port map (
            O => \N__19143\,
            I => \N__19125\
        );

    \I__2780\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19125\
        );

    \I__2779\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19118\
        );

    \I__2778\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19118\
        );

    \I__2777\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19118\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__19134\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_9\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__19125\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_9\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__19118\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_9\
        );

    \I__2773\ : InMux
    port map (
            O => \N__19111\,
            I => \N__19108\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__19108\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_7\
        );

    \I__2771\ : InMux
    port map (
            O => \N__19105\,
            I => \N__19102\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__19102\,
            I => \b2v_inst11.dutycycle_RNI_8Z0Z_9\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__19099\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_7_cascade_\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__19096\,
            I => \N__19093\
        );

    \I__2767\ : InMux
    port map (
            O => \N__19093\,
            I => \N__19090\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__19090\,
            I => \N__19087\
        );

    \I__2765\ : Odrv12
    port map (
            O => \N__19087\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_11\
        );

    \I__2764\ : InMux
    port map (
            O => \N__19084\,
            I => \N__19081\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__19081\,
            I => \b2v_inst11.un1_dutycycle_53_13_1\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__19078\,
            I => \b2v_inst11.un1_dutycycle_53_39_0_0_1_cascade_\
        );

    \I__2761\ : InMux
    port map (
            O => \N__19075\,
            I => \N__19072\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__19072\,
            I => \b2v_inst11.un1_dutycycle_53_39_0_0\
        );

    \I__2759\ : CascadeMux
    port map (
            O => \N__19069\,
            I => \b2v_inst11.un1_dutycycle_53_39_1_cascade_\
        );

    \I__2758\ : InMux
    port map (
            O => \N__19066\,
            I => \N__19063\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__19063\,
            I => \b2v_inst11.un1_dutycycle_53_41_0\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__19060\,
            I => \N__19057\
        );

    \I__2755\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19054\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__19054\,
            I => \N__19051\
        );

    \I__2753\ : Odrv4
    port map (
            O => \N__19051\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_13\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__19048\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_9_cascade_\
        );

    \I__2751\ : CascadeMux
    port map (
            O => \N__19045\,
            I => \b2v_inst11.un1_dutycycle_53_10_1_0_cascade_\
        );

    \I__2750\ : CascadeMux
    port map (
            O => \N__19042\,
            I => \b2v_inst11.un1_dutycycle_53_44_0_1_cascade_\
        );

    \I__2749\ : CascadeMux
    port map (
            O => \N__19039\,
            I => \b2v_inst11.dutycycle_RNI_6Z0Z_9_cascade_\
        );

    \I__2748\ : CascadeMux
    port map (
            O => \N__19036\,
            I => \N__19033\
        );

    \I__2747\ : InMux
    port map (
            O => \N__19033\,
            I => \N__19030\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__19030\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_11\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__19027\,
            I => \N__19024\
        );

    \I__2744\ : InMux
    port map (
            O => \N__19024\,
            I => \N__19021\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__19021\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_15\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__19018\,
            I => \b2v_inst11.un1_m7_1_0_cascade_\
        );

    \I__2741\ : InMux
    port map (
            O => \N__19015\,
            I => \N__19012\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__19012\,
            I => \N__19008\
        );

    \I__2739\ : InMux
    port map (
            O => \N__19011\,
            I => \N__19005\
        );

    \I__2738\ : Span4Mux_v
    port map (
            O => \N__19008\,
            I => \N__19002\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__19005\,
            I => \b2v_inst11.un1_i3_mux\
        );

    \I__2736\ : Odrv4
    port map (
            O => \N__19002\,
            I => \b2v_inst11.un1_i3_mux\
        );

    \I__2735\ : InMux
    port map (
            O => \N__18997\,
            I => \N__18994\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__18994\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_11\
        );

    \I__2733\ : InMux
    port map (
            O => \N__18991\,
            I => \N__18988\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__18988\,
            I => \b2v_inst11.un1_dutycycle_53_44_0_2_tz\
        );

    \I__2731\ : InMux
    port map (
            O => \N__18985\,
            I => \b2v_inst11.un1_dutycycle_53_cry_11\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__18982\,
            I => \N__18979\
        );

    \I__2729\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18976\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__18976\,
            I => \N__18973\
        );

    \I__2727\ : Span4Mux_v
    port map (
            O => \N__18973\,
            I => \N__18970\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__18970\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_13\
        );

    \I__2725\ : InMux
    port map (
            O => \N__18967\,
            I => \b2v_inst11.un1_dutycycle_53_cry_12\
        );

    \I__2724\ : InMux
    port map (
            O => \N__18964\,
            I => \N__18961\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__18961\,
            I => \N__18958\
        );

    \I__2722\ : Odrv4
    port map (
            O => \N__18958\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_13\
        );

    \I__2721\ : CascadeMux
    port map (
            O => \N__18955\,
            I => \N__18952\
        );

    \I__2720\ : InMux
    port map (
            O => \N__18952\,
            I => \N__18948\
        );

    \I__2719\ : InMux
    port map (
            O => \N__18951\,
            I => \N__18945\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__18948\,
            I => \N__18942\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__18945\,
            I => \b2v_inst11.mult1_un47_sum\
        );

    \I__2716\ : Odrv4
    port map (
            O => \N__18942\,
            I => \b2v_inst11.mult1_un47_sum\
        );

    \I__2715\ : InMux
    port map (
            O => \N__18937\,
            I => \b2v_inst11.un1_dutycycle_53_cry_13\
        );

    \I__2714\ : InMux
    port map (
            O => \N__18934\,
            I => \N__18931\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__18931\,
            I => \N__18928\
        );

    \I__2712\ : Span4Mux_h
    port map (
            O => \N__18928\,
            I => \N__18922\
        );

    \I__2711\ : InMux
    port map (
            O => \N__18927\,
            I => \N__18915\
        );

    \I__2710\ : InMux
    port map (
            O => \N__18926\,
            I => \N__18915\
        );

    \I__2709\ : InMux
    port map (
            O => \N__18925\,
            I => \N__18915\
        );

    \I__2708\ : Odrv4
    port map (
            O => \N__18922\,
            I => \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__18915\,
            I => \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0\
        );

    \I__2706\ : InMux
    port map (
            O => \N__18910\,
            I => \b2v_inst11.un1_dutycycle_53_cry_14\
        );

    \I__2705\ : CascadeMux
    port map (
            O => \N__18907\,
            I => \N__18904\
        );

    \I__2704\ : InMux
    port map (
            O => \N__18904\,
            I => \N__18901\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__18901\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_14\
        );

    \I__2702\ : InMux
    port map (
            O => \N__18898\,
            I => \N__18893\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__18897\,
            I => \N__18890\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__18896\,
            I => \N__18887\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__18893\,
            I => \N__18884\
        );

    \I__2698\ : InMux
    port map (
            O => \N__18890\,
            I => \N__18879\
        );

    \I__2697\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18879\
        );

    \I__2696\ : Span4Mux_h
    port map (
            O => \N__18884\,
            I => \N__18874\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__18879\,
            I => \N__18874\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__18874\,
            I => \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\
        );

    \I__2693\ : InMux
    port map (
            O => \N__18871\,
            I => \bfn_5_9_0_\
        );

    \I__2692\ : InMux
    port map (
            O => \N__18868\,
            I => \b2v_inst11.CO2\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__18865\,
            I => \N__18862\
        );

    \I__2690\ : InMux
    port map (
            O => \N__18862\,
            I => \N__18859\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__18859\,
            I => \N__18855\
        );

    \I__2688\ : InMux
    port map (
            O => \N__18858\,
            I => \N__18852\
        );

    \I__2687\ : Span4Mux_h
    port map (
            O => \N__18855\,
            I => \N__18847\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__18852\,
            I => \N__18847\
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__18847\,
            I => \b2v_inst11.CO2_THRU_CO\
        );

    \I__2684\ : InMux
    port map (
            O => \N__18844\,
            I => \N__18841\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__18841\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_10\
        );

    \I__2682\ : InMux
    port map (
            O => \N__18838\,
            I => \N__18835\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__18835\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_15\
        );

    \I__2680\ : InMux
    port map (
            O => \N__18832\,
            I => \b2v_inst11.un1_dutycycle_53_cry_2_cZ0\
        );

    \I__2679\ : InMux
    port map (
            O => \N__18829\,
            I => \b2v_inst11.un1_dutycycle_53_cry_3_cZ0\
        );

    \I__2678\ : InMux
    port map (
            O => \N__18826\,
            I => \N__18822\
        );

    \I__2677\ : InMux
    port map (
            O => \N__18825\,
            I => \N__18819\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__18822\,
            I => \N__18814\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__18819\,
            I => \N__18814\
        );

    \I__2674\ : Odrv12
    port map (
            O => \N__18814\,
            I => \b2v_inst11.mult1_un110_sum\
        );

    \I__2673\ : InMux
    port map (
            O => \N__18811\,
            I => \b2v_inst11.un1_dutycycle_53_cry_4_cZ0\
        );

    \I__2672\ : InMux
    port map (
            O => \N__18808\,
            I => \N__18804\
        );

    \I__2671\ : InMux
    port map (
            O => \N__18807\,
            I => \N__18801\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__18804\,
            I => \N__18796\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__18801\,
            I => \N__18796\
        );

    \I__2668\ : Odrv12
    port map (
            O => \N__18796\,
            I => \b2v_inst11.mult1_un103_sum\
        );

    \I__2667\ : InMux
    port map (
            O => \N__18793\,
            I => \b2v_inst11.un1_dutycycle_53_cry_5_cZ0\
        );

    \I__2666\ : InMux
    port map (
            O => \N__18790\,
            I => \N__18787\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__18787\,
            I => \N__18784\
        );

    \I__2664\ : Span4Mux_s3_v
    port map (
            O => \N__18784\,
            I => \N__18780\
        );

    \I__2663\ : InMux
    port map (
            O => \N__18783\,
            I => \N__18777\
        );

    \I__2662\ : Odrv4
    port map (
            O => \N__18780\,
            I => \b2v_inst11.mult1_un96_sum\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__18777\,
            I => \b2v_inst11.mult1_un96_sum\
        );

    \I__2660\ : InMux
    port map (
            O => \N__18772\,
            I => \b2v_inst11.un1_dutycycle_53_cry_6_cZ0\
        );

    \I__2659\ : InMux
    port map (
            O => \N__18769\,
            I => \bfn_5_8_0_\
        );

    \I__2658\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18763\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__18763\,
            I => \N__18759\
        );

    \I__2656\ : InMux
    port map (
            O => \N__18762\,
            I => \N__18756\
        );

    \I__2655\ : Sp12to4
    port map (
            O => \N__18759\,
            I => \N__18751\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__18756\,
            I => \N__18751\
        );

    \I__2653\ : Odrv12
    port map (
            O => \N__18751\,
            I => \b2v_inst11.mult1_un82_sum\
        );

    \I__2652\ : InMux
    port map (
            O => \N__18748\,
            I => \b2v_inst11.un1_dutycycle_53_cry_8_cZ0\
        );

    \I__2651\ : InMux
    port map (
            O => \N__18745\,
            I => \N__18742\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__18742\,
            I => \N__18738\
        );

    \I__2649\ : InMux
    port map (
            O => \N__18741\,
            I => \N__18735\
        );

    \I__2648\ : Sp12to4
    port map (
            O => \N__18738\,
            I => \N__18730\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__18735\,
            I => \N__18730\
        );

    \I__2646\ : Odrv12
    port map (
            O => \N__18730\,
            I => \b2v_inst11.mult1_un75_sum\
        );

    \I__2645\ : InMux
    port map (
            O => \N__18727\,
            I => \b2v_inst11.un1_dutycycle_53_cry_9_cZ0\
        );

    \I__2644\ : InMux
    port map (
            O => \N__18724\,
            I => \b2v_inst11.un1_dutycycle_53_cry_10\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__18721\,
            I => \N__18718\
        );

    \I__2642\ : InMux
    port map (
            O => \N__18718\,
            I => \N__18715\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__18715\,
            I => \b2v_inst11.mult1_un47_sum_cry_4_s\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__18712\,
            I => \N__18709\
        );

    \I__2639\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18706\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__18706\,
            I => \b2v_inst11.mult1_un54_sum_cry_5_s\
        );

    \I__2637\ : InMux
    port map (
            O => \N__18703\,
            I => \b2v_inst11.mult1_un54_sum_cry_4\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__18700\,
            I => \N__18697\
        );

    \I__2635\ : InMux
    port map (
            O => \N__18697\,
            I => \N__18694\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__18694\,
            I => \b2v_inst11.mult1_un47_sum_cry_5_s\
        );

    \I__2633\ : InMux
    port map (
            O => \N__18691\,
            I => \N__18688\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__18688\,
            I => \b2v_inst11.mult1_un54_sum_cry_6_s\
        );

    \I__2631\ : InMux
    port map (
            O => \N__18685\,
            I => \b2v_inst11.mult1_un54_sum_cry_5\
        );

    \I__2630\ : InMux
    port map (
            O => \N__18682\,
            I => \N__18679\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__18679\,
            I => \b2v_inst11.mult1_un47_sum_l_fx_6\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__18676\,
            I => \N__18673\
        );

    \I__2627\ : InMux
    port map (
            O => \N__18673\,
            I => \N__18668\
        );

    \I__2626\ : InMux
    port map (
            O => \N__18672\,
            I => \N__18665\
        );

    \I__2625\ : InMux
    port map (
            O => \N__18671\,
            I => \N__18662\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__18668\,
            I => \b2v_inst11.mult1_un47_sum_s_6\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__18665\,
            I => \b2v_inst11.mult1_un47_sum_s_6\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__18662\,
            I => \b2v_inst11.mult1_un47_sum_s_6\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__18655\,
            I => \N__18652\
        );

    \I__2620\ : InMux
    port map (
            O => \N__18652\,
            I => \N__18649\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__18649\,
            I => \b2v_inst11.mult1_un61_sum_axb_8\
        );

    \I__2618\ : InMux
    port map (
            O => \N__18646\,
            I => \b2v_inst11.mult1_un54_sum_cry_6\
        );

    \I__2617\ : InMux
    port map (
            O => \N__18643\,
            I => \N__18640\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__18640\,
            I => \b2v_inst11.mult1_un40_sum_i_5\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__18637\,
            I => \N__18634\
        );

    \I__2614\ : InMux
    port map (
            O => \N__18634\,
            I => \N__18630\
        );

    \I__2613\ : InMux
    port map (
            O => \N__18633\,
            I => \N__18627\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__18630\,
            I => \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__18627\,
            I => \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__2610\ : InMux
    port map (
            O => \N__18622\,
            I => \b2v_inst11.mult1_un54_sum_cry_7\
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__18619\,
            I => \N__18615\
        );

    \I__2608\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18609\
        );

    \I__2607\ : InMux
    port map (
            O => \N__18615\,
            I => \N__18609\
        );

    \I__2606\ : InMux
    port map (
            O => \N__18614\,
            I => \N__18606\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__18609\,
            I => \b2v_inst11.mult1_un54_sum_s_8\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__18606\,
            I => \b2v_inst11.mult1_un54_sum_s_8\
        );

    \I__2603\ : CascadeMux
    port map (
            O => \N__18601\,
            I => \b2v_inst11.mult1_un54_sum_s_8_cascade_\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__18598\,
            I => \N__18594\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__18597\,
            I => \N__18590\
        );

    \I__2600\ : InMux
    port map (
            O => \N__18594\,
            I => \N__18583\
        );

    \I__2599\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18583\
        );

    \I__2598\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18583\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__18583\,
            I => \b2v_inst11.mult1_un54_sum_i_8\
        );

    \I__2596\ : InMux
    port map (
            O => \N__18580\,
            I => \N__18577\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__18577\,
            I => \N__18574\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__18574\,
            I => \N__18571\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__18571\,
            I => \b2v_inst11.m15_e_2\
        );

    \I__2592\ : InMux
    port map (
            O => \N__18568\,
            I => \b2v_inst11.un1_dutycycle_53_cry_0_cZ0\
        );

    \I__2591\ : InMux
    port map (
            O => \N__18565\,
            I => \b2v_inst11.un1_dutycycle_53_cry_1_cZ0\
        );

    \I__2590\ : InMux
    port map (
            O => \N__18562\,
            I => \N__18559\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__18559\,
            I => \b2v_inst11.mult1_un61_sum_cry_4_s\
        );

    \I__2588\ : InMux
    port map (
            O => \N__18556\,
            I => \b2v_inst11.mult1_un61_sum_cry_3\
        );

    \I__2587\ : InMux
    port map (
            O => \N__18553\,
            I => \N__18550\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__18550\,
            I => \b2v_inst11.mult1_un61_sum_cry_5_s\
        );

    \I__2585\ : InMux
    port map (
            O => \N__18547\,
            I => \b2v_inst11.mult1_un61_sum_cry_4\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__18544\,
            I => \N__18541\
        );

    \I__2583\ : InMux
    port map (
            O => \N__18541\,
            I => \N__18538\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__18538\,
            I => \b2v_inst11.mult1_un61_sum_cry_6_s\
        );

    \I__2581\ : InMux
    port map (
            O => \N__18535\,
            I => \b2v_inst11.mult1_un61_sum_cry_5\
        );

    \I__2580\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18529\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__18529\,
            I => \b2v_inst11.mult1_un68_sum_axb_8\
        );

    \I__2578\ : InMux
    port map (
            O => \N__18526\,
            I => \b2v_inst11.mult1_un61_sum_cry_6\
        );

    \I__2577\ : InMux
    port map (
            O => \N__18523\,
            I => \b2v_inst11.mult1_un61_sum_cry_7\
        );

    \I__2576\ : InMux
    port map (
            O => \N__18520\,
            I => \N__18517\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__18517\,
            I => \b2v_inst11.mult1_un47_sum_i\
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__18514\,
            I => \N__18511\
        );

    \I__2573\ : InMux
    port map (
            O => \N__18511\,
            I => \N__18508\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__18508\,
            I => \b2v_inst11.mult1_un54_sum_cry_3_s\
        );

    \I__2571\ : InMux
    port map (
            O => \N__18505\,
            I => \b2v_inst11.mult1_un54_sum_cry_2\
        );

    \I__2570\ : InMux
    port map (
            O => \N__18502\,
            I => \N__18497\
        );

    \I__2569\ : InMux
    port map (
            O => \N__18501\,
            I => \N__18494\
        );

    \I__2568\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18491\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__18497\,
            I => \b2v_inst11.mult1_un47_sum_cry_3_s\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__18494\,
            I => \b2v_inst11.mult1_un47_sum_cry_3_s\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__18491\,
            I => \b2v_inst11.mult1_un47_sum_cry_3_s\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__18484\,
            I => \N__18481\
        );

    \I__2563\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18478\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__18478\,
            I => \b2v_inst11.mult1_un47_sum_l_fx_3\
        );

    \I__2561\ : InMux
    port map (
            O => \N__18475\,
            I => \N__18472\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__18472\,
            I => \b2v_inst11.mult1_un54_sum_cry_4_s\
        );

    \I__2559\ : InMux
    port map (
            O => \N__18469\,
            I => \b2v_inst11.mult1_un54_sum_cry_3\
        );

    \I__2558\ : InMux
    port map (
            O => \N__18466\,
            I => \N__18463\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__18463\,
            I => \b2v_inst11.mult1_un68_sum_cry_3_s\
        );

    \I__2556\ : InMux
    port map (
            O => \N__18460\,
            I => \b2v_inst11.mult1_un68_sum_cry_2_c\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__18457\,
            I => \N__18454\
        );

    \I__2554\ : InMux
    port map (
            O => \N__18454\,
            I => \N__18451\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__18451\,
            I => \b2v_inst11.mult1_un68_sum_cry_4_s\
        );

    \I__2552\ : InMux
    port map (
            O => \N__18448\,
            I => \b2v_inst11.mult1_un68_sum_cry_3_c\
        );

    \I__2551\ : InMux
    port map (
            O => \N__18445\,
            I => \N__18442\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__18442\,
            I => \b2v_inst11.mult1_un68_sum_cry_5_s\
        );

    \I__2549\ : InMux
    port map (
            O => \N__18439\,
            I => \b2v_inst11.mult1_un68_sum_cry_4_c\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__18436\,
            I => \N__18433\
        );

    \I__2547\ : InMux
    port map (
            O => \N__18433\,
            I => \N__18430\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__18430\,
            I => \b2v_inst11.mult1_un68_sum_cry_6_s\
        );

    \I__2545\ : InMux
    port map (
            O => \N__18427\,
            I => \b2v_inst11.mult1_un68_sum_cry_5_c\
        );

    \I__2544\ : InMux
    port map (
            O => \N__18424\,
            I => \N__18421\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__18421\,
            I => \b2v_inst11.mult1_un75_sum_axb_8\
        );

    \I__2542\ : InMux
    port map (
            O => \N__18418\,
            I => \b2v_inst11.mult1_un68_sum_cry_6_c\
        );

    \I__2541\ : InMux
    port map (
            O => \N__18415\,
            I => \b2v_inst11.mult1_un68_sum_cry_7\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__18412\,
            I => \b2v_inst11.mult1_un68_sum_s_8_cascade_\
        );

    \I__2539\ : CascadeMux
    port map (
            O => \N__18409\,
            I => \N__18405\
        );

    \I__2538\ : InMux
    port map (
            O => \N__18408\,
            I => \N__18397\
        );

    \I__2537\ : InMux
    port map (
            O => \N__18405\,
            I => \N__18397\
        );

    \I__2536\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18397\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__18397\,
            I => \b2v_inst11.mult1_un68_sum_i_0_8\
        );

    \I__2534\ : InMux
    port map (
            O => \N__18394\,
            I => \N__18391\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__18391\,
            I => \b2v_inst11.mult1_un61_sum_cry_3_s\
        );

    \I__2532\ : InMux
    port map (
            O => \N__18388\,
            I => \b2v_inst11.mult1_un61_sum_cry_2\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__18385\,
            I => \N__18382\
        );

    \I__2530\ : InMux
    port map (
            O => \N__18382\,
            I => \N__18379\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__18379\,
            I => \b2v_inst11.mult1_un82_sum_i\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__18376\,
            I => \N__18373\
        );

    \I__2527\ : InMux
    port map (
            O => \N__18373\,
            I => \N__18370\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__18370\,
            I => \b2v_inst11.mult1_un75_sum_i\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__18367\,
            I => \N__18364\
        );

    \I__2524\ : InMux
    port map (
            O => \N__18364\,
            I => \N__18361\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__18361\,
            I => \N__18358\
        );

    \I__2522\ : Odrv12
    port map (
            O => \N__18358\,
            I => \b2v_inst11.mult1_un103_sum_i\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__18355\,
            I => \N__18352\
        );

    \I__2520\ : InMux
    port map (
            O => \N__18352\,
            I => \N__18344\
        );

    \I__2519\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18344\
        );

    \I__2518\ : InMux
    port map (
            O => \N__18350\,
            I => \N__18341\
        );

    \I__2517\ : InMux
    port map (
            O => \N__18349\,
            I => \N__18338\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__18344\,
            I => \b2v_inst11.mult1_un103_sum_s_8\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__18341\,
            I => \b2v_inst11.mult1_un103_sum_s_8\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__18338\,
            I => \b2v_inst11.mult1_un103_sum_s_8\
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__18331\,
            I => \N__18328\
        );

    \I__2512\ : InMux
    port map (
            O => \N__18328\,
            I => \N__18319\
        );

    \I__2511\ : InMux
    port map (
            O => \N__18327\,
            I => \N__18319\
        );

    \I__2510\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18319\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__18319\,
            I => \b2v_inst11.mult1_un89_sum_i_0_8\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__18316\,
            I => \N__18313\
        );

    \I__2507\ : InMux
    port map (
            O => \N__18313\,
            I => \N__18310\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__18310\,
            I => \N__18307\
        );

    \I__2505\ : Span4Mux_s3_v
    port map (
            O => \N__18307\,
            I => \N__18304\
        );

    \I__2504\ : Span4Mux_v
    port map (
            O => \N__18304\,
            I => \N__18301\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__18301\,
            I => \b2v_inst11.mult1_un96_sum_i\
        );

    \I__2502\ : InMux
    port map (
            O => \N__18298\,
            I => \N__18295\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__18295\,
            I => \b2v_inst11.mult1_un103_sum_cry_3_s\
        );

    \I__2500\ : InMux
    port map (
            O => \N__18292\,
            I => \b2v_inst11.mult1_un103_sum_cry_2\
        );

    \I__2499\ : InMux
    port map (
            O => \N__18289\,
            I => \N__18286\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__18286\,
            I => \b2v_inst11.mult1_un96_sum_cry_3_s\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__18283\,
            I => \N__18280\
        );

    \I__2496\ : InMux
    port map (
            O => \N__18280\,
            I => \N__18277\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__18277\,
            I => \b2v_inst11.mult1_un103_sum_cry_4_s\
        );

    \I__2494\ : InMux
    port map (
            O => \N__18274\,
            I => \b2v_inst11.mult1_un103_sum_cry_3\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__18271\,
            I => \N__18268\
        );

    \I__2492\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18265\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__18265\,
            I => \b2v_inst11.mult1_un96_sum_cry_4_s\
        );

    \I__2490\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18259\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__18259\,
            I => \b2v_inst11.mult1_un103_sum_cry_5_s\
        );

    \I__2488\ : InMux
    port map (
            O => \N__18256\,
            I => \b2v_inst11.mult1_un103_sum_cry_4\
        );

    \I__2487\ : InMux
    port map (
            O => \N__18253\,
            I => \N__18250\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__18250\,
            I => \b2v_inst11.mult1_un96_sum_cry_5_s\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__18247\,
            I => \N__18244\
        );

    \I__2484\ : InMux
    port map (
            O => \N__18244\,
            I => \N__18241\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__18241\,
            I => \b2v_inst11.mult1_un103_sum_cry_6_s\
        );

    \I__2482\ : InMux
    port map (
            O => \N__18238\,
            I => \b2v_inst11.mult1_un103_sum_cry_5\
        );

    \I__2481\ : CascadeMux
    port map (
            O => \N__18235\,
            I => \N__18231\
        );

    \I__2480\ : InMux
    port map (
            O => \N__18234\,
            I => \N__18223\
        );

    \I__2479\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18223\
        );

    \I__2478\ : InMux
    port map (
            O => \N__18230\,
            I => \N__18223\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__18223\,
            I => \b2v_inst11.mult1_un96_sum_i_0_8\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__18220\,
            I => \N__18217\
        );

    \I__2475\ : InMux
    port map (
            O => \N__18217\,
            I => \N__18214\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__18214\,
            I => \b2v_inst11.mult1_un96_sum_cry_6_s\
        );

    \I__2473\ : InMux
    port map (
            O => \N__18211\,
            I => \N__18208\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__18208\,
            I => \b2v_inst11.mult1_un110_sum_axb_8\
        );

    \I__2471\ : InMux
    port map (
            O => \N__18205\,
            I => \b2v_inst11.mult1_un103_sum_cry_6\
        );

    \I__2470\ : InMux
    port map (
            O => \N__18202\,
            I => \N__18199\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__18199\,
            I => \b2v_inst11.mult1_un103_sum_axb_8\
        );

    \I__2468\ : InMux
    port map (
            O => \N__18196\,
            I => \b2v_inst11.mult1_un103_sum_cry_7\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__18193\,
            I => \b2v_inst11.mult1_un103_sum_s_8_cascade_\
        );

    \I__2466\ : CascadeMux
    port map (
            O => \N__18190\,
            I => \N__18186\
        );

    \I__2465\ : InMux
    port map (
            O => \N__18189\,
            I => \N__18178\
        );

    \I__2464\ : InMux
    port map (
            O => \N__18186\,
            I => \N__18178\
        );

    \I__2463\ : InMux
    port map (
            O => \N__18185\,
            I => \N__18178\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__18178\,
            I => \b2v_inst11.mult1_un103_sum_i_0_8\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__18175\,
            I => \N__18172\
        );

    \I__2460\ : InMux
    port map (
            O => \N__18172\,
            I => \N__18169\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__18169\,
            I => \N__18166\
        );

    \I__2458\ : Odrv4
    port map (
            O => \N__18166\,
            I => \b2v_inst11.count_off_0_13\
        );

    \I__2457\ : CascadeMux
    port map (
            O => \N__18163\,
            I => \N__18159\
        );

    \I__2456\ : InMux
    port map (
            O => \N__18162\,
            I => \N__18144\
        );

    \I__2455\ : InMux
    port map (
            O => \N__18159\,
            I => \N__18144\
        );

    \I__2454\ : CEMux
    port map (
            O => \N__18158\,
            I => \N__18144\
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__18157\,
            I => \N__18140\
        );

    \I__2452\ : CEMux
    port map (
            O => \N__18156\,
            I => \N__18127\
        );

    \I__2451\ : InMux
    port map (
            O => \N__18155\,
            I => \N__18120\
        );

    \I__2450\ : InMux
    port map (
            O => \N__18154\,
            I => \N__18120\
        );

    \I__2449\ : CEMux
    port map (
            O => \N__18153\,
            I => \N__18120\
        );

    \I__2448\ : InMux
    port map (
            O => \N__18152\,
            I => \N__18115\
        );

    \I__2447\ : CEMux
    port map (
            O => \N__18151\,
            I => \N__18115\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__18144\,
            I => \N__18112\
        );

    \I__2445\ : InMux
    port map (
            O => \N__18143\,
            I => \N__18109\
        );

    \I__2444\ : InMux
    port map (
            O => \N__18140\,
            I => \N__18106\
        );

    \I__2443\ : InMux
    port map (
            O => \N__18139\,
            I => \N__18103\
        );

    \I__2442\ : InMux
    port map (
            O => \N__18138\,
            I => \N__18097\
        );

    \I__2441\ : InMux
    port map (
            O => \N__18137\,
            I => \N__18094\
        );

    \I__2440\ : InMux
    port map (
            O => \N__18136\,
            I => \N__18083\
        );

    \I__2439\ : CEMux
    port map (
            O => \N__18135\,
            I => \N__18083\
        );

    \I__2438\ : InMux
    port map (
            O => \N__18134\,
            I => \N__18083\
        );

    \I__2437\ : InMux
    port map (
            O => \N__18133\,
            I => \N__18083\
        );

    \I__2436\ : InMux
    port map (
            O => \N__18132\,
            I => \N__18083\
        );

    \I__2435\ : InMux
    port map (
            O => \N__18131\,
            I => \N__18078\
        );

    \I__2434\ : InMux
    port map (
            O => \N__18130\,
            I => \N__18078\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__18127\,
            I => \N__18074\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__18120\,
            I => \N__18071\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__18115\,
            I => \N__18068\
        );

    \I__2430\ : Span4Mux_s2_v
    port map (
            O => \N__18112\,
            I => \N__18065\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__18109\,
            I => \N__18062\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__18106\,
            I => \N__18057\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__18103\,
            I => \N__18057\
        );

    \I__2426\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18050\
        );

    \I__2425\ : InMux
    port map (
            O => \N__18101\,
            I => \N__18050\
        );

    \I__2424\ : InMux
    port map (
            O => \N__18100\,
            I => \N__18050\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__18097\,
            I => \N__18047\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__18094\,
            I => \N__18042\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__18083\,
            I => \N__18042\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__18078\,
            I => \N__18039\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__18077\,
            I => \N__18034\
        );

    \I__2418\ : Span4Mux_s3_h
    port map (
            O => \N__18074\,
            I => \N__18030\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__18071\,
            I => \N__18027\
        );

    \I__2416\ : Span4Mux_s2_h
    port map (
            O => \N__18068\,
            I => \N__18018\
        );

    \I__2415\ : Span4Mux_s2_h
    port map (
            O => \N__18065\,
            I => \N__18018\
        );

    \I__2414\ : Span4Mux_s2_v
    port map (
            O => \N__18062\,
            I => \N__18018\
        );

    \I__2413\ : Span4Mux_s2_v
    port map (
            O => \N__18057\,
            I => \N__18018\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__18050\,
            I => \N__18011\
        );

    \I__2411\ : Span4Mux_v
    port map (
            O => \N__18047\,
            I => \N__18011\
        );

    \I__2410\ : Span4Mux_s2_v
    port map (
            O => \N__18042\,
            I => \N__18011\
        );

    \I__2409\ : Span4Mux_s3_h
    port map (
            O => \N__18039\,
            I => \N__18008\
        );

    \I__2408\ : InMux
    port map (
            O => \N__18038\,
            I => \N__17999\
        );

    \I__2407\ : CEMux
    port map (
            O => \N__18037\,
            I => \N__17999\
        );

    \I__2406\ : InMux
    port map (
            O => \N__18034\,
            I => \N__17999\
        );

    \I__2405\ : InMux
    port map (
            O => \N__18033\,
            I => \N__17999\
        );

    \I__2404\ : Odrv4
    port map (
            O => \N__18030\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__18027\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__18018\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__18011\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__2400\ : Odrv4
    port map (
            O => \N__18008\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__17999\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__2398\ : InMux
    port map (
            O => \N__17986\,
            I => \N__17983\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__17983\,
            I => \N__17980\
        );

    \I__2396\ : Odrv12
    port map (
            O => \N__17980\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2\
        );

    \I__2395\ : InMux
    port map (
            O => \N__17977\,
            I => \b2v_inst11.mult1_un110_sum_cry_2\
        );

    \I__2394\ : InMux
    port map (
            O => \N__17974\,
            I => \b2v_inst11.mult1_un110_sum_cry_3\
        );

    \I__2393\ : InMux
    port map (
            O => \N__17971\,
            I => \b2v_inst11.mult1_un110_sum_cry_4\
        );

    \I__2392\ : InMux
    port map (
            O => \N__17968\,
            I => \b2v_inst11.mult1_un110_sum_cry_5\
        );

    \I__2391\ : InMux
    port map (
            O => \N__17965\,
            I => \b2v_inst11.mult1_un110_sum_cry_6\
        );

    \I__2390\ : InMux
    port map (
            O => \N__17962\,
            I => \b2v_inst11.mult1_un110_sum_cry_7\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__17959\,
            I => \N__17955\
        );

    \I__2388\ : InMux
    port map (
            O => \N__17958\,
            I => \N__17949\
        );

    \I__2387\ : InMux
    port map (
            O => \N__17955\,
            I => \N__17944\
        );

    \I__2386\ : InMux
    port map (
            O => \N__17954\,
            I => \N__17944\
        );

    \I__2385\ : InMux
    port map (
            O => \N__17953\,
            I => \N__17941\
        );

    \I__2384\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17938\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__17949\,
            I => \b2v_inst11.mult1_un89_sum_s_8\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__17944\,
            I => \b2v_inst11.mult1_un89_sum_s_8\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__17941\,
            I => \b2v_inst11.mult1_un89_sum_s_8\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__17938\,
            I => \b2v_inst11.mult1_un89_sum_s_8\
        );

    \I__2379\ : InMux
    port map (
            O => \N__17929\,
            I => \N__17926\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__17926\,
            I => \N__17923\
        );

    \I__2377\ : Span4Mux_s2_h
    port map (
            O => \N__17923\,
            I => \N__17920\
        );

    \I__2376\ : Span4Mux_v
    port map (
            O => \N__17920\,
            I => \N__17917\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__17917\,
            I => \b2v_inst11.N_322\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__17914\,
            I => \b2v_inst11.count_offZ0Z_0_cascade_\
        );

    \I__2373\ : InMux
    port map (
            O => \N__17911\,
            I => \N__17907\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__17910\,
            I => \N__17904\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__17907\,
            I => \N__17901\
        );

    \I__2370\ : InMux
    port map (
            O => \N__17904\,
            I => \N__17898\
        );

    \I__2369\ : Span4Mux_v
    port map (
            O => \N__17901\,
            I => \N__17894\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__17898\,
            I => \N__17891\
        );

    \I__2367\ : InMux
    port map (
            O => \N__17897\,
            I => \N__17888\
        );

    \I__2366\ : Span4Mux_s1_v
    port map (
            O => \N__17894\,
            I => \N__17883\
        );

    \I__2365\ : Span4Mux_v
    port map (
            O => \N__17891\,
            I => \N__17883\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__17888\,
            I => \b2v_inst11.count_offZ0Z_1\
        );

    \I__2363\ : Odrv4
    port map (
            O => \N__17883\,
            I => \b2v_inst11.count_offZ0Z_1\
        );

    \I__2362\ : InMux
    port map (
            O => \N__17878\,
            I => \N__17875\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__17875\,
            I => \b2v_inst11.count_off_RNIZ0Z_1\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__17872\,
            I => \b2v_inst11.count_off_RNIZ0Z_1_cascade_\
        );

    \I__2359\ : InMux
    port map (
            O => \N__17869\,
            I => \N__17866\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__17866\,
            I => \b2v_inst11.count_off_0_1\
        );

    \I__2357\ : InMux
    port map (
            O => \N__17863\,
            I => \N__17859\
        );

    \I__2356\ : InMux
    port map (
            O => \N__17862\,
            I => \N__17856\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__17859\,
            I => \N__17853\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__17856\,
            I => \N__17849\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__17853\,
            I => \N__17846\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__17852\,
            I => \N__17842\
        );

    \I__2351\ : Span4Mux_s1_v
    port map (
            O => \N__17849\,
            I => \N__17837\
        );

    \I__2350\ : Span4Mux_s1_h
    port map (
            O => \N__17846\,
            I => \N__17837\
        );

    \I__2349\ : InMux
    port map (
            O => \N__17845\,
            I => \N__17832\
        );

    \I__2348\ : InMux
    port map (
            O => \N__17842\,
            I => \N__17832\
        );

    \I__2347\ : Odrv4
    port map (
            O => \N__17837\,
            I => \b2v_inst11.count_offZ0Z_0\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__17832\,
            I => \b2v_inst11.count_offZ0Z_0\
        );

    \I__2345\ : InMux
    port map (
            O => \N__17827\,
            I => \N__17824\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__17824\,
            I => \b2v_inst11.count_off_0_0\
        );

    \I__2343\ : InMux
    port map (
            O => \N__17821\,
            I => \N__17818\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__17818\,
            I => \b2v_inst11.count_off_0_10\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__17815\,
            I => \N__17812\
        );

    \I__2340\ : InMux
    port map (
            O => \N__17812\,
            I => \N__17806\
        );

    \I__2339\ : InMux
    port map (
            O => \N__17811\,
            I => \N__17806\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__17806\,
            I => \N__17803\
        );

    \I__2337\ : Odrv4
    port map (
            O => \N__17803\,
            I => \b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__17800\,
            I => \N__17796\
        );

    \I__2335\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17793\
        );

    \I__2334\ : InMux
    port map (
            O => \N__17796\,
            I => \N__17790\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__17793\,
            I => \N__17787\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__17790\,
            I => \N__17784\
        );

    \I__2331\ : Span4Mux_s3_h
    port map (
            O => \N__17787\,
            I => \N__17781\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__17784\,
            I => \b2v_inst11.count_offZ0Z_10\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__17781\,
            I => \b2v_inst11.count_offZ0Z_10\
        );

    \I__2328\ : InMux
    port map (
            O => \N__17776\,
            I => \N__17773\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__17773\,
            I => \N__17769\
        );

    \I__2326\ : InMux
    port map (
            O => \N__17772\,
            I => \N__17766\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__17769\,
            I => \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__17766\,
            I => \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5\
        );

    \I__2323\ : InMux
    port map (
            O => \N__17761\,
            I => \N__17758\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__17758\,
            I => \b2v_inst11.dutycycle_RNIGKEF3Z0Z_12\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__17755\,
            I => \N__17752\
        );

    \I__2320\ : InMux
    port map (
            O => \N__17752\,
            I => \N__17746\
        );

    \I__2319\ : InMux
    port map (
            O => \N__17751\,
            I => \N__17746\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__17746\,
            I => \b2v_inst11.dutycycleZ1Z_12\
        );

    \I__2317\ : CascadeMux
    port map (
            O => \N__17743\,
            I => \b2v_inst11.dutycycle_RNIGKEF3Z0Z_12_cascade_\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__17740\,
            I => \b2v_inst11.dutycycleZ0Z_10_cascade_\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__17737\,
            I => \b2v_inst11.un1_dutycycle_53_56_a0_3_0_cascade_\
        );

    \I__2314\ : InMux
    port map (
            O => \N__17734\,
            I => \N__17728\
        );

    \I__2313\ : InMux
    port map (
            O => \N__17733\,
            I => \N__17728\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__17728\,
            I => \b2v_inst11.N_232_N\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__17725\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_325_N_cascade_\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__17722\,
            I => \b2v_inst11.un1_func_state25_6_0_1_cascade_\
        );

    \I__2309\ : InMux
    port map (
            O => \N__17719\,
            I => \N__17716\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__17716\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_323_N\
        );

    \I__2307\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17710\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__17710\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_324_N\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__17707\,
            I => \b2v_inst11.N_289_cascade_\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__17704\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_0_2_cascade_\
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__17701\,
            I => \b2v_inst11.N_302_cascade_\
        );

    \I__2302\ : CascadeMux
    port map (
            O => \N__17698\,
            I => \b2v_inst11.N_301_cascade_\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__17695\,
            I => \b2v_inst11.dutycycle_RNIJU083Z0Z_8_cascade_\
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__17692\,
            I => \b2v_inst11.N_108_f0_cascade_\
        );

    \I__2299\ : InMux
    port map (
            O => \N__17689\,
            I => \N__17686\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__17686\,
            I => \b2v_inst11.dutycycle_RNIHTFQZ0Z_8\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__17683\,
            I => \b2v_inst11.dutycycle_RNI2NK31Z0Z_8_cascade_\
        );

    \I__2296\ : InMux
    port map (
            O => \N__17680\,
            I => \N__17677\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__17677\,
            I => \b2v_inst11.dutycycle_e_1_8\
        );

    \I__2294\ : InMux
    port map (
            O => \N__17674\,
            I => \N__17662\
        );

    \I__2293\ : InMux
    port map (
            O => \N__17673\,
            I => \N__17662\
        );

    \I__2292\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17662\
        );

    \I__2291\ : InMux
    port map (
            O => \N__17671\,
            I => \N__17662\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__17662\,
            I => \b2v_inst11.dutycycleZ1Z_8\
        );

    \I__2289\ : InMux
    port map (
            O => \N__17659\,
            I => \N__17656\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__17656\,
            I => \b2v_inst11.N_108_f0\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__17653\,
            I => \b2v_inst11.dutycycle_e_1_8_cascade_\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__17650\,
            I => \b2v_inst11.dutycycleZ0Z_1_cascade_\
        );

    \I__2285\ : InMux
    port map (
            O => \N__17647\,
            I => \N__17644\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__17644\,
            I => \b2v_inst11.dutycycle_RNIJU083_0Z0Z_8\
        );

    \I__2283\ : IoInMux
    port map (
            O => \N__17641\,
            I => \N__17637\
        );

    \I__2282\ : IoInMux
    port map (
            O => \N__17640\,
            I => \N__17634\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__17637\,
            I => \N__17629\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__17634\,
            I => \N__17629\
        );

    \I__2279\ : IoSpan4Mux
    port map (
            O => \N__17629\,
            I => \N__17626\
        );

    \I__2278\ : Span4Mux_s0_h
    port map (
            O => \N__17626\,
            I => \N__17622\
        );

    \I__2277\ : IoInMux
    port map (
            O => \N__17625\,
            I => \N__17619\
        );

    \I__2276\ : Sp12to4
    port map (
            O => \N__17622\,
            I => \N__17614\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__17619\,
            I => \N__17614\
        );

    \I__2274\ : Odrv12
    port map (
            O => \N__17614\,
            I => \delayed_vccin_vccinaux_ok_RNIM6F44_0\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__17611\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_12_cascade_\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__17608\,
            I => \b2v_inst11.dutycycle_RNI_10Z0Z_9_cascade_\
        );

    \I__2271\ : InMux
    port map (
            O => \N__17605\,
            I => \N__17599\
        );

    \I__2270\ : InMux
    port map (
            O => \N__17604\,
            I => \N__17599\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__17599\,
            I => \b2v_inst11.dutycycle_en_10\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__17596\,
            I => \N__17592\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__17595\,
            I => \N__17589\
        );

    \I__2266\ : InMux
    port map (
            O => \N__17592\,
            I => \N__17584\
        );

    \I__2265\ : InMux
    port map (
            O => \N__17589\,
            I => \N__17584\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__17584\,
            I => \b2v_inst11.dutycycleZ1Z_13\
        );

    \I__2263\ : CascadeMux
    port map (
            O => \N__17581\,
            I => \b2v_inst11.dutycycleZ0Z_9_cascade_\
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__17578\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_13_cascade_\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__17575\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_10_cascade_\
        );

    \I__2260\ : InMux
    port map (
            O => \N__17572\,
            I => \N__17569\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__17569\,
            I => \N__17566\
        );

    \I__2258\ : Span4Mux_v
    port map (
            O => \N__17566\,
            I => \N__17562\
        );

    \I__2257\ : InMux
    port map (
            O => \N__17565\,
            I => \N__17559\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__17562\,
            I => \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__17559\,
            I => \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5\
        );

    \I__2254\ : InMux
    port map (
            O => \N__17554\,
            I => \N__17551\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__17551\,
            I => \N__17548\
        );

    \I__2252\ : Span4Mux_s3_h
    port map (
            O => \N__17548\,
            I => \N__17545\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__17545\,
            I => \b2v_inst11.count_clk_0_3\
        );

    \I__2250\ : CEMux
    port map (
            O => \N__17542\,
            I => \N__17539\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__17539\,
            I => \N__17534\
        );

    \I__2248\ : CEMux
    port map (
            O => \N__17538\,
            I => \N__17531\
        );

    \I__2247\ : CEMux
    port map (
            O => \N__17537\,
            I => \N__17528\
        );

    \I__2246\ : Span4Mux_s2_h
    port map (
            O => \N__17534\,
            I => \N__17520\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__17531\,
            I => \N__17515\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__17528\,
            I => \N__17515\
        );

    \I__2243\ : CEMux
    port map (
            O => \N__17527\,
            I => \N__17512\
        );

    \I__2242\ : CEMux
    port map (
            O => \N__17526\,
            I => \N__17508\
        );

    \I__2241\ : InMux
    port map (
            O => \N__17525\,
            I => \N__17501\
        );

    \I__2240\ : InMux
    port map (
            O => \N__17524\,
            I => \N__17501\
        );

    \I__2239\ : InMux
    port map (
            O => \N__17523\,
            I => \N__17501\
        );

    \I__2238\ : Span4Mux_v
    port map (
            O => \N__17520\,
            I => \N__17496\
        );

    \I__2237\ : Span4Mux_v
    port map (
            O => \N__17515\,
            I => \N__17489\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__17512\,
            I => \N__17489\
        );

    \I__2235\ : CEMux
    port map (
            O => \N__17511\,
            I => \N__17486\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__17508\,
            I => \N__17477\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__17501\,
            I => \N__17474\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__17500\,
            I => \N__17471\
        );

    \I__2231\ : CascadeMux
    port map (
            O => \N__17499\,
            I => \N__17468\
        );

    \I__2230\ : IoSpan4Mux
    port map (
            O => \N__17496\,
            I => \N__17463\
        );

    \I__2229\ : InMux
    port map (
            O => \N__17495\,
            I => \N__17458\
        );

    \I__2228\ : InMux
    port map (
            O => \N__17494\,
            I => \N__17458\
        );

    \I__2227\ : Span4Mux_h
    port map (
            O => \N__17489\,
            I => \N__17455\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__17486\,
            I => \N__17452\
        );

    \I__2225\ : InMux
    port map (
            O => \N__17485\,
            I => \N__17447\
        );

    \I__2224\ : InMux
    port map (
            O => \N__17484\,
            I => \N__17447\
        );

    \I__2223\ : InMux
    port map (
            O => \N__17483\,
            I => \N__17438\
        );

    \I__2222\ : InMux
    port map (
            O => \N__17482\,
            I => \N__17438\
        );

    \I__2221\ : InMux
    port map (
            O => \N__17481\,
            I => \N__17438\
        );

    \I__2220\ : InMux
    port map (
            O => \N__17480\,
            I => \N__17438\
        );

    \I__2219\ : Span4Mux_h
    port map (
            O => \N__17477\,
            I => \N__17433\
        );

    \I__2218\ : Span4Mux_s2_h
    port map (
            O => \N__17474\,
            I => \N__17433\
        );

    \I__2217\ : InMux
    port map (
            O => \N__17471\,
            I => \N__17430\
        );

    \I__2216\ : InMux
    port map (
            O => \N__17468\,
            I => \N__17423\
        );

    \I__2215\ : InMux
    port map (
            O => \N__17467\,
            I => \N__17423\
        );

    \I__2214\ : InMux
    port map (
            O => \N__17466\,
            I => \N__17423\
        );

    \I__2213\ : Span4Mux_s3_v
    port map (
            O => \N__17463\,
            I => \N__17418\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__17458\,
            I => \N__17418\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__17455\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2210\ : Odrv12
    port map (
            O => \N__17452\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__17447\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__17438\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2207\ : Odrv4
    port map (
            O => \N__17433\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__17430\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__17423\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2204\ : Odrv4
    port map (
            O => \N__17418\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__17401\,
            I => \N__17398\
        );

    \I__2202\ : InMux
    port map (
            O => \N__17398\,
            I => \N__17395\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__17395\,
            I => \b2v_inst11.N_150_N\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__17392\,
            I => \b2v_inst11.N_152_N_cascade_\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__17389\,
            I => \b2v_inst11.dutycycleZ0Z_12_cascade_\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__17386\,
            I => \b2v_inst11.N_155_N_cascade_\
        );

    \I__2197\ : InMux
    port map (
            O => \N__17383\,
            I => \N__17380\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__17380\,
            I => \b2v_inst11.dutycycle_en_12\
        );

    \I__2195\ : CascadeMux
    port map (
            O => \N__17377\,
            I => \b2v_inst11.dutycycle_en_12_cascade_\
        );

    \I__2194\ : InMux
    port map (
            O => \N__17374\,
            I => \N__17370\
        );

    \I__2193\ : InMux
    port map (
            O => \N__17373\,
            I => \N__17367\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__17370\,
            I => \b2v_inst11.dutycycleZ0Z_15\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__17367\,
            I => \b2v_inst11.dutycycleZ0Z_15\
        );

    \I__2190\ : IoInMux
    port map (
            O => \N__17362\,
            I => \N__17359\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__17359\,
            I => \N__17356\
        );

    \I__2188\ : Span4Mux_s3_h
    port map (
            O => \N__17356\,
            I => \N__17353\
        );

    \I__2187\ : Odrv4
    port map (
            O => \N__17353\,
            I => \b2v_inst200.count_enZ0\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__17350\,
            I => \N__17347\
        );

    \I__2185\ : InMux
    port map (
            O => \N__17347\,
            I => \N__17344\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__17344\,
            I => \b2v_inst11.un1_dutycycle_53_i_29\
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__17341\,
            I => \N__17338\
        );

    \I__2182\ : InMux
    port map (
            O => \N__17338\,
            I => \N__17335\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__17335\,
            I => \b2v_inst11.mult1_un40_sum_i_l_ofx_4\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__17332\,
            I => \N__17329\
        );

    \I__2179\ : InMux
    port map (
            O => \N__17329\,
            I => \N__17326\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__17326\,
            I => \b2v_inst11.mult1_un47_sum_s_4_sf\
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__17323\,
            I => \b2v_inst11.mult1_un40_sum_i_5_cascade_\
        );

    \I__2176\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17316\
        );

    \I__2175\ : InMux
    port map (
            O => \N__17319\,
            I => \N__17313\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__17316\,
            I => \N__17310\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__17313\,
            I => \N__17307\
        );

    \I__2172\ : Span4Mux_s3_h
    port map (
            O => \N__17310\,
            I => \N__17304\
        );

    \I__2171\ : Span4Mux_s3_h
    port map (
            O => \N__17307\,
            I => \N__17301\
        );

    \I__2170\ : Odrv4
    port map (
            O => \N__17304\,
            I => \b2v_inst16.countZ0Z_10\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__17301\,
            I => \b2v_inst16.countZ0Z_10\
        );

    \I__2168\ : InMux
    port map (
            O => \N__17296\,
            I => \N__17290\
        );

    \I__2167\ : InMux
    port map (
            O => \N__17295\,
            I => \N__17290\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__17290\,
            I => \N__17287\
        );

    \I__2165\ : Span4Mux_h
    port map (
            O => \N__17287\,
            I => \N__17284\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__17284\,
            I => \b2v_inst16.count_rst\
        );

    \I__2163\ : InMux
    port map (
            O => \N__17281\,
            I => \N__17278\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__17278\,
            I => \b2v_inst16.count_4_10\
        );

    \I__2161\ : InMux
    port map (
            O => \N__17275\,
            I => \b2v_inst11.mult1_un47_sum_cry_2\
        );

    \I__2160\ : InMux
    port map (
            O => \N__17272\,
            I => \b2v_inst11.mult1_un47_sum_cry_3\
        );

    \I__2159\ : InMux
    port map (
            O => \N__17269\,
            I => \b2v_inst11.mult1_un47_sum_cry_4\
        );

    \I__2158\ : InMux
    port map (
            O => \N__17266\,
            I => \b2v_inst11.mult1_un47_sum_cry_5\
        );

    \I__2157\ : InMux
    port map (
            O => \N__17263\,
            I => \N__17260\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__17260\,
            I => \b2v_inst11.mult1_un75_sum_cry_3_s\
        );

    \I__2155\ : InMux
    port map (
            O => \N__17257\,
            I => \b2v_inst11.mult1_un75_sum_cry_2\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__17254\,
            I => \N__17251\
        );

    \I__2153\ : InMux
    port map (
            O => \N__17251\,
            I => \N__17248\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__17248\,
            I => \b2v_inst11.mult1_un75_sum_cry_4_s\
        );

    \I__2151\ : InMux
    port map (
            O => \N__17245\,
            I => \b2v_inst11.mult1_un75_sum_cry_3\
        );

    \I__2150\ : InMux
    port map (
            O => \N__17242\,
            I => \N__17239\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__17239\,
            I => \b2v_inst11.mult1_un75_sum_cry_5_s\
        );

    \I__2148\ : InMux
    port map (
            O => \N__17236\,
            I => \b2v_inst11.mult1_un75_sum_cry_4\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__17233\,
            I => \N__17230\
        );

    \I__2146\ : InMux
    port map (
            O => \N__17230\,
            I => \N__17227\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__17227\,
            I => \b2v_inst11.mult1_un75_sum_cry_6_s\
        );

    \I__2144\ : InMux
    port map (
            O => \N__17224\,
            I => \b2v_inst11.mult1_un75_sum_cry_5\
        );

    \I__2143\ : InMux
    port map (
            O => \N__17221\,
            I => \N__17218\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__17218\,
            I => \b2v_inst11.mult1_un82_sum_axb_8\
        );

    \I__2141\ : InMux
    port map (
            O => \N__17215\,
            I => \b2v_inst11.mult1_un75_sum_cry_6\
        );

    \I__2140\ : InMux
    port map (
            O => \N__17212\,
            I => \b2v_inst11.mult1_un75_sum_cry_7\
        );

    \I__2139\ : CascadeMux
    port map (
            O => \N__17209\,
            I => \b2v_inst11.mult1_un75_sum_s_8_cascade_\
        );

    \I__2138\ : CascadeMux
    port map (
            O => \N__17206\,
            I => \N__17202\
        );

    \I__2137\ : InMux
    port map (
            O => \N__17205\,
            I => \N__17194\
        );

    \I__2136\ : InMux
    port map (
            O => \N__17202\,
            I => \N__17194\
        );

    \I__2135\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17194\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__17194\,
            I => \b2v_inst11.mult1_un75_sum_i_0_8\
        );

    \I__2133\ : InMux
    port map (
            O => \N__17191\,
            I => \b2v_inst11.mult1_un89_sum_cry_7\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__17188\,
            I => \N__17184\
        );

    \I__2131\ : InMux
    port map (
            O => \N__17187\,
            I => \N__17176\
        );

    \I__2130\ : InMux
    port map (
            O => \N__17184\,
            I => \N__17176\
        );

    \I__2129\ : InMux
    port map (
            O => \N__17183\,
            I => \N__17176\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__17176\,
            I => \b2v_inst11.mult1_un82_sum_i_0_8\
        );

    \I__2127\ : InMux
    port map (
            O => \N__17173\,
            I => \N__17170\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__17170\,
            I => \b2v_inst11.mult1_un82_sum_cry_3_s\
        );

    \I__2125\ : InMux
    port map (
            O => \N__17167\,
            I => \b2v_inst11.mult1_un82_sum_cry_2\
        );

    \I__2124\ : CascadeMux
    port map (
            O => \N__17164\,
            I => \N__17161\
        );

    \I__2123\ : InMux
    port map (
            O => \N__17161\,
            I => \N__17158\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__17158\,
            I => \b2v_inst11.mult1_un82_sum_cry_4_s\
        );

    \I__2121\ : InMux
    port map (
            O => \N__17155\,
            I => \b2v_inst11.mult1_un82_sum_cry_3\
        );

    \I__2120\ : InMux
    port map (
            O => \N__17152\,
            I => \N__17149\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__17149\,
            I => \b2v_inst11.mult1_un82_sum_cry_5_s\
        );

    \I__2118\ : InMux
    port map (
            O => \N__17146\,
            I => \b2v_inst11.mult1_un82_sum_cry_4\
        );

    \I__2117\ : CascadeMux
    port map (
            O => \N__17143\,
            I => \N__17140\
        );

    \I__2116\ : InMux
    port map (
            O => \N__17140\,
            I => \N__17137\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__17137\,
            I => \b2v_inst11.mult1_un82_sum_cry_6_s\
        );

    \I__2114\ : InMux
    port map (
            O => \N__17134\,
            I => \b2v_inst11.mult1_un82_sum_cry_5\
        );

    \I__2113\ : InMux
    port map (
            O => \N__17131\,
            I => \N__17128\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__17128\,
            I => \b2v_inst11.mult1_un89_sum_axb_8\
        );

    \I__2111\ : InMux
    port map (
            O => \N__17125\,
            I => \b2v_inst11.mult1_un82_sum_cry_6\
        );

    \I__2110\ : InMux
    port map (
            O => \N__17122\,
            I => \b2v_inst11.mult1_un82_sum_cry_7\
        );

    \I__2109\ : InMux
    port map (
            O => \N__17119\,
            I => \b2v_inst11.mult1_un96_sum_cry_6\
        );

    \I__2108\ : InMux
    port map (
            O => \N__17116\,
            I => \b2v_inst11.mult1_un96_sum_cry_7\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__17113\,
            I => \b2v_inst11.mult1_un96_sum_s_8_cascade_\
        );

    \I__2106\ : InMux
    port map (
            O => \N__17110\,
            I => \N__17107\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__17107\,
            I => \b2v_inst11.mult1_un89_sum_cry_3_s\
        );

    \I__2104\ : InMux
    port map (
            O => \N__17104\,
            I => \b2v_inst11.mult1_un89_sum_cry_2\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__17101\,
            I => \N__17098\
        );

    \I__2102\ : InMux
    port map (
            O => \N__17098\,
            I => \N__17095\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__17095\,
            I => \b2v_inst11.mult1_un89_sum_cry_4_s\
        );

    \I__2100\ : InMux
    port map (
            O => \N__17092\,
            I => \b2v_inst11.mult1_un89_sum_cry_3\
        );

    \I__2099\ : InMux
    port map (
            O => \N__17089\,
            I => \N__17086\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__17086\,
            I => \b2v_inst11.mult1_un89_sum_cry_5_s\
        );

    \I__2097\ : InMux
    port map (
            O => \N__17083\,
            I => \b2v_inst11.mult1_un89_sum_cry_4\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__17080\,
            I => \N__17077\
        );

    \I__2095\ : InMux
    port map (
            O => \N__17077\,
            I => \N__17074\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__17074\,
            I => \b2v_inst11.mult1_un89_sum_cry_6_s\
        );

    \I__2093\ : InMux
    port map (
            O => \N__17071\,
            I => \b2v_inst11.mult1_un89_sum_cry_5\
        );

    \I__2092\ : InMux
    port map (
            O => \N__17068\,
            I => \N__17065\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__17065\,
            I => \b2v_inst11.mult1_un96_sum_axb_8\
        );

    \I__2090\ : InMux
    port map (
            O => \N__17062\,
            I => \b2v_inst11.mult1_un89_sum_cry_6\
        );

    \I__2089\ : InMux
    port map (
            O => \N__17059\,
            I => \N__17056\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__17056\,
            I => \b2v_inst11.count_off_0_8\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__17053\,
            I => \N__17050\
        );

    \I__2086\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17044\
        );

    \I__2085\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17044\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__17044\,
            I => \N__17041\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__17041\,
            I => \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2\
        );

    \I__2082\ : CascadeMux
    port map (
            O => \N__17038\,
            I => \N__17035\
        );

    \I__2081\ : InMux
    port map (
            O => \N__17035\,
            I => \N__17032\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__17032\,
            I => \N__17029\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__17029\,
            I => \b2v_inst11.count_offZ0Z_8\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__17026\,
            I => \b2v_inst11.count_offZ0Z_8_cascade_\
        );

    \I__2077\ : InMux
    port map (
            O => \N__17023\,
            I => \N__17020\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__17020\,
            I => \N__17017\
        );

    \I__2075\ : Span4Mux_v
    port map (
            O => \N__17017\,
            I => \N__17014\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__17014\,
            I => \b2v_inst11.un34_clk_100khz_3\
        );

    \I__2073\ : InMux
    port map (
            O => \N__17011\,
            I => \N__17005\
        );

    \I__2072\ : InMux
    port map (
            O => \N__17010\,
            I => \N__17005\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__17005\,
            I => \b2v_inst11.count_offZ0Z_7\
        );

    \I__2070\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16998\
        );

    \I__2069\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16995\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__16998\,
            I => \b2v_inst11.count_off_1_7\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__16995\,
            I => \b2v_inst11.count_off_1_7\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__16990\,
            I => \N__16987\
        );

    \I__2065\ : InMux
    port map (
            O => \N__16987\,
            I => \N__16984\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__16984\,
            I => \N__16981\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__16981\,
            I => \b2v_inst11.un3_count_off_1_axb_7\
        );

    \I__2062\ : InMux
    port map (
            O => \N__16978\,
            I => \b2v_inst11.mult1_un96_sum_cry_2\
        );

    \I__2061\ : InMux
    port map (
            O => \N__16975\,
            I => \b2v_inst11.mult1_un96_sum_cry_3\
        );

    \I__2060\ : InMux
    port map (
            O => \N__16972\,
            I => \b2v_inst11.mult1_un96_sum_cry_4\
        );

    \I__2059\ : InMux
    port map (
            O => \N__16969\,
            I => \b2v_inst11.mult1_un96_sum_cry_5\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__16966\,
            I => \b2v_inst11.count_off_1_9_cascade_\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__16963\,
            I => \N__16959\
        );

    \I__2056\ : InMux
    port map (
            O => \N__16962\,
            I => \N__16956\
        );

    \I__2055\ : InMux
    port map (
            O => \N__16959\,
            I => \N__16953\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__16956\,
            I => \b2v_inst11.count_offZ0Z_9\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__16953\,
            I => \b2v_inst11.count_offZ0Z_9\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__16948\,
            I => \N__16945\
        );

    \I__2051\ : InMux
    port map (
            O => \N__16945\,
            I => \N__16942\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__16942\,
            I => \b2v_inst11.un3_count_off_1_axb_9\
        );

    \I__2049\ : InMux
    port map (
            O => \N__16939\,
            I => \N__16933\
        );

    \I__2048\ : InMux
    port map (
            O => \N__16938\,
            I => \N__16933\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__16933\,
            I => \b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__16930\,
            I => \N__16927\
        );

    \I__2045\ : InMux
    port map (
            O => \N__16927\,
            I => \N__16924\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__16924\,
            I => \N__16920\
        );

    \I__2043\ : InMux
    port map (
            O => \N__16923\,
            I => \N__16917\
        );

    \I__2042\ : Span4Mux_s1_h
    port map (
            O => \N__16920\,
            I => \N__16914\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__16917\,
            I => \N__16911\
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__16914\,
            I => \b2v_inst11.count_off_1_6\
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__16911\,
            I => \b2v_inst11.count_off_1_6\
        );

    \I__2038\ : InMux
    port map (
            O => \N__16906\,
            I => \N__16902\
        );

    \I__2037\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16899\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__16902\,
            I => \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__16899\,
            I => \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2\
        );

    \I__2034\ : InMux
    port map (
            O => \N__16894\,
            I => \N__16891\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__16891\,
            I => \b2v_inst11.count_off_0_15\
        );

    \I__2032\ : InMux
    port map (
            O => \N__16888\,
            I => \N__16884\
        );

    \I__2031\ : InMux
    port map (
            O => \N__16887\,
            I => \N__16881\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__16884\,
            I => \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__16881\,
            I => \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5\
        );

    \I__2028\ : InMux
    port map (
            O => \N__16876\,
            I => \N__16873\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__16873\,
            I => \b2v_inst11.count_offZ0Z_15\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__16870\,
            I => \N__16866\
        );

    \I__2025\ : InMux
    port map (
            O => \N__16869\,
            I => \N__16863\
        );

    \I__2024\ : InMux
    port map (
            O => \N__16866\,
            I => \N__16860\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__16863\,
            I => \b2v_inst11.count_offZ0Z_13\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__16860\,
            I => \b2v_inst11.count_offZ0Z_13\
        );

    \I__2021\ : InMux
    port map (
            O => \N__16855\,
            I => \N__16851\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__16854\,
            I => \N__16848\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__16851\,
            I => \N__16845\
        );

    \I__2018\ : InMux
    port map (
            O => \N__16848\,
            I => \N__16842\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__16845\,
            I => \b2v_inst11.count_offZ0Z_14\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__16842\,
            I => \b2v_inst11.count_offZ0Z_14\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__16837\,
            I => \b2v_inst11.count_offZ0Z_15_cascade_\
        );

    \I__2014\ : InMux
    port map (
            O => \N__16834\,
            I => \N__16831\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__16831\,
            I => \N__16828\
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__16828\,
            I => \b2v_inst11.un34_clk_100khz_11\
        );

    \I__2011\ : InMux
    port map (
            O => \N__16825\,
            I => \N__16819\
        );

    \I__2010\ : InMux
    port map (
            O => \N__16824\,
            I => \N__16819\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__16819\,
            I => \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5\
        );

    \I__2008\ : InMux
    port map (
            O => \N__16816\,
            I => \N__16813\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__16813\,
            I => \b2v_inst11.un34_clk_100khz_12\
        );

    \I__2006\ : CascadeMux
    port map (
            O => \N__16810\,
            I => \b2v_inst11.un34_clk_100khz_4_cascade_\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__16807\,
            I => \N__16804\
        );

    \I__2004\ : InMux
    port map (
            O => \N__16804\,
            I => \N__16801\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__16801\,
            I => \b2v_inst11.count_off_0_12\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__16798\,
            I => \N__16795\
        );

    \I__2001\ : InMux
    port map (
            O => \N__16795\,
            I => \N__16789\
        );

    \I__2000\ : InMux
    port map (
            O => \N__16794\,
            I => \N__16789\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__16789\,
            I => \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__16786\,
            I => \N__16783\
        );

    \I__1997\ : InMux
    port map (
            O => \N__16783\,
            I => \N__16780\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__16780\,
            I => \b2v_inst11.count_offZ0Z_12\
        );

    \I__1995\ : InMux
    port map (
            O => \N__16777\,
            I => \N__16774\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__16774\,
            I => \b2v_inst11.count_off_1_11\
        );

    \I__1993\ : InMux
    port map (
            O => \N__16771\,
            I => \N__16765\
        );

    \I__1992\ : InMux
    port map (
            O => \N__16770\,
            I => \N__16765\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__16765\,
            I => \b2v_inst11.count_offZ0Z_11\
        );

    \I__1990\ : CascadeMux
    port map (
            O => \N__16762\,
            I => \b2v_inst11.count_offZ0Z_12_cascade_\
        );

    \I__1989\ : InMux
    port map (
            O => \N__16759\,
            I => \N__16756\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__16756\,
            I => \b2v_inst11.un34_clk_100khz_5\
        );

    \I__1987\ : InMux
    port map (
            O => \N__16753\,
            I => \N__16749\
        );

    \I__1986\ : InMux
    port map (
            O => \N__16752\,
            I => \N__16746\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__16749\,
            I => \N__16743\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__16746\,
            I => \N__16740\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__16743\,
            I => \b2v_inst11.count_offZ0Z_6\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__16740\,
            I => \b2v_inst11.count_offZ0Z_6\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__16735\,
            I => \N__16732\
        );

    \I__1980\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16726\
        );

    \I__1979\ : InMux
    port map (
            O => \N__16731\,
            I => \N__16726\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__16726\,
            I => \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2\
        );

    \I__1977\ : InMux
    port map (
            O => \N__16723\,
            I => \N__16720\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__16720\,
            I => \b2v_inst11.count_off_1_9\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__16717\,
            I => \N__16714\
        );

    \I__1974\ : InMux
    port map (
            O => \N__16714\,
            I => \N__16709\
        );

    \I__1973\ : InMux
    port map (
            O => \N__16713\,
            I => \N__16704\
        );

    \I__1972\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16704\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__16709\,
            I => \N__16701\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__16704\,
            I => \b2v_inst11.count_clkZ0Z_9\
        );

    \I__1969\ : Odrv4
    port map (
            O => \N__16701\,
            I => \b2v_inst11.count_clkZ0Z_9\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__16696\,
            I => \N__16693\
        );

    \I__1967\ : InMux
    port map (
            O => \N__16693\,
            I => \N__16687\
        );

    \I__1966\ : InMux
    port map (
            O => \N__16692\,
            I => \N__16680\
        );

    \I__1965\ : InMux
    port map (
            O => \N__16691\,
            I => \N__16680\
        );

    \I__1964\ : InMux
    port map (
            O => \N__16690\,
            I => \N__16680\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__16687\,
            I => \N__16677\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__16680\,
            I => \b2v_inst11.count_clkZ0Z_1\
        );

    \I__1961\ : Odrv4
    port map (
            O => \N__16677\,
            I => \b2v_inst11.count_clkZ0Z_1\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__16672\,
            I => \N__16669\
        );

    \I__1959\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16666\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__16666\,
            I => \b2v_inst11.count_clk_RNIZ0Z_5\
        );

    \I__1957\ : InMux
    port map (
            O => \N__16663\,
            I => \N__16657\
        );

    \I__1956\ : InMux
    port map (
            O => \N__16662\,
            I => \N__16657\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__16657\,
            I => \N__16654\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__16654\,
            I => \b2v_inst11.N_172\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__16651\,
            I => \N__16648\
        );

    \I__1952\ : InMux
    port map (
            O => \N__16648\,
            I => \N__16645\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__16645\,
            I => \N__16642\
        );

    \I__1950\ : Span4Mux_v
    port map (
            O => \N__16642\,
            I => \N__16638\
        );

    \I__1949\ : InMux
    port map (
            O => \N__16641\,
            I => \N__16635\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__16638\,
            I => \b2v_inst11.N_421\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__16635\,
            I => \b2v_inst11.N_421\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__16630\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\
        );

    \I__1945\ : InMux
    port map (
            O => \N__16627\,
            I => \N__16624\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__16624\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_i_1\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__16621\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_0_cascade_\
        );

    \I__1942\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16614\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__16617\,
            I => \N__16607\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__16614\,
            I => \N__16596\
        );

    \I__1939\ : InMux
    port map (
            O => \N__16613\,
            I => \N__16582\
        );

    \I__1938\ : InMux
    port map (
            O => \N__16612\,
            I => \N__16582\
        );

    \I__1937\ : InMux
    port map (
            O => \N__16611\,
            I => \N__16582\
        );

    \I__1936\ : InMux
    port map (
            O => \N__16610\,
            I => \N__16582\
        );

    \I__1935\ : InMux
    port map (
            O => \N__16607\,
            I => \N__16582\
        );

    \I__1934\ : InMux
    port map (
            O => \N__16606\,
            I => \N__16573\
        );

    \I__1933\ : InMux
    port map (
            O => \N__16605\,
            I => \N__16573\
        );

    \I__1932\ : InMux
    port map (
            O => \N__16604\,
            I => \N__16573\
        );

    \I__1931\ : InMux
    port map (
            O => \N__16603\,
            I => \N__16573\
        );

    \I__1930\ : InMux
    port map (
            O => \N__16602\,
            I => \N__16566\
        );

    \I__1929\ : InMux
    port map (
            O => \N__16601\,
            I => \N__16566\
        );

    \I__1928\ : InMux
    port map (
            O => \N__16600\,
            I => \N__16566\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__16599\,
            I => \N__16561\
        );

    \I__1926\ : Span4Mux_v
    port map (
            O => \N__16596\,
            I => \N__16558\
        );

    \I__1925\ : InMux
    port map (
            O => \N__16595\,
            I => \N__16551\
        );

    \I__1924\ : InMux
    port map (
            O => \N__16594\,
            I => \N__16551\
        );

    \I__1923\ : InMux
    port map (
            O => \N__16593\,
            I => \N__16551\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__16582\,
            I => \N__16544\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__16573\,
            I => \N__16544\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__16566\,
            I => \N__16544\
        );

    \I__1919\ : InMux
    port map (
            O => \N__16565\,
            I => \N__16535\
        );

    \I__1918\ : InMux
    port map (
            O => \N__16564\,
            I => \N__16535\
        );

    \I__1917\ : InMux
    port map (
            O => \N__16561\,
            I => \N__16535\
        );

    \I__1916\ : Span4Mux_s1_h
    port map (
            O => \N__16558\,
            I => \N__16530\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__16551\,
            I => \N__16530\
        );

    \I__1914\ : Span4Mux_s2_h
    port map (
            O => \N__16544\,
            I => \N__16527\
        );

    \I__1913\ : InMux
    port map (
            O => \N__16543\,
            I => \N__16522\
        );

    \I__1912\ : InMux
    port map (
            O => \N__16542\,
            I => \N__16522\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__16535\,
            I => \b2v_inst11.func_state_RNICC5V2_0_1\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__16530\,
            I => \b2v_inst11.func_state_RNICC5V2_0_1\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__16527\,
            I => \b2v_inst11.func_state_RNICC5V2_0_1\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__16522\,
            I => \b2v_inst11.func_state_RNICC5V2_0_1\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__16513\,
            I => \b2v_inst11.count_off_1_11_cascade_\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__16510\,
            I => \N__16507\
        );

    \I__1905\ : InMux
    port map (
            O => \N__16507\,
            I => \N__16504\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__16504\,
            I => \b2v_inst11.un3_count_off_1_axb_11\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__16501\,
            I => \b2v_inst11.count_clk_RNIZ0Z_3_cascade_\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__16498\,
            I => \N__16495\
        );

    \I__1901\ : InMux
    port map (
            O => \N__16495\,
            I => \N__16492\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__16492\,
            I => \b2v_inst11.count_clk_en_0\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__16489\,
            I => \N__16485\
        );

    \I__1898\ : InMux
    port map (
            O => \N__16488\,
            I => \N__16482\
        );

    \I__1897\ : InMux
    port map (
            O => \N__16485\,
            I => \N__16479\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__16482\,
            I => \N__16474\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__16479\,
            I => \N__16474\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__16474\,
            I => \b2v_inst11.count_clkZ0Z_12\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__16471\,
            I => \N__16468\
        );

    \I__1892\ : InMux
    port map (
            O => \N__16468\,
            I => \N__16462\
        );

    \I__1891\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16462\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__16462\,
            I => \N__16459\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__16459\,
            I => \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BAZ0\
        );

    \I__1888\ : InMux
    port map (
            O => \N__16456\,
            I => \N__16453\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__16453\,
            I => \b2v_inst11.count_clk_0_12\
        );

    \I__1886\ : InMux
    port map (
            O => \N__16450\,
            I => \N__16447\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__16447\,
            I => \N__16444\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__16444\,
            I => \b2v_inst11.count_clk_RNI_0Z0Z_0\
        );

    \I__1883\ : InMux
    port map (
            O => \N__16441\,
            I => \N__16432\
        );

    \I__1882\ : InMux
    port map (
            O => \N__16440\,
            I => \N__16432\
        );

    \I__1881\ : InMux
    port map (
            O => \N__16439\,
            I => \N__16432\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__16432\,
            I => \N__16427\
        );

    \I__1879\ : InMux
    port map (
            O => \N__16431\,
            I => \N__16424\
        );

    \I__1878\ : InMux
    port map (
            O => \N__16430\,
            I => \N__16421\
        );

    \I__1877\ : Odrv12
    port map (
            O => \N__16427\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__16424\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__16421\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__1874\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16411\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__16411\,
            I => \b2v_inst11.count_clk_0_1\
        );

    \I__1872\ : CascadeMux
    port map (
            O => \N__16408\,
            I => \b2v_inst11.count_clk_RNIZ0Z_0_cascade_\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__16405\,
            I => \b2v_inst11.count_clkZ0Z_1_cascade_\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__16402\,
            I => \N__16399\
        );

    \I__1869\ : InMux
    port map (
            O => \N__16399\,
            I => \N__16394\
        );

    \I__1868\ : InMux
    port map (
            O => \N__16398\,
            I => \N__16391\
        );

    \I__1867\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16388\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__16394\,
            I => \N__16385\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__16391\,
            I => \b2v_inst11.count_clkZ0Z_5\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__16388\,
            I => \b2v_inst11.count_clkZ0Z_5\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__16385\,
            I => \b2v_inst11.count_clkZ0Z_5\
        );

    \I__1862\ : InMux
    port map (
            O => \N__16378\,
            I => \N__16372\
        );

    \I__1861\ : InMux
    port map (
            O => \N__16377\,
            I => \N__16372\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__16372\,
            I => \b2v_inst11.N_187\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__16369\,
            I => \b2v_inst11.count_clk_en_cascade_\
        );

    \I__1858\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16360\
        );

    \I__1857\ : InMux
    port map (
            O => \N__16365\,
            I => \N__16360\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__16360\,
            I => \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5\
        );

    \I__1855\ : InMux
    port map (
            O => \N__16357\,
            I => \N__16354\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__16354\,
            I => \b2v_inst11.count_clk_0_2\
        );

    \I__1853\ : CascadeMux
    port map (
            O => \N__16351\,
            I => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_\
        );

    \I__1852\ : InMux
    port map (
            O => \N__16348\,
            I => \N__16345\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__16345\,
            I => \b2v_inst11.N_373\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__16342\,
            I => \b2v_inst11.N_373_cascade_\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__16339\,
            I => \N__16336\
        );

    \I__1848\ : InMux
    port map (
            O => \N__16336\,
            I => \N__16331\
        );

    \I__1847\ : InMux
    port map (
            O => \N__16335\,
            I => \N__16326\
        );

    \I__1846\ : InMux
    port map (
            O => \N__16334\,
            I => \N__16326\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__16331\,
            I => \N__16323\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__16326\,
            I => \b2v_inst11.count_clkZ0Z_8\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__16323\,
            I => \b2v_inst11.count_clkZ0Z_8\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__16318\,
            I => \N__16315\
        );

    \I__1841\ : InMux
    port map (
            O => \N__16315\,
            I => \N__16310\
        );

    \I__1840\ : InMux
    port map (
            O => \N__16314\,
            I => \N__16305\
        );

    \I__1839\ : InMux
    port map (
            O => \N__16313\,
            I => \N__16305\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__16310\,
            I => \N__16302\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__16305\,
            I => \b2v_inst11.count_clkZ0Z_6\
        );

    \I__1836\ : Odrv4
    port map (
            O => \N__16302\,
            I => \b2v_inst11.count_clkZ0Z_6\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__16297\,
            I => \N__16293\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__16296\,
            I => \N__16290\
        );

    \I__1833\ : InMux
    port map (
            O => \N__16293\,
            I => \N__16286\
        );

    \I__1832\ : InMux
    port map (
            O => \N__16290\,
            I => \N__16283\
        );

    \I__1831\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16280\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__16286\,
            I => \N__16277\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__16283\,
            I => \b2v_inst11.count_clkZ0Z_4\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__16280\,
            I => \b2v_inst11.count_clkZ0Z_4\
        );

    \I__1827\ : Odrv4
    port map (
            O => \N__16277\,
            I => \b2v_inst11.count_clkZ0Z_4\
        );

    \I__1826\ : InMux
    port map (
            O => \N__16270\,
            I => \N__16265\
        );

    \I__1825\ : InMux
    port map (
            O => \N__16269\,
            I => \N__16260\
        );

    \I__1824\ : InMux
    port map (
            O => \N__16268\,
            I => \N__16260\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__16265\,
            I => \b2v_inst11.count_clkZ0Z_2\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__16260\,
            I => \b2v_inst11.count_clkZ0Z_2\
        );

    \I__1821\ : InMux
    port map (
            O => \N__16255\,
            I => \N__16248\
        );

    \I__1820\ : InMux
    port map (
            O => \N__16254\,
            I => \N__16248\
        );

    \I__1819\ : InMux
    port map (
            O => \N__16253\,
            I => \N__16245\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__16248\,
            I => \b2v_inst11.count_clkZ0Z_3\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__16245\,
            I => \b2v_inst11.count_clkZ0Z_3\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__16240\,
            I => \b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__16237\,
            I => \N__16234\
        );

    \I__1814\ : InMux
    port map (
            O => \N__16234\,
            I => \N__16228\
        );

    \I__1813\ : InMux
    port map (
            O => \N__16233\,
            I => \N__16221\
        );

    \I__1812\ : InMux
    port map (
            O => \N__16232\,
            I => \N__16221\
        );

    \I__1811\ : InMux
    port map (
            O => \N__16231\,
            I => \N__16221\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__16228\,
            I => \N__16218\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__16221\,
            I => \b2v_inst11.count_clkZ0Z_7\
        );

    \I__1808\ : Odrv4
    port map (
            O => \N__16218\,
            I => \b2v_inst11.count_clkZ0Z_7\
        );

    \I__1807\ : InMux
    port map (
            O => \N__16213\,
            I => \N__16210\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__16210\,
            I => \b2v_inst11.count_clk_0_0\
        );

    \I__1805\ : InMux
    port map (
            O => \N__16207\,
            I => \N__16204\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__16204\,
            I => \b2v_inst11.count_clk_0_10\
        );

    \I__1803\ : InMux
    port map (
            O => \N__16201\,
            I => \N__16195\
        );

    \I__1802\ : InMux
    port map (
            O => \N__16200\,
            I => \N__16195\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__16195\,
            I => \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__16192\,
            I => \N__16189\
        );

    \I__1799\ : InMux
    port map (
            O => \N__16189\,
            I => \N__16186\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__16186\,
            I => \b2v_inst11.count_clkZ0Z_10\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__16183\,
            I => \N__16179\
        );

    \I__1796\ : InMux
    port map (
            O => \N__16182\,
            I => \N__16176\
        );

    \I__1795\ : InMux
    port map (
            O => \N__16179\,
            I => \N__16173\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__16176\,
            I => \b2v_inst11.count_clkZ0Z_11\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__16173\,
            I => \b2v_inst11.count_clkZ0Z_11\
        );

    \I__1792\ : CascadeMux
    port map (
            O => \N__16168\,
            I => \b2v_inst11.count_clkZ0Z_10_cascade_\
        );

    \I__1791\ : InMux
    port map (
            O => \N__16165\,
            I => \N__16161\
        );

    \I__1790\ : InMux
    port map (
            O => \N__16164\,
            I => \N__16158\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__16161\,
            I => \N__16155\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__16158\,
            I => \b2v_inst11.count_clkZ0Z_15\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__16155\,
            I => \b2v_inst11.count_clkZ0Z_15\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__16150\,
            I => \b2v_inst11.un2_count_clk_17_0_o2_1_4_cascade_\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__16147\,
            I => \N__16143\
        );

    \I__1784\ : InMux
    port map (
            O => \N__16146\,
            I => \N__16140\
        );

    \I__1783\ : InMux
    port map (
            O => \N__16143\,
            I => \N__16137\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__16140\,
            I => \b2v_inst11.count_clkZ0Z_14\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__16137\,
            I => \b2v_inst11.count_clkZ0Z_14\
        );

    \I__1780\ : InMux
    port map (
            O => \N__16132\,
            I => \N__16129\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__16129\,
            I => \b2v_inst11.count_clk_0_13\
        );

    \I__1778\ : InMux
    port map (
            O => \N__16126\,
            I => \N__16120\
        );

    \I__1777\ : InMux
    port map (
            O => \N__16125\,
            I => \N__16120\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__16120\,
            I => \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CAZ0\
        );

    \I__1775\ : CascadeMux
    port map (
            O => \N__16117\,
            I => \N__16113\
        );

    \I__1774\ : InMux
    port map (
            O => \N__16116\,
            I => \N__16110\
        );

    \I__1773\ : InMux
    port map (
            O => \N__16113\,
            I => \N__16107\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__16110\,
            I => \b2v_inst11.count_clkZ0Z_13\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__16107\,
            I => \b2v_inst11.count_clkZ0Z_13\
        );

    \I__1770\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16096\
        );

    \I__1769\ : InMux
    port map (
            O => \N__16101\,
            I => \N__16096\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__16096\,
            I => \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DAZ0\
        );

    \I__1767\ : InMux
    port map (
            O => \N__16093\,
            I => \N__16090\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__16090\,
            I => \b2v_inst11.count_clk_0_14\
        );

    \I__1765\ : InMux
    port map (
            O => \N__16087\,
            I => \N__16083\
        );

    \I__1764\ : InMux
    port map (
            O => \N__16086\,
            I => \N__16080\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__16083\,
            I => \b2v_inst200.countZ0Z_14\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__16080\,
            I => \b2v_inst200.countZ0Z_14\
        );

    \I__1761\ : InMux
    port map (
            O => \N__16075\,
            I => \N__16069\
        );

    \I__1760\ : InMux
    port map (
            O => \N__16074\,
            I => \N__16069\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__16069\,
            I => \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59\
        );

    \I__1758\ : InMux
    port map (
            O => \N__16066\,
            I => \b2v_inst200.un2_count_1_cry_13\
        );

    \I__1757\ : InMux
    port map (
            O => \N__16063\,
            I => \N__16059\
        );

    \I__1756\ : InMux
    port map (
            O => \N__16062\,
            I => \N__16056\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__16059\,
            I => \b2v_inst200.countZ0Z_15\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__16056\,
            I => \b2v_inst200.countZ0Z_15\
        );

    \I__1753\ : InMux
    port map (
            O => \N__16051\,
            I => \N__16048\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__16048\,
            I => \N__16044\
        );

    \I__1751\ : InMux
    port map (
            O => \N__16047\,
            I => \N__16041\
        );

    \I__1750\ : Odrv12
    port map (
            O => \N__16044\,
            I => \b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__16041\,
            I => \b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69\
        );

    \I__1748\ : InMux
    port map (
            O => \N__16036\,
            I => \b2v_inst200.un2_count_1_cry_14\
        );

    \I__1747\ : InMux
    port map (
            O => \N__16033\,
            I => \N__16030\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__16030\,
            I => \N__16027\
        );

    \I__1745\ : Span4Mux_v
    port map (
            O => \N__16027\,
            I => \N__16023\
        );

    \I__1744\ : InMux
    port map (
            O => \N__16026\,
            I => \N__16020\
        );

    \I__1743\ : Odrv4
    port map (
            O => \N__16023\,
            I => \b2v_inst200.countZ0Z_16\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__16020\,
            I => \b2v_inst200.countZ0Z_16\
        );

    \I__1741\ : InMux
    port map (
            O => \N__16015\,
            I => \N__16009\
        );

    \I__1740\ : InMux
    port map (
            O => \N__16014\,
            I => \N__16009\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__16009\,
            I => \N__16006\
        );

    \I__1738\ : Odrv4
    port map (
            O => \N__16006\,
            I => \b2v_inst200.count_1_16\
        );

    \I__1737\ : InMux
    port map (
            O => \N__16003\,
            I => \bfn_2_8_0_\
        );

    \I__1736\ : InMux
    port map (
            O => \N__16000\,
            I => \N__15997\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__15997\,
            I => \N__15993\
        );

    \I__1734\ : InMux
    port map (
            O => \N__15996\,
            I => \N__15990\
        );

    \I__1733\ : Odrv12
    port map (
            O => \N__15993\,
            I => \b2v_inst200.countZ0Z_17\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__15990\,
            I => \b2v_inst200.countZ0Z_17\
        );

    \I__1731\ : InMux
    port map (
            O => \N__15985\,
            I => \b2v_inst200.un2_count_1_cry_16\
        );

    \I__1730\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15976\
        );

    \I__1729\ : InMux
    port map (
            O => \N__15981\,
            I => \N__15976\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__15976\,
            I => \N__15973\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__15973\,
            I => \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\
        );

    \I__1726\ : InMux
    port map (
            O => \N__15970\,
            I => \N__15964\
        );

    \I__1725\ : InMux
    port map (
            O => \N__15969\,
            I => \N__15964\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__15964\,
            I => \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AAZ0\
        );

    \I__1723\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15958\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__15958\,
            I => \b2v_inst11.count_clk_0_11\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__15955\,
            I => \b2v_inst11.count_clkZ0Z_0_cascade_\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__15952\,
            I => \N__15949\
        );

    \I__1719\ : InMux
    port map (
            O => \N__15949\,
            I => \N__15945\
        );

    \I__1718\ : InMux
    port map (
            O => \N__15948\,
            I => \N__15942\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__15945\,
            I => \b2v_inst200.countZ0Z_6\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__15942\,
            I => \b2v_inst200.countZ0Z_6\
        );

    \I__1715\ : InMux
    port map (
            O => \N__15937\,
            I => \N__15933\
        );

    \I__1714\ : InMux
    port map (
            O => \N__15936\,
            I => \N__15930\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__15933\,
            I => \b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__15930\,
            I => \b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0\
        );

    \I__1711\ : InMux
    port map (
            O => \N__15925\,
            I => \b2v_inst200.un2_count_1_cry_5\
        );

    \I__1710\ : InMux
    port map (
            O => \N__15922\,
            I => \N__15918\
        );

    \I__1709\ : InMux
    port map (
            O => \N__15921\,
            I => \N__15915\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__15918\,
            I => \b2v_inst200.countZ0Z_7\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__15915\,
            I => \b2v_inst200.countZ0Z_7\
        );

    \I__1706\ : InMux
    port map (
            O => \N__15910\,
            I => \N__15907\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__15907\,
            I => \N__15903\
        );

    \I__1704\ : InMux
    port map (
            O => \N__15906\,
            I => \N__15900\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__15903\,
            I => \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__15900\,
            I => \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\
        );

    \I__1701\ : InMux
    port map (
            O => \N__15895\,
            I => \b2v_inst200.un2_count_1_cry_6\
        );

    \I__1700\ : InMux
    port map (
            O => \N__15892\,
            I => \N__15888\
        );

    \I__1699\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15885\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__15888\,
            I => \b2v_inst200.countZ0Z_8\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__15885\,
            I => \b2v_inst200.countZ0Z_8\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__15880\,
            I => \N__15877\
        );

    \I__1695\ : InMux
    port map (
            O => \N__15877\,
            I => \N__15871\
        );

    \I__1694\ : InMux
    port map (
            O => \N__15876\,
            I => \N__15871\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__15871\,
            I => \b2v_inst200.un2_count_1_cry_7_c_RNIP33EZ0\
        );

    \I__1692\ : InMux
    port map (
            O => \N__15868\,
            I => \bfn_2_7_0_\
        );

    \I__1691\ : InMux
    port map (
            O => \N__15865\,
            I => \N__15862\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__15862\,
            I => \b2v_inst200.countZ0Z_9\
        );

    \I__1689\ : InMux
    port map (
            O => \N__15859\,
            I => \N__15853\
        );

    \I__1688\ : InMux
    port map (
            O => \N__15858\,
            I => \N__15853\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__15853\,
            I => \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0\
        );

    \I__1686\ : InMux
    port map (
            O => \N__15850\,
            I => \b2v_inst200.un2_count_1_cry_8\
        );

    \I__1685\ : InMux
    port map (
            O => \N__15847\,
            I => \N__15844\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__15844\,
            I => \N__15840\
        );

    \I__1683\ : InMux
    port map (
            O => \N__15843\,
            I => \N__15837\
        );

    \I__1682\ : Odrv4
    port map (
            O => \N__15840\,
            I => \b2v_inst200.countZ0Z_10\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__15837\,
            I => \b2v_inst200.countZ0Z_10\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__15832\,
            I => \N__15829\
        );

    \I__1679\ : InMux
    port map (
            O => \N__15829\,
            I => \N__15823\
        );

    \I__1678\ : InMux
    port map (
            O => \N__15828\,
            I => \N__15823\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__15823\,
            I => \N__15820\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__15820\,
            I => \b2v_inst200.un2_count_1_cry_9_c_RNIR75EZ0\
        );

    \I__1675\ : InMux
    port map (
            O => \N__15817\,
            I => \b2v_inst200.un2_count_1_cry_9\
        );

    \I__1674\ : InMux
    port map (
            O => \N__15814\,
            I => \N__15810\
        );

    \I__1673\ : CascadeMux
    port map (
            O => \N__15813\,
            I => \N__15807\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__15810\,
            I => \N__15804\
        );

    \I__1671\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15801\
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__15804\,
            I => \b2v_inst200.countZ0Z_11\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__15801\,
            I => \b2v_inst200.countZ0Z_11\
        );

    \I__1668\ : InMux
    port map (
            O => \N__15796\,
            I => \N__15790\
        );

    \I__1667\ : InMux
    port map (
            O => \N__15795\,
            I => \N__15790\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__15790\,
            I => \N__15787\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__15787\,
            I => \b2v_inst200.un2_count_1_cry_10_c_RNI3AZ0Z29\
        );

    \I__1664\ : InMux
    port map (
            O => \N__15784\,
            I => \b2v_inst200.un2_count_1_cry_10\
        );

    \I__1663\ : InMux
    port map (
            O => \N__15781\,
            I => \N__15777\
        );

    \I__1662\ : InMux
    port map (
            O => \N__15780\,
            I => \N__15774\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__15777\,
            I => \b2v_inst200.countZ0Z_12\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__15774\,
            I => \b2v_inst200.countZ0Z_12\
        );

    \I__1659\ : InMux
    port map (
            O => \N__15769\,
            I => \N__15763\
        );

    \I__1658\ : InMux
    port map (
            O => \N__15768\,
            I => \N__15763\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__15763\,
            I => \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39\
        );

    \I__1656\ : InMux
    port map (
            O => \N__15760\,
            I => \b2v_inst200.un2_count_1_cry_11\
        );

    \I__1655\ : InMux
    port map (
            O => \N__15757\,
            I => \N__15753\
        );

    \I__1654\ : InMux
    port map (
            O => \N__15756\,
            I => \N__15750\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__15753\,
            I => \b2v_inst200.countZ0Z_13\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__15750\,
            I => \b2v_inst200.countZ0Z_13\
        );

    \I__1651\ : InMux
    port map (
            O => \N__15745\,
            I => \N__15739\
        );

    \I__1650\ : InMux
    port map (
            O => \N__15744\,
            I => \N__15739\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__15739\,
            I => \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49\
        );

    \I__1648\ : InMux
    port map (
            O => \N__15736\,
            I => \b2v_inst200.un2_count_1_cry_12\
        );

    \I__1647\ : InMux
    port map (
            O => \N__15733\,
            I => \N__15730\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__15730\,
            I => \b2v_inst200.count_2_1\
        );

    \I__1645\ : InMux
    port map (
            O => \N__15727\,
            I => \N__15724\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__15724\,
            I => \b2v_inst200.count_2_2\
        );

    \I__1643\ : InMux
    port map (
            O => \N__15721\,
            I => \N__15701\
        );

    \I__1642\ : InMux
    port map (
            O => \N__15720\,
            I => \N__15696\
        );

    \I__1641\ : InMux
    port map (
            O => \N__15719\,
            I => \N__15696\
        );

    \I__1640\ : InMux
    port map (
            O => \N__15718\,
            I => \N__15689\
        );

    \I__1639\ : InMux
    port map (
            O => \N__15717\,
            I => \N__15689\
        );

    \I__1638\ : InMux
    port map (
            O => \N__15716\,
            I => \N__15689\
        );

    \I__1637\ : InMux
    port map (
            O => \N__15715\,
            I => \N__15680\
        );

    \I__1636\ : InMux
    port map (
            O => \N__15714\,
            I => \N__15680\
        );

    \I__1635\ : InMux
    port map (
            O => \N__15713\,
            I => \N__15680\
        );

    \I__1634\ : InMux
    port map (
            O => \N__15712\,
            I => \N__15680\
        );

    \I__1633\ : InMux
    port map (
            O => \N__15711\,
            I => \N__15671\
        );

    \I__1632\ : InMux
    port map (
            O => \N__15710\,
            I => \N__15671\
        );

    \I__1631\ : InMux
    port map (
            O => \N__15709\,
            I => \N__15671\
        );

    \I__1630\ : InMux
    port map (
            O => \N__15708\,
            I => \N__15671\
        );

    \I__1629\ : InMux
    port map (
            O => \N__15707\,
            I => \N__15662\
        );

    \I__1628\ : InMux
    port map (
            O => \N__15706\,
            I => \N__15662\
        );

    \I__1627\ : InMux
    port map (
            O => \N__15705\,
            I => \N__15662\
        );

    \I__1626\ : InMux
    port map (
            O => \N__15704\,
            I => \N__15662\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__15701\,
            I => \N__15653\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__15696\,
            I => \N__15650\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__15689\,
            I => \N__15647\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__15680\,
            I => \N__15644\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__15671\,
            I => \N__15641\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__15662\,
            I => \N__15638\
        );

    \I__1619\ : CEMux
    port map (
            O => \N__15661\,
            I => \N__15613\
        );

    \I__1618\ : CEMux
    port map (
            O => \N__15660\,
            I => \N__15613\
        );

    \I__1617\ : CEMux
    port map (
            O => \N__15659\,
            I => \N__15613\
        );

    \I__1616\ : CEMux
    port map (
            O => \N__15658\,
            I => \N__15613\
        );

    \I__1615\ : CEMux
    port map (
            O => \N__15657\,
            I => \N__15613\
        );

    \I__1614\ : CEMux
    port map (
            O => \N__15656\,
            I => \N__15613\
        );

    \I__1613\ : Glb2LocalMux
    port map (
            O => \N__15653\,
            I => \N__15613\
        );

    \I__1612\ : Glb2LocalMux
    port map (
            O => \N__15650\,
            I => \N__15613\
        );

    \I__1611\ : Glb2LocalMux
    port map (
            O => \N__15647\,
            I => \N__15613\
        );

    \I__1610\ : Glb2LocalMux
    port map (
            O => \N__15644\,
            I => \N__15613\
        );

    \I__1609\ : Glb2LocalMux
    port map (
            O => \N__15641\,
            I => \N__15613\
        );

    \I__1608\ : Glb2LocalMux
    port map (
            O => \N__15638\,
            I => \N__15613\
        );

    \I__1607\ : GlobalMux
    port map (
            O => \N__15613\,
            I => \N__15610\
        );

    \I__1606\ : gio2CtrlBuf
    port map (
            O => \N__15610\,
            I => \b2v_inst200.count_en_g\
        );

    \I__1605\ : InMux
    port map (
            O => \N__15607\,
            I => \N__15603\
        );

    \I__1604\ : InMux
    port map (
            O => \N__15606\,
            I => \N__15600\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__15603\,
            I => \b2v_inst200.countZ0Z_0\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__15600\,
            I => \b2v_inst200.countZ0Z_0\
        );

    \I__1601\ : InMux
    port map (
            O => \N__15595\,
            I => \N__15592\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__15592\,
            I => \b2v_inst200.count_1_0\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__15589\,
            I => \N__15586\
        );

    \I__1598\ : InMux
    port map (
            O => \N__15586\,
            I => \N__15582\
        );

    \I__1597\ : InMux
    port map (
            O => \N__15585\,
            I => \N__15579\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__15582\,
            I => \b2v_inst200.countZ0Z_1\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__15579\,
            I => \b2v_inst200.countZ0Z_1\
        );

    \I__1594\ : InMux
    port map (
            O => \N__15574\,
            I => \N__15568\
        );

    \I__1593\ : InMux
    port map (
            O => \N__15573\,
            I => \N__15568\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__15568\,
            I => \b2v_inst200.count_RNIC03N_5Z0Z_0\
        );

    \I__1591\ : InMux
    port map (
            O => \N__15565\,
            I => \b2v_inst200.un2_count_1_cry_1_cy\
        );

    \I__1590\ : InMux
    port map (
            O => \N__15562\,
            I => \N__15558\
        );

    \I__1589\ : InMux
    port map (
            O => \N__15561\,
            I => \N__15555\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__15558\,
            I => \b2v_inst200.countZ0Z_2\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__15555\,
            I => \b2v_inst200.countZ0Z_2\
        );

    \I__1586\ : InMux
    port map (
            O => \N__15550\,
            I => \N__15546\
        );

    \I__1585\ : InMux
    port map (
            O => \N__15549\,
            I => \N__15543\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__15546\,
            I => \N__15540\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__15543\,
            I => \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__15540\,
            I => \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\
        );

    \I__1581\ : InMux
    port map (
            O => \N__15535\,
            I => \b2v_inst200.un2_count_1_cry_1\
        );

    \I__1580\ : InMux
    port map (
            O => \N__15532\,
            I => \N__15528\
        );

    \I__1579\ : InMux
    port map (
            O => \N__15531\,
            I => \N__15525\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__15528\,
            I => \b2v_inst200.countZ0Z_3\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__15525\,
            I => \b2v_inst200.countZ0Z_3\
        );

    \I__1576\ : InMux
    port map (
            O => \N__15520\,
            I => \N__15514\
        );

    \I__1575\ : InMux
    port map (
            O => \N__15519\,
            I => \N__15514\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__15514\,
            I => \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0\
        );

    \I__1573\ : InMux
    port map (
            O => \N__15511\,
            I => \b2v_inst200.un2_count_1_cry_2\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__15508\,
            I => \N__15505\
        );

    \I__1571\ : InMux
    port map (
            O => \N__15505\,
            I => \N__15501\
        );

    \I__1570\ : InMux
    port map (
            O => \N__15504\,
            I => \N__15498\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__15501\,
            I => \b2v_inst200.countZ0Z_4\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__15498\,
            I => \b2v_inst200.countZ0Z_4\
        );

    \I__1567\ : InMux
    port map (
            O => \N__15493\,
            I => \N__15487\
        );

    \I__1566\ : InMux
    port map (
            O => \N__15492\,
            I => \N__15487\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__15487\,
            I => \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\
        );

    \I__1564\ : InMux
    port map (
            O => \N__15484\,
            I => \b2v_inst200.un2_count_1_cry_3\
        );

    \I__1563\ : InMux
    port map (
            O => \N__15481\,
            I => \N__15477\
        );

    \I__1562\ : InMux
    port map (
            O => \N__15480\,
            I => \N__15474\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__15477\,
            I => \b2v_inst200.countZ0Z_5\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__15474\,
            I => \b2v_inst200.countZ0Z_5\
        );

    \I__1559\ : InMux
    port map (
            O => \N__15469\,
            I => \N__15463\
        );

    \I__1558\ : InMux
    port map (
            O => \N__15468\,
            I => \N__15463\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__15463\,
            I => \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\
        );

    \I__1556\ : InMux
    port map (
            O => \N__15460\,
            I => \b2v_inst200.un2_count_1_cry_4\
        );

    \I__1555\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15454\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__15454\,
            I => \N__15451\
        );

    \I__1553\ : Span4Mux_v
    port map (
            O => \N__15451\,
            I => \N__15448\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__15448\,
            I => \b2v_inst200.count_2_15\
        );

    \I__1551\ : InMux
    port map (
            O => \N__15445\,
            I => \N__15442\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__15442\,
            I => \N__15439\
        );

    \I__1549\ : Span4Mux_s1_h
    port map (
            O => \N__15439\,
            I => \N__15436\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__15436\,
            I => \b2v_inst200.count_2_7\
        );

    \I__1547\ : InMux
    port map (
            O => \N__15433\,
            I => \N__15430\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__15430\,
            I => \b2v_inst200.un25_clk_100khz_11\
        );

    \I__1545\ : InMux
    port map (
            O => \N__15427\,
            I => \N__15424\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__15424\,
            I => \b2v_inst200.count_0_16\
        );

    \I__1543\ : InMux
    port map (
            O => \N__15421\,
            I => \N__15418\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__15418\,
            I => \b2v_inst200.count_0_17\
        );

    \I__1541\ : CascadeMux
    port map (
            O => \N__15415\,
            I => \b2v_inst16.un13_clk_100khz_i_cascade_\
        );

    \I__1540\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15409\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__15409\,
            I => \b2v_inst16.count_4_0\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__15406\,
            I => \b2v_inst16.count_rst_5_cascade_\
        );

    \I__1537\ : InMux
    port map (
            O => \N__15403\,
            I => \N__15400\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__15400\,
            I => \b2v_inst16.count_4_13\
        );

    \I__1535\ : InMux
    port map (
            O => \N__15397\,
            I => \N__15391\
        );

    \I__1534\ : InMux
    port map (
            O => \N__15396\,
            I => \N__15391\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__15391\,
            I => \b2v_inst16.count_rst_2\
        );

    \I__1532\ : InMux
    port map (
            O => \N__15388\,
            I => \N__15385\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__15385\,
            I => \b2v_inst16.countZ0Z_13\
        );

    \I__1530\ : InMux
    port map (
            O => \N__15382\,
            I => \N__15372\
        );

    \I__1529\ : InMux
    port map (
            O => \N__15381\,
            I => \N__15372\
        );

    \I__1528\ : InMux
    port map (
            O => \N__15380\,
            I => \N__15369\
        );

    \I__1527\ : InMux
    port map (
            O => \N__15379\,
            I => \N__15362\
        );

    \I__1526\ : InMux
    port map (
            O => \N__15378\,
            I => \N__15362\
        );

    \I__1525\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15362\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__15372\,
            I => \b2v_inst16.countZ0Z_0\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__15369\,
            I => \b2v_inst16.countZ0Z_0\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__15362\,
            I => \b2v_inst16.countZ0Z_0\
        );

    \I__1521\ : CascadeMux
    port map (
            O => \N__15355\,
            I => \b2v_inst16.countZ0Z_13_cascade_\
        );

    \I__1520\ : InMux
    port map (
            O => \N__15352\,
            I => \N__15349\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__15349\,
            I => \b2v_inst16.un13_clk_100khz_11\
        );

    \I__1518\ : InMux
    port map (
            O => \N__15346\,
            I => \N__15342\
        );

    \I__1517\ : InMux
    port map (
            O => \N__15345\,
            I => \N__15339\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__15342\,
            I => \b2v_inst16.countZ0Z_15\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__15339\,
            I => \b2v_inst16.countZ0Z_15\
        );

    \I__1514\ : InMux
    port map (
            O => \N__15334\,
            I => \N__15328\
        );

    \I__1513\ : InMux
    port map (
            O => \N__15333\,
            I => \N__15328\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__15328\,
            I => \b2v_inst16.count_rst_4\
        );

    \I__1511\ : InMux
    port map (
            O => \N__15325\,
            I => \N__15322\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__15322\,
            I => \b2v_inst16.count_4_15\
        );

    \I__1509\ : InMux
    port map (
            O => \N__15319\,
            I => \N__15316\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__15316\,
            I => \b2v_inst16.count_4_14\
        );

    \I__1507\ : InMux
    port map (
            O => \N__15313\,
            I => \N__15309\
        );

    \I__1506\ : InMux
    port map (
            O => \N__15312\,
            I => \N__15306\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__15309\,
            I => \b2v_inst16.count_rst_3\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__15306\,
            I => \b2v_inst16.count_rst_3\
        );

    \I__1503\ : InMux
    port map (
            O => \N__15301\,
            I => \N__15297\
        );

    \I__1502\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15294\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__15297\,
            I => \b2v_inst16.countZ0Z_14\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__15294\,
            I => \b2v_inst16.countZ0Z_14\
        );

    \I__1499\ : InMux
    port map (
            O => \N__15289\,
            I => \N__15285\
        );

    \I__1498\ : InMux
    port map (
            O => \N__15288\,
            I => \N__15282\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__15285\,
            I => \b2v_inst16.count_rst_12\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__15282\,
            I => \b2v_inst16.count_rst_12\
        );

    \I__1495\ : InMux
    port map (
            O => \N__15277\,
            I => \N__15274\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__15274\,
            I => \b2v_inst16.count_4_7\
        );

    \I__1493\ : InMux
    port map (
            O => \N__15271\,
            I => \N__15267\
        );

    \I__1492\ : InMux
    port map (
            O => \N__15270\,
            I => \N__15264\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__15267\,
            I => \b2v_inst16.count_rst_9\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__15264\,
            I => \b2v_inst16.count_rst_9\
        );

    \I__1489\ : InMux
    port map (
            O => \N__15259\,
            I => \N__15256\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__15256\,
            I => \b2v_inst16.count_4_4\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__15253\,
            I => \b2v_inst16.count_rst_6_cascade_\
        );

    \I__1486\ : InMux
    port map (
            O => \N__15250\,
            I => \N__15247\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__15247\,
            I => \b2v_inst16.count_rst_6\
        );

    \I__1484\ : InMux
    port map (
            O => \N__15244\,
            I => \N__15241\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__15241\,
            I => \N__15237\
        );

    \I__1482\ : InMux
    port map (
            O => \N__15240\,
            I => \N__15234\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__15237\,
            I => \b2v_inst16.countZ0Z_11\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__15234\,
            I => \b2v_inst16.countZ0Z_11\
        );

    \I__1479\ : CascadeMux
    port map (
            O => \N__15229\,
            I => \b2v_inst16.countZ0Z_1_cascade_\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__15226\,
            I => \N__15223\
        );

    \I__1477\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15218\
        );

    \I__1476\ : InMux
    port map (
            O => \N__15222\,
            I => \N__15213\
        );

    \I__1475\ : InMux
    port map (
            O => \N__15221\,
            I => \N__15213\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__15218\,
            I => \N__15210\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__15213\,
            I => \b2v_inst16.un4_count_1_axb_1\
        );

    \I__1472\ : Odrv4
    port map (
            O => \N__15210\,
            I => \b2v_inst16.un4_count_1_axb_1\
        );

    \I__1471\ : InMux
    port map (
            O => \N__15205\,
            I => \N__15199\
        );

    \I__1470\ : InMux
    port map (
            O => \N__15204\,
            I => \N__15199\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__15199\,
            I => \b2v_inst16.count_4_1\
        );

    \I__1468\ : InMux
    port map (
            O => \N__15196\,
            I => \N__15193\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__15193\,
            I => \N__15189\
        );

    \I__1466\ : InMux
    port map (
            O => \N__15192\,
            I => \N__15186\
        );

    \I__1465\ : Span4Mux_s1_v
    port map (
            O => \N__15189\,
            I => \N__15183\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__15186\,
            I => \N__15180\
        );

    \I__1463\ : Odrv4
    port map (
            O => \N__15183\,
            I => \b2v_inst16.countZ0Z_2\
        );

    \I__1462\ : Odrv4
    port map (
            O => \N__15180\,
            I => \b2v_inst16.countZ0Z_2\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__15175\,
            I => \N__15172\
        );

    \I__1460\ : InMux
    port map (
            O => \N__15172\,
            I => \N__15168\
        );

    \I__1459\ : InMux
    port map (
            O => \N__15171\,
            I => \N__15165\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__15168\,
            I => \N__15162\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__15165\,
            I => \N__15159\
        );

    \I__1456\ : Odrv4
    port map (
            O => \N__15162\,
            I => \b2v_inst16.countZ0Z_6\
        );

    \I__1455\ : Odrv4
    port map (
            O => \N__15159\,
            I => \b2v_inst16.countZ0Z_6\
        );

    \I__1454\ : InMux
    port map (
            O => \N__15154\,
            I => \N__15151\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__15151\,
            I => \N__15147\
        );

    \I__1452\ : InMux
    port map (
            O => \N__15150\,
            I => \N__15144\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__15147\,
            I => \b2v_inst16.countZ0Z_12\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__15144\,
            I => \b2v_inst16.countZ0Z_12\
        );

    \I__1449\ : InMux
    port map (
            O => \N__15139\,
            I => \N__15136\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__15136\,
            I => \b2v_inst16.un13_clk_100khz_9\
        );

    \I__1447\ : InMux
    port map (
            O => \N__15133\,
            I => \N__15130\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__15130\,
            I => \b2v_inst16.un13_clk_100khz_8\
        );

    \I__1445\ : CascadeMux
    port map (
            O => \N__15127\,
            I => \b2v_inst16.un13_clk_100khz_10_cascade_\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__15124\,
            I => \b2v_inst11.count_off_1_3_cascade_\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__15121\,
            I => \N__15118\
        );

    \I__1442\ : InMux
    port map (
            O => \N__15118\,
            I => \N__15115\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__15115\,
            I => \N__15112\
        );

    \I__1440\ : Odrv4
    port map (
            O => \N__15112\,
            I => \b2v_inst11.un3_count_off_1_axb_3\
        );

    \I__1439\ : CascadeMux
    port map (
            O => \N__15109\,
            I => \N__15106\
        );

    \I__1438\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15103\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__15103\,
            I => \N__15100\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__15100\,
            I => \b2v_inst11.count_offZ0Z_4\
        );

    \I__1435\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15094\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__15094\,
            I => \b2v_inst11.count_off_1_3\
        );

    \I__1433\ : CascadeMux
    port map (
            O => \N__15091\,
            I => \b2v_inst11.count_offZ0Z_4_cascade_\
        );

    \I__1432\ : InMux
    port map (
            O => \N__15088\,
            I => \N__15085\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__15085\,
            I => \N__15082\
        );

    \I__1430\ : Odrv4
    port map (
            O => \N__15082\,
            I => \b2v_inst11.un34_clk_100khz_2\
        );

    \I__1429\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15073\
        );

    \I__1428\ : InMux
    port map (
            O => \N__15078\,
            I => \N__15073\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__15073\,
            I => \N__15070\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__15070\,
            I => \b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362\
        );

    \I__1425\ : InMux
    port map (
            O => \N__15067\,
            I => \N__15061\
        );

    \I__1424\ : InMux
    port map (
            O => \N__15066\,
            I => \N__15061\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__15061\,
            I => \b2v_inst11.count_offZ0Z_3\
        );

    \I__1422\ : InMux
    port map (
            O => \N__15058\,
            I => \N__15052\
        );

    \I__1421\ : InMux
    port map (
            O => \N__15057\,
            I => \N__15052\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__15052\,
            I => \N__15049\
        );

    \I__1419\ : Odrv4
    port map (
            O => \N__15049\,
            I => \b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__15046\,
            I => \N__15043\
        );

    \I__1417\ : InMux
    port map (
            O => \N__15043\,
            I => \N__15040\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__15040\,
            I => \b2v_inst11.count_off_0_4\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__15037\,
            I => \N__15034\
        );

    \I__1414\ : InMux
    port map (
            O => \N__15034\,
            I => \N__15031\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__15031\,
            I => \b2v_inst11.count_off_0_14\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__15028\,
            I => \N__15025\
        );

    \I__1411\ : InMux
    port map (
            O => \N__15025\,
            I => \N__15019\
        );

    \I__1410\ : InMux
    port map (
            O => \N__15024\,
            I => \N__15019\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__15019\,
            I => \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5\
        );

    \I__1408\ : InMux
    port map (
            O => \N__15016\,
            I => \b2v_inst11.un3_count_off_1_cry_6\
        );

    \I__1407\ : InMux
    port map (
            O => \N__15013\,
            I => \b2v_inst11.un3_count_off_1_cry_7\
        );

    \I__1406\ : InMux
    port map (
            O => \N__15010\,
            I => \bfn_1_15_0_\
        );

    \I__1405\ : InMux
    port map (
            O => \N__15007\,
            I => \b2v_inst11.un3_count_off_1_cry_9\
        );

    \I__1404\ : InMux
    port map (
            O => \N__15004\,
            I => \b2v_inst11.un3_count_off_1_cry_10\
        );

    \I__1403\ : InMux
    port map (
            O => \N__15001\,
            I => \b2v_inst11.un3_count_off_1_cry_11\
        );

    \I__1402\ : InMux
    port map (
            O => \N__14998\,
            I => \b2v_inst11.un3_count_off_1_cry_12\
        );

    \I__1401\ : InMux
    port map (
            O => \N__14995\,
            I => \b2v_inst11.un3_count_off_1_cry_13\
        );

    \I__1400\ : InMux
    port map (
            O => \N__14992\,
            I => \b2v_inst11.un3_count_off_1_cry_14\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__14989\,
            I => \b2v_inst11.un34_clk_100khz_1_cascade_\
        );

    \I__1398\ : InMux
    port map (
            O => \N__14986\,
            I => \N__14983\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__14983\,
            I => \b2v_inst11.un34_clk_100khz_0\
        );

    \I__1396\ : InMux
    port map (
            O => \N__14980\,
            I => \N__14977\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__14977\,
            I => \b2v_inst11.count_off_0_5\
        );

    \I__1394\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14971\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__14971\,
            I => \b2v_inst11.un3_count_off_1_axb_2\
        );

    \I__1392\ : InMux
    port map (
            O => \N__14968\,
            I => \N__14962\
        );

    \I__1391\ : InMux
    port map (
            O => \N__14967\,
            I => \N__14962\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__14962\,
            I => \b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152\
        );

    \I__1389\ : InMux
    port map (
            O => \N__14959\,
            I => \b2v_inst11.un3_count_off_1_cry_1\
        );

    \I__1388\ : InMux
    port map (
            O => \N__14956\,
            I => \b2v_inst11.un3_count_off_1_cry_2_cZ0\
        );

    \I__1387\ : InMux
    port map (
            O => \N__14953\,
            I => \b2v_inst11.un3_count_off_1_cry_3_cZ0\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__14950\,
            I => \N__14946\
        );

    \I__1385\ : InMux
    port map (
            O => \N__14949\,
            I => \N__14943\
        );

    \I__1384\ : InMux
    port map (
            O => \N__14946\,
            I => \N__14940\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__14943\,
            I => \b2v_inst11.count_offZ0Z_5\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__14940\,
            I => \b2v_inst11.count_offZ0Z_5\
        );

    \I__1381\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14929\
        );

    \I__1380\ : InMux
    port map (
            O => \N__14934\,
            I => \N__14929\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__14929\,
            I => \b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882\
        );

    \I__1378\ : InMux
    port map (
            O => \N__14926\,
            I => \b2v_inst11.un3_count_off_1_cry_4_cZ0\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__14923\,
            I => \N__14920\
        );

    \I__1376\ : InMux
    port map (
            O => \N__14920\,
            I => \N__14917\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__14917\,
            I => \N__14914\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__14914\,
            I => \b2v_inst11.un3_count_off_1_axb_6\
        );

    \I__1373\ : InMux
    port map (
            O => \N__14911\,
            I => \b2v_inst11.un3_count_off_1_cry_5\
        );

    \I__1372\ : InMux
    port map (
            O => \N__14908\,
            I => \N__14902\
        );

    \I__1371\ : InMux
    port map (
            O => \N__14907\,
            I => \N__14902\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__14902\,
            I => \N__14899\
        );

    \I__1369\ : Odrv4
    port map (
            O => \N__14899\,
            I => \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5\
        );

    \I__1368\ : InMux
    port map (
            O => \N__14896\,
            I => \N__14893\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__14893\,
            I => \b2v_inst11.count_clk_0_4\
        );

    \I__1366\ : InMux
    port map (
            O => \N__14890\,
            I => \N__14887\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__14887\,
            I => \b2v_inst11.count_off_1_2\
        );

    \I__1364\ : InMux
    port map (
            O => \N__14884\,
            I => \N__14878\
        );

    \I__1363\ : InMux
    port map (
            O => \N__14883\,
            I => \N__14878\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__14878\,
            I => \b2v_inst11.count_offZ0Z_2\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__14875\,
            I => \b2v_inst11.count_off_1_2_cascade_\
        );

    \I__1360\ : InMux
    port map (
            O => \N__14872\,
            I => \N__14869\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__14869\,
            I => \N__14865\
        );

    \I__1358\ : InMux
    port map (
            O => \N__14868\,
            I => \N__14862\
        );

    \I__1357\ : Odrv4
    port map (
            O => \N__14865\,
            I => \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__14862\,
            I => \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0\
        );

    \I__1355\ : InMux
    port map (
            O => \N__14857\,
            I => \N__14854\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__14854\,
            I => \b2v_inst11.count_clk_0_15\
        );

    \I__1353\ : InMux
    port map (
            O => \N__14851\,
            I => \N__14845\
        );

    \I__1352\ : InMux
    port map (
            O => \N__14850\,
            I => \N__14845\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__14845\,
            I => \N__14842\
        );

    \I__1350\ : Odrv4
    port map (
            O => \N__14842\,
            I => \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\
        );

    \I__1349\ : InMux
    port map (
            O => \N__14839\,
            I => \N__14836\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__14836\,
            I => \b2v_inst11.count_clk_0_6\
        );

    \I__1347\ : CascadeMux
    port map (
            O => \N__14833\,
            I => \N__14829\
        );

    \I__1346\ : InMux
    port map (
            O => \N__14832\,
            I => \N__14824\
        );

    \I__1345\ : InMux
    port map (
            O => \N__14829\,
            I => \N__14824\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__14824\,
            I => \N__14821\
        );

    \I__1343\ : Odrv4
    port map (
            O => \N__14821\,
            I => \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5\
        );

    \I__1342\ : InMux
    port map (
            O => \N__14818\,
            I => \N__14815\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__14815\,
            I => \b2v_inst11.count_clk_0_8\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__14812\,
            I => \N__14808\
        );

    \I__1339\ : InMux
    port map (
            O => \N__14811\,
            I => \N__14803\
        );

    \I__1338\ : InMux
    port map (
            O => \N__14808\,
            I => \N__14803\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__14803\,
            I => \N__14800\
        );

    \I__1336\ : Odrv4
    port map (
            O => \N__14800\,
            I => \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5\
        );

    \I__1335\ : InMux
    port map (
            O => \N__14797\,
            I => \N__14794\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__14794\,
            I => \b2v_inst11.count_clk_0_7\
        );

    \I__1333\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14785\
        );

    \I__1332\ : InMux
    port map (
            O => \N__14790\,
            I => \N__14785\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__14785\,
            I => \N__14782\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__14782\,
            I => \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5\
        );

    \I__1329\ : InMux
    port map (
            O => \N__14779\,
            I => \N__14776\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__14776\,
            I => \b2v_inst11.count_clk_0_9\
        );

    \I__1327\ : InMux
    port map (
            O => \N__14773\,
            I => \b2v_inst11.un1_count_clk_2_cry_9_cZ0\
        );

    \I__1326\ : InMux
    port map (
            O => \N__14770\,
            I => \b2v_inst11.un1_count_clk_2_cry_10_cZ0\
        );

    \I__1325\ : InMux
    port map (
            O => \N__14767\,
            I => \b2v_inst11.un1_count_clk_2_cry_11\
        );

    \I__1324\ : InMux
    port map (
            O => \N__14764\,
            I => \b2v_inst11.un1_count_clk_2_cry_12\
        );

    \I__1323\ : InMux
    port map (
            O => \N__14761\,
            I => \b2v_inst11.un1_count_clk_2_cry_13\
        );

    \I__1322\ : InMux
    port map (
            O => \N__14758\,
            I => \b2v_inst11.un1_count_clk_2_cry_14\
        );

    \I__1321\ : InMux
    port map (
            O => \N__14755\,
            I => \N__14749\
        );

    \I__1320\ : InMux
    port map (
            O => \N__14754\,
            I => \N__14749\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__14749\,
            I => \N__14746\
        );

    \I__1318\ : Odrv4
    port map (
            O => \N__14746\,
            I => \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5\
        );

    \I__1317\ : InMux
    port map (
            O => \N__14743\,
            I => \N__14740\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__14740\,
            I => \b2v_inst11.count_clk_0_5\
        );

    \I__1315\ : InMux
    port map (
            O => \N__14737\,
            I => \b2v_inst11.un1_count_clk_2_cry_1\
        );

    \I__1314\ : InMux
    port map (
            O => \N__14734\,
            I => \b2v_inst11.un1_count_clk_2_cry_2\
        );

    \I__1313\ : InMux
    port map (
            O => \N__14731\,
            I => \b2v_inst11.un1_count_clk_2_cry_3\
        );

    \I__1312\ : InMux
    port map (
            O => \N__14728\,
            I => \b2v_inst11.un1_count_clk_2_cry_4\
        );

    \I__1311\ : InMux
    port map (
            O => \N__14725\,
            I => \b2v_inst11.un1_count_clk_2_cry_5\
        );

    \I__1310\ : InMux
    port map (
            O => \N__14722\,
            I => \b2v_inst11.un1_count_clk_2_cry_6\
        );

    \I__1309\ : InMux
    port map (
            O => \N__14719\,
            I => \b2v_inst11.un1_count_clk_2_cry_7_cZ0\
        );

    \I__1308\ : InMux
    port map (
            O => \N__14716\,
            I => \bfn_1_10_0_\
        );

    \I__1307\ : InMux
    port map (
            O => \N__14713\,
            I => \N__14710\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__14710\,
            I => \b2v_inst200.count_2_5\
        );

    \I__1305\ : InMux
    port map (
            O => \N__14707\,
            I => \N__14704\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__14704\,
            I => \b2v_inst200.count_2_9\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__14701\,
            I => \b2v_inst200.countZ0Z_9_cascade_\
        );

    \I__1302\ : InMux
    port map (
            O => \N__14698\,
            I => \N__14695\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__14695\,
            I => \N__14692\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__14692\,
            I => \b2v_inst200.un25_clk_100khz_9\
        );

    \I__1299\ : InMux
    port map (
            O => \N__14689\,
            I => \N__14686\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__14686\,
            I => \b2v_inst200.count_2_12\
        );

    \I__1297\ : InMux
    port map (
            O => \N__14683\,
            I => \N__14680\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__14680\,
            I => \b2v_inst200.count_2_13\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__14677\,
            I => \b2v_inst200.countZ0Z_0_cascade_\
        );

    \I__1294\ : InMux
    port map (
            O => \N__14674\,
            I => \N__14671\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__14671\,
            I => \b2v_inst200.un25_clk_100khz_13\
        );

    \I__1292\ : InMux
    port map (
            O => \N__14668\,
            I => \N__14665\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__14665\,
            I => \b2v_inst200.count_2_6\
        );

    \I__1290\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14659\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__14659\,
            I => \b2v_inst200.count_2_14\
        );

    \I__1288\ : InMux
    port map (
            O => \N__14656\,
            I => \N__14653\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__14653\,
            I => \N__14650\
        );

    \I__1286\ : Odrv4
    port map (
            O => \N__14650\,
            I => \b2v_inst200.un25_clk_100khz_10\
        );

    \I__1285\ : InMux
    port map (
            O => \N__14647\,
            I => \N__14644\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__14644\,
            I => \b2v_inst200.count_2_3\
        );

    \I__1283\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14638\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__14638\,
            I => \b2v_inst200.count_2_4\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__14635\,
            I => \b2v_inst200.count_RNI_0_0_cascade_\
        );

    \I__1280\ : InMux
    port map (
            O => \N__14632\,
            I => \N__14629\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__14629\,
            I => \b2v_inst200.count_2_11\
        );

    \I__1278\ : InMux
    port map (
            O => \N__14626\,
            I => \N__14623\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__14623\,
            I => \b2v_inst200.count_2_10\
        );

    \I__1276\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14617\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__14617\,
            I => \b2v_inst200.count_2_8\
        );

    \I__1274\ : InMux
    port map (
            O => \N__14614\,
            I => \N__14611\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__14611\,
            I => \b2v_inst200.count_2_0\
        );

    \I__1272\ : InMux
    port map (
            O => \N__14608\,
            I => \N__14602\
        );

    \I__1271\ : InMux
    port map (
            O => \N__14607\,
            I => \N__14602\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__14602\,
            I => \b2v_inst16.count_rst_1\
        );

    \I__1269\ : InMux
    port map (
            O => \N__14599\,
            I => \N__14596\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__14596\,
            I => \b2v_inst16.count_4_12\
        );

    \I__1267\ : InMux
    port map (
            O => \N__14593\,
            I => \N__14587\
        );

    \I__1266\ : InMux
    port map (
            O => \N__14592\,
            I => \N__14587\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__14587\,
            I => \b2v_inst16.count_rst_0\
        );

    \I__1264\ : InMux
    port map (
            O => \N__14584\,
            I => \N__14581\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__14581\,
            I => \b2v_inst16.count_4_11\
        );

    \I__1262\ : InMux
    port map (
            O => \N__14578\,
            I => \N__14572\
        );

    \I__1261\ : InMux
    port map (
            O => \N__14577\,
            I => \N__14572\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__14572\,
            I => \N__14569\
        );

    \I__1259\ : Odrv4
    port map (
            O => \N__14569\,
            I => \b2v_inst16.count_rst_11\
        );

    \I__1258\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14563\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__14563\,
            I => \b2v_inst16.count_4_6\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__14560\,
            I => \b2v_inst200.un25_clk_100khz_12_cascade_\
        );

    \I__1255\ : CascadeMux
    port map (
            O => \N__14557\,
            I => \b2v_inst200.count_RNIC03N_3Z0Z_0_cascade_\
        );

    \I__1254\ : InMux
    port map (
            O => \N__14554\,
            I => \b2v_inst16.un4_count_1_cry_9\
        );

    \I__1253\ : InMux
    port map (
            O => \N__14551\,
            I => \b2v_inst16.un4_count_1_cry_10_cZ0\
        );

    \I__1252\ : InMux
    port map (
            O => \N__14548\,
            I => \b2v_inst16.un4_count_1_cry_11\
        );

    \I__1251\ : InMux
    port map (
            O => \N__14545\,
            I => \b2v_inst16.un4_count_1_cry_12\
        );

    \I__1250\ : InMux
    port map (
            O => \N__14542\,
            I => \b2v_inst16.un4_count_1_cry_13\
        );

    \I__1249\ : InMux
    port map (
            O => \N__14539\,
            I => \b2v_inst16.un4_count_1_cry_14\
        );

    \I__1248\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14530\
        );

    \I__1247\ : InMux
    port map (
            O => \N__14535\,
            I => \N__14530\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__14530\,
            I => \N__14527\
        );

    \I__1245\ : Odrv4
    port map (
            O => \N__14527\,
            I => \b2v_inst16.count_rst_7\
        );

    \I__1244\ : InMux
    port map (
            O => \N__14524\,
            I => \N__14521\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__14521\,
            I => \b2v_inst16.count_4_2\
        );

    \I__1242\ : InMux
    port map (
            O => \N__14518\,
            I => \b2v_inst16.un4_count_1_cry_1\
        );

    \I__1241\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14511\
        );

    \I__1240\ : InMux
    port map (
            O => \N__14514\,
            I => \N__14508\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__14511\,
            I => \b2v_inst16.countZ0Z_3\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__14508\,
            I => \b2v_inst16.countZ0Z_3\
        );

    \I__1237\ : InMux
    port map (
            O => \N__14503\,
            I => \N__14497\
        );

    \I__1236\ : InMux
    port map (
            O => \N__14502\,
            I => \N__14497\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__14497\,
            I => \b2v_inst16.count_rst_8\
        );

    \I__1234\ : InMux
    port map (
            O => \N__14494\,
            I => \b2v_inst16.un4_count_1_cry_2_cZ0\
        );

    \I__1233\ : InMux
    port map (
            O => \N__14491\,
            I => \N__14487\
        );

    \I__1232\ : InMux
    port map (
            O => \N__14490\,
            I => \N__14484\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__14487\,
            I => \b2v_inst16.countZ0Z_4\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__14484\,
            I => \b2v_inst16.countZ0Z_4\
        );

    \I__1229\ : InMux
    port map (
            O => \N__14479\,
            I => \b2v_inst16.un4_count_1_cry_3\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__14476\,
            I => \N__14473\
        );

    \I__1227\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14469\
        );

    \I__1226\ : InMux
    port map (
            O => \N__14472\,
            I => \N__14466\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__14469\,
            I => \b2v_inst16.countZ0Z_5\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__14466\,
            I => \b2v_inst16.countZ0Z_5\
        );

    \I__1223\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14455\
        );

    \I__1222\ : InMux
    port map (
            O => \N__14460\,
            I => \N__14455\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__14455\,
            I => \b2v_inst16.count_rst_10\
        );

    \I__1220\ : InMux
    port map (
            O => \N__14452\,
            I => \b2v_inst16.un4_count_1_cry_4\
        );

    \I__1219\ : InMux
    port map (
            O => \N__14449\,
            I => \b2v_inst16.un4_count_1_cry_5\
        );

    \I__1218\ : InMux
    port map (
            O => \N__14446\,
            I => \N__14442\
        );

    \I__1217\ : InMux
    port map (
            O => \N__14445\,
            I => \N__14439\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__14442\,
            I => \b2v_inst16.countZ0Z_7\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__14439\,
            I => \b2v_inst16.countZ0Z_7\
        );

    \I__1214\ : InMux
    port map (
            O => \N__14434\,
            I => \b2v_inst16.un4_count_1_cry_6\
        );

    \I__1213\ : InMux
    port map (
            O => \N__14431\,
            I => \b2v_inst16.un4_count_1_cry_7\
        );

    \I__1212\ : InMux
    port map (
            O => \N__14428\,
            I => \bfn_1_3_0_\
        );

    \I__1211\ : InMux
    port map (
            O => \N__14425\,
            I => \N__14422\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__14422\,
            I => \b2v_inst16.count_4_3\
        );

    \I__1209\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14416\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__14416\,
            I => \b2v_inst16.count_4_5\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst6.un2_count_1_cry_8\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst5.un2_count_1_cry_8\,
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_9_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_1_0_\
        );

    \IN_MUX_bfv_9_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst36.un2_count_1_cry_8\,
            carryinitout => \bfn_9_2_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => b2v_inst20_un4_counter_7,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst20.counter_1_cry_8\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst20.counter_1_cry_16\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst20.counter_1_cry_24\,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_1_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_2_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst16.un4_count_1_cry_8\,
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un3_count_off_1_cry_8\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_4_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_1_0_\
        );

    \IN_MUX_bfv_4_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_2_0_\
        );

    \IN_MUX_bfv_4_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_3_0_\
        );

    \IN_MUX_bfv_4_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_4_0_\
        );

    \IN_MUX_bfv_5_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_4_0_\
        );

    \IN_MUX_bfv_5_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_5_0_\
        );

    \IN_MUX_bfv_5_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_6_0_\
        );

    \IN_MUX_bfv_4_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_6_0_\
        );

    \IN_MUX_bfv_9_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_4_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_7_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_2_0_\
        );

    \IN_MUX_bfv_7_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_3_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_6_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_2_0_\
        );

    \IN_MUX_bfv_6_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_1_0_\
        );

    \IN_MUX_bfv_5_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_1_0_\
        );

    \IN_MUX_bfv_5_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_2_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_count_cry_8\,
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_count_clk_2_cry_8_cZ0\,
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_2_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_6_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst200.un2_count_1_cry_7\,
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst200.un2_count_1_cry_15\,
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_7_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_5_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un85_clk_100khz_cry_7\,
            carryinitout => \bfn_7_6_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un85_clk_100khz_cry_15_cZ0\,
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_6_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_13_0_\
        );

    \IN_MUX_bfv_6_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_dutycycle_94_cry_7_cZ0\,
            carryinitout => \bfn_6_14_0_\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_dutycycle_53_cry_7_cZ0\,
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_dutycycle_53_cry_15\,
            carryinitout => \bfn_5_9_0_\
        );

    \b2v_inst200.count_en_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__17362\,
            GLOBALBUFFEROUTPUT => \b2v_inst200.count_en_g\
        );

    \b2v_inst16.delayed_vddq_pwrgd_en_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__27625\,
            GLOBALBUFFEROUTPUT => b2v_inst16_delayed_vddq_pwrgd_en_g
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_3_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14491\,
            in1 => \N__14446\,
            in2 => \N__14476\,
            in3 => \N__14515\,
            lcout => \b2v_inst16.un13_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIF7UJ1_3_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14425\,
            in1 => \N__14502\,
            in2 => \_gnd_net_\,
            in3 => \N__30624\,
            lcout => \b2v_inst16.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_3_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14503\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34638\,
            ce => \N__30629\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIHAVJ1_4_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15259\,
            in1 => \N__15270\,
            in2 => \_gnd_net_\,
            in3 => \N__30625\,
            lcout => \b2v_inst16.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIJD0K1_5_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14419\,
            in1 => \N__14460\,
            in2 => \_gnd_net_\,
            in3 => \N__30626\,
            lcout => \b2v_inst16.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_5_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14461\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34638\,
            ce => \N__30629\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNINJ2K1_7_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15277\,
            in1 => \N__15288\,
            in2 => \_gnd_net_\,
            in3 => \N__30627\,
            lcout => \b2v_inst16.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_1_c_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15380\,
            in2 => \N__15226\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_2_0_\,
            carryout => \b2v_inst16.un4_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15192\,
            in2 => \_gnd_net_\,
            in3 => \N__14518\,
            lcout => \b2v_inst16.count_rst_7\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_1\,
            carryout => \b2v_inst16.un4_count_1_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20340\,
            in1 => \N__14514\,
            in2 => \_gnd_net_\,
            in3 => \N__14494\,
            lcout => \b2v_inst16.count_rst_8\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_2_cZ0\,
            carryout => \b2v_inst16.un4_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20343\,
            in1 => \N__14490\,
            in2 => \_gnd_net_\,
            in3 => \N__14479\,
            lcout => \b2v_inst16.count_rst_9\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_3\,
            carryout => \b2v_inst16.un4_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20341\,
            in1 => \N__14472\,
            in2 => \_gnd_net_\,
            in3 => \N__14452\,
            lcout => \b2v_inst16.count_rst_10\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_4\,
            carryout => \b2v_inst16.un4_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15171\,
            in2 => \_gnd_net_\,
            in3 => \N__14449\,
            lcout => \b2v_inst16.count_rst_11\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_5\,
            carryout => \b2v_inst16.un4_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20342\,
            in1 => \N__14445\,
            in2 => \_gnd_net_\,
            in3 => \N__14434\,
            lcout => \b2v_inst16.count_rst_12\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_6\,
            carryout => \b2v_inst16.un4_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20344\,
            in1 => \N__30198\,
            in2 => \_gnd_net_\,
            in3 => \N__14431\,
            lcout => \b2v_inst16.count_rst_13\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_7\,
            carryout => \b2v_inst16.un4_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20346\,
            in1 => \_gnd_net_\,
            in2 => \N__30150\,
            in3 => \N__14428\,
            lcout => \b2v_inst16.count_rst_14\,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => \b2v_inst16.un4_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17319\,
            in2 => \_gnd_net_\,
            in3 => \N__14554\,
            lcout => \b2v_inst16.count_rst\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_9\,
            carryout => \b2v_inst16.un4_count_1_cry_10_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_10_c_RNIDGU31_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20345\,
            in1 => \N__15240\,
            in2 => \_gnd_net_\,
            in3 => \N__14551\,
            lcout => \b2v_inst16.count_rst_0\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_10_cZ0\,
            carryout => \b2v_inst16.un4_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15150\,
            in2 => \_gnd_net_\,
            in3 => \N__14548\,
            lcout => \b2v_inst16.count_rst_1\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_11\,
            carryout => \b2v_inst16.un4_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15388\,
            in2 => \_gnd_net_\,
            in3 => \N__14545\,
            lcout => \b2v_inst16.count_rst_2\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_12\,
            carryout => \b2v_inst16.un4_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15300\,
            in2 => \_gnd_net_\,
            in3 => \N__14542\,
            lcout => \b2v_inst16.count_rst_3\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_13\,
            carryout => \b2v_inst16.un4_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15346\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14539\,
            lcout => \b2v_inst16.count_rst_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_14_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15313\,
            lcout => \b2v_inst16.count_4_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34626\,
            ce => \N__30622\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNID4TJ1_2_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14524\,
            in1 => \N__14535\,
            in2 => \_gnd_net_\,
            in3 => \N__30630\,
            lcout => \b2v_inst16.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_2_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14536\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34622\,
            ce => \N__30628\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIFJV31_12_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14599\,
            in1 => \N__14607\,
            in2 => \_gnd_net_\,
            in3 => \N__30633\,
            lcout => \b2v_inst16.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_12_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14608\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34622\,
            ce => \N__30628\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIJM901_11_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14584\,
            in1 => \N__14592\,
            in2 => \_gnd_net_\,
            in3 => \N__30632\,
            lcout => \b2v_inst16.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_11_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14593\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34622\,
            ce => \N__30628\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNILG1K1_6_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14577\,
            in1 => \N__14566\,
            in2 => \_gnd_net_\,
            in3 => \N__30631\,
            lcout => \b2v_inst16.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_6_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14578\,
            lcout => \b2v_inst16.count_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34622\,
            ce => \N__30628\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_6_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15948\,
            in1 => \N__15843\,
            in2 => \N__15813\,
            in3 => \N__15891\,
            lcout => OPEN,
            ltout => \b2v_inst200.un25_clk_100khz_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIC03N_3_0_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14656\,
            in1 => \N__14674\,
            in2 => \N__14560\,
            in3 => \N__15433\,
            lcout => \b2v_inst200.count_RNIC03N_3Z0Z_0\,
            ltout => \b2v_inst200.count_RNIC03N_3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_0_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14557\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_RNI_0_0\,
            ltout => \b2v_inst200.count_RNI_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI96451_6_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__14668\,
            in1 => \N__15937\,
            in2 => \N__14635\,
            in3 => \N__15719\,
            lcout => \b2v_inst200.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI1QM71_11_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__15796\,
            in1 => \N__14632\,
            in2 => \N__33604\,
            in3 => \N__15721\,
            lcout => \b2v_inst200.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_11_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15795\,
            in2 => \_gnd_net_\,
            in3 => \N__33591\,
            lcout => \b2v_inst200.count_2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34617\,
            ce => \N__15659\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_10_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33590\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15828\,
            lcout => \b2v_inst200.count_2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34617\,
            ce => \N__15659\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIOMPC1_10_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__14626\,
            in1 => \N__33586\,
            in2 => \N__15832\,
            in3 => \N__15720\,
            lcout => \b2v_inst200.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIDC651_8_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__14620\,
            in1 => \N__33592\,
            in2 => \N__15880\,
            in3 => \N__15718\,
            lcout => \b2v_inst200.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_8_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33594\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15876\,
            lcout => \b2v_inst200.count_2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34615\,
            ce => \N__15658\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI73Q71_14_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14662\,
            in1 => \N__16074\,
            in2 => \_gnd_net_\,
            in3 => \N__15716\,
            lcout => \b2v_inst200.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_0_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__33593\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15607\,
            lcout => \b2v_inst200.count_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34615\,
            ce => \N__15658\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIC03N_0_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14614\,
            in1 => \N__15595\,
            in2 => \_gnd_net_\,
            in3 => \N__15717\,
            lcout => \b2v_inst200.countZ0Z_0\,
            ltout => \b2v_inst200.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIC03N_1_0_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14698\,
            in2 => \N__14677\,
            in3 => \N__16087\,
            lcout => \b2v_inst200.un25_clk_100khz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_6_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15936\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33595\,
            lcout => \b2v_inst200.count_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34615\,
            ce => \N__15658\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_14_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16075\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34615\,
            ce => \N__15658\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_3_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15481\,
            in1 => \N__15922\,
            in2 => \N__15508\,
            in3 => \N__15532\,
            lcout => \b2v_inst200.un25_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI3T051_3_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14647\,
            in1 => \N__15519\,
            in2 => \_gnd_net_\,
            in3 => \N__15708\,
            lcout => \b2v_inst200.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_3_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15520\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34611\,
            ce => \N__15657\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI50251_4_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15492\,
            in1 => \N__14641\,
            in2 => \_gnd_net_\,
            in3 => \N__15709\,
            lcout => \b2v_inst200.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_4_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15493\,
            lcout => \b2v_inst200.count_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34611\,
            ce => \N__15657\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI73351_5_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14713\,
            in1 => \N__15468\,
            in2 => \_gnd_net_\,
            in3 => \N__15710\,
            lcout => \b2v_inst200.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_5_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34611\,
            ce => \N__15657\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIB9551_7_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15445\,
            in1 => \N__15906\,
            in2 => \_gnd_net_\,
            in3 => \N__15711\,
            lcout => \b2v_inst200.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_9_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15859\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34609\,
            ce => \N__15656\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIFF751_9_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14707\,
            in1 => \N__15858\,
            in2 => \_gnd_net_\,
            in3 => \N__15712\,
            lcout => \b2v_inst200.countZ0Z_9\,
            ltout => \b2v_inst200.countZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_9_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15781\,
            in1 => \N__15757\,
            in2 => \N__14701\,
            in3 => \N__16063\,
            lcout => \b2v_inst200.un25_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI3TN71_12_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15768\,
            in1 => \N__14689\,
            in2 => \_gnd_net_\,
            in3 => \N__15713\,
            lcout => \b2v_inst200.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_12_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15769\,
            lcout => \b2v_inst200.count_2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34609\,
            ce => \N__15656\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI50P71_13_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14683\,
            in1 => \N__15744\,
            in2 => \_gnd_net_\,
            in3 => \N__15714\,
            lcout => \b2v_inst200.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_13_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15745\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_2_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34609\,
            ce => \N__15656\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI96R71_15_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15457\,
            in1 => \N__16047\,
            in2 => \_gnd_net_\,
            in3 => \N__15715\,
            lcout => \b2v_inst200.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_1_c_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16430\,
            in2 => \N__16696\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16606\,
            in1 => \N__16270\,
            in2 => \_gnd_net_\,
            in3 => \N__14737\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_1\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16600\,
            in1 => \N__16253\,
            in2 => \_gnd_net_\,
            in3 => \N__14734\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_2\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__16603\,
            in1 => \_gnd_net_\,
            in2 => \N__16297\,
            in3 => \N__14731\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_3\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__16601\,
            in1 => \_gnd_net_\,
            in2 => \N__16402\,
            in3 => \N__14728\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_4\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__16604\,
            in1 => \_gnd_net_\,
            in2 => \N__16318\,
            in3 => \N__14725\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_5\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__16602\,
            in1 => \_gnd_net_\,
            in2 => \N__16237\,
            in3 => \N__14722\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_6\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__16605\,
            in1 => \_gnd_net_\,
            in2 => \N__16339\,
            in3 => \N__14719\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_7_cZ0\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__16593\,
            in1 => \_gnd_net_\,
            in2 => \N__16717\,
            in3 => \N__14716\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_9_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16192\,
            in3 => \N__14773\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_9_cZ0\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_10_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16183\,
            in3 => \N__14770\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AAZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_10_cZ0\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16489\,
            in3 => \N__14767\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BAZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_11\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__16594\,
            in1 => \_gnd_net_\,
            in2 => \N__16117\,
            in3 => \N__14764\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CAZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_12\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__16618\,
            in1 => \_gnd_net_\,
            in2 => \N__16147\,
            in3 => \N__14761\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DAZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_13\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16595\,
            in1 => \N__16164\,
            in2 => \_gnd_net_\,
            in3 => \N__14758\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI0JFF5_5_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14743\,
            in1 => \N__17480\,
            in2 => \_gnd_net_\,
            in3 => \N__14754\,
            lcout => \b2v_inst11.count_clkZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_5_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14755\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34610\,
            ce => \N__17542\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI281F5_15_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14857\,
            in1 => \N__17483\,
            in2 => \_gnd_net_\,
            in3 => \N__14868\,
            lcout => \b2v_inst11.count_clkZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_15_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14872\,
            lcout => \b2v_inst11.count_clk_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34610\,
            ce => \N__17542\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI2MGF5_6_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14839\,
            in1 => \N__17481\,
            in2 => \_gnd_net_\,
            in3 => \N__14850\,
            lcout => \b2v_inst11.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_6_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14851\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34610\,
            ce => \N__17542\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI6SIF5_8_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__14818\,
            in1 => \N__17482\,
            in2 => \N__14833\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clkZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_8_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14832\,
            lcout => \b2v_inst11.count_clk_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34610\,
            ce => \N__17542\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI4PHF5_7_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14797\,
            in2 => \N__14812\,
            in3 => \N__17524\,
            lcout => \b2v_inst11.count_clkZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_7_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14811\,
            lcout => \b2v_inst11.count_clk_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34614\,
            ce => \N__17537\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI8VJF5_9_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14779\,
            in1 => \N__17525\,
            in2 => \_gnd_net_\,
            in3 => \N__14790\,
            lcout => \b2v_inst11.count_clkZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_9_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14791\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34614\,
            ce => \N__17537\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIUFEF5_4_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14896\,
            in1 => \N__17523\,
            in2 => \_gnd_net_\,
            in3 => \N__14907\,
            lcout => \b2v_inst11.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_4_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14908\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34614\,
            ce => \N__17537\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNINJ641_7_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__24328\,
            in1 => \N__23043\,
            in2 => \_gnd_net_\,
            in3 => \N__16641\,
            lcout => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNICG51A_6_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16752\,
            in1 => \N__18138\,
            in2 => \_gnd_net_\,
            in3 => \N__16923\,
            lcout => \b2v_inst11.un3_count_off_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_5_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14935\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19562\,
            lcout => \b2v_inst11.count_off_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34616\,
            ce => \N__18153\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI4411A_2_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14883\,
            in1 => \N__18130\,
            in2 => \_gnd_net_\,
            in3 => \N__14890\,
            lcout => \b2v_inst11.un3_count_off_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_2_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14968\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19561\,
            lcout => \b2v_inst11.count_offZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34616\,
            ce => \N__18153\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_1_c_RNIIQOD2_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19541\,
            in2 => \_gnd_net_\,
            in3 => \N__14967\,
            lcout => \b2v_inst11.count_off_1_2\,
            ltout => \b2v_inst11.count_off_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI4411A_0_2_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__18154\,
            in1 => \N__14884\,
            in2 => \N__14875\,
            in3 => \N__14949\,
            lcout => \b2v_inst11.un34_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNICG51A_0_6_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__16753\,
            in1 => \N__17911\,
            in2 => \N__16930\,
            in3 => \N__18155\,
            lcout => OPEN,
            ltout => \b2v_inst11.un34_clk_100khz_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI4FF481_2_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15088\,
            in1 => \N__17023\,
            in2 => \N__14989\,
            in3 => \N__14986\,
            lcout => \b2v_inst11.un34_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIAD41A_5_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__14980\,
            in1 => \N__18131\,
            in2 => \N__19581\,
            in3 => \N__14934\,
            lcout => \b2v_inst11.count_offZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_1_c_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17863\,
            in2 => \N__17910\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \b2v_inst11.un3_count_off_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14974\,
            in2 => \_gnd_net_\,
            in3 => \N__14959\,
            lcout => \b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_1\,
            carryout => \b2v_inst11.un3_count_off_1_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15121\,
            in3 => \N__14956\,
            lcout => \b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_2_cZ0\,
            carryout => \b2v_inst11.un3_count_off_1_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15109\,
            in3 => \N__14953\,
            lcout => \b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_3_cZ0\,
            carryout => \b2v_inst11.un3_count_off_1_cry_4_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14950\,
            in3 => \N__14926\,
            lcout => \b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_4_cZ0\,
            carryout => \b2v_inst11.un3_count_off_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14923\,
            in3 => \N__14911\,
            lcout => \b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_5\,
            carryout => \b2v_inst11.un3_count_off_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16990\,
            in3 => \N__15016\,
            lcout => \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_6\,
            carryout => \b2v_inst11.un3_count_off_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17038\,
            in3 => \N__15013\,
            lcout => \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_7\,
            carryout => \b2v_inst11.un3_count_off_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16948\,
            in3 => \N__15010\,
            lcout => \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \b2v_inst11.un3_count_off_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17800\,
            in3 => \N__15007\,
            lcout => \b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_9\,
            carryout => \b2v_inst11.un3_count_off_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16510\,
            in3 => \N__15004\,
            lcout => \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_10\,
            carryout => \b2v_inst11.un3_count_off_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16786\,
            in3 => \N__15001\,
            lcout => \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_11\,
            carryout => \b2v_inst11.un3_count_off_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16870\,
            in3 => \N__14998\,
            lcout => \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_12\,
            carryout => \b2v_inst11.un3_count_off_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16854\,
            in3 => \N__14995\,
            lcout => \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_13\,
            carryout => \b2v_inst11.un3_count_off_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16876\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14992\,
            lcout => \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI8V45A_13_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__19580\,
            in1 => \N__18137\,
            in2 => \N__18175\,
            in3 => \N__17772\,
            lcout => \b2v_inst11.count_offZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_2_c_RNIJSPD2_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19572\,
            in2 => \_gnd_net_\,
            in3 => \N__15078\,
            lcout => \b2v_inst11.count_off_1_3\,
            ltout => \b2v_inst11.count_off_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI6721A_3_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15066\,
            in2 => \N__15124\,
            in3 => \N__18132\,
            lcout => \b2v_inst11.un3_count_off_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI8A31A_4_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__18133\,
            in1 => \N__19573\,
            in2 => \N__15046\,
            in3 => \N__15057\,
            lcout => \b2v_inst11.count_offZ0Z_4\,
            ltout => \b2v_inst11.count_offZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI6721A_0_3_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__15097\,
            in1 => \N__15067\,
            in2 => \N__15091\,
            in3 => \N__18136\,
            lcout => \b2v_inst11.un34_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_3_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19575\,
            in2 => \_gnd_net_\,
            in3 => \N__15079\,
            lcout => \b2v_inst11.count_offZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34630\,
            ce => \N__18135\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_4_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__15058\,
            in1 => \_gnd_net_\,
            in2 => \N__19582\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34630\,
            ce => \N__18135\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_14_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15028\,
            in3 => \N__19579\,
            lcout => \b2v_inst11.count_off_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34630\,
            ce => \N__18135\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIA265A_14_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__19574\,
            in1 => \N__18134\,
            in2 => \N__15037\,
            in3 => \N__15024\,
            lcout => \b2v_inst11.count_offZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_7_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15289\,
            lcout => \b2v_inst16.count_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34647\,
            ce => \N__30623\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_4_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15271\,
            lcout => \b2v_inst16.count_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34647\,
            ce => \N__30623\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_1_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15222\,
            in2 => \_gnd_net_\,
            in3 => \N__15377\,
            lcout => \b2v_inst16.count_rst_6\,
            ltout => \b2v_inst16.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI2J651_0_1_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15204\,
            in2 => \N__15253\,
            in3 => \N__30609\,
            lcout => \b2v_inst16.un4_count_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI2J651_1_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__15205\,
            in1 => \_gnd_net_\,
            in2 => \N__30643\,
            in3 => \N__15250\,
            lcout => OPEN,
            ltout => \b2v_inst16.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIL9G52_1_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__15244\,
            in1 => \N__30199\,
            in2 => \N__15229\,
            in3 => \N__30151\,
            lcout => \b2v_inst16.un13_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_1_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15221\,
            in2 => \_gnd_net_\,
            in3 => \N__15379\,
            lcout => \b2v_inst16.count_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34640\,
            ce => \N__30639\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_10_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15196\,
            in1 => \N__17320\,
            in2 => \N__15175\,
            in3 => \N__15154\,
            lcout => OPEN,
            ltout => \b2v_inst16.un13_clk_100khz_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIL9G52_0_1_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__15139\,
            in1 => \N__15133\,
            in2 => \N__15127\,
            in3 => \N__15352\,
            lcout => \b2v_inst16.un13_clk_100khz_i\,
            ltout => \b2v_inst16.un13_clk_100khz_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_0_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__15378\,
            in1 => \_gnd_net_\,
            in2 => \N__15415\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34640\,
            ce => \N__30639\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_13_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15397\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34632\,
            ce => \N__30598\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_0_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__20339\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15382\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI1I651_0_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15412\,
            in2 => \N__15406\,
            in3 => \N__30571\,
            lcout => \b2v_inst16.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIHM041_13_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30572\,
            in1 => \N__15403\,
            in2 => \_gnd_net_\,
            in3 => \N__15396\,
            lcout => \b2v_inst16.countZ0Z_13\,
            ltout => \b2v_inst16.countZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_15_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15381\,
            in1 => \N__15301\,
            in2 => \N__15355\,
            in3 => \N__15345\,
            lcout => \b2v_inst16.un13_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNILS241_15_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30574\,
            in1 => \N__15325\,
            in2 => \_gnd_net_\,
            in3 => \N__15333\,
            lcout => \b2v_inst16.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_15_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15334\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34632\,
            ce => \N__30598\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIJP141_14_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30573\,
            in1 => \N__15319\,
            in2 => \_gnd_net_\,
            in3 => \N__15312\,
            lcout => \b2v_inst16.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_15_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16051\,
            lcout => \b2v_inst200.count_2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34628\,
            ce => \N__15661\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_2_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15550\,
            lcout => \b2v_inst200.count_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34628\,
            ce => \N__15661\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_7_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15910\,
            lcout => \b2v_inst200.count_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34628\,
            ce => \N__15661\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_17_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__16026\,
            in1 => \N__15562\,
            in2 => \N__15589\,
            in3 => \N__15996\,
            lcout => \b2v_inst200.un25_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIB9S71_16_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15427\,
            in1 => \N__16015\,
            in2 => \_gnd_net_\,
            in3 => \N__15707\,
            lcout => \b2v_inst200.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_16_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16014\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34623\,
            ce => \N__15660\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIDCT71_17_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15421\,
            in1 => \N__15981\,
            in2 => \_gnd_net_\,
            in3 => \N__15705\,
            lcout => \b2v_inst200.countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_17_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15982\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34623\,
            ce => \N__15660\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIP16E1_1_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15733\,
            in1 => \N__15573\,
            in2 => \_gnd_net_\,
            in3 => \N__15706\,
            lcout => \b2v_inst200.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_1_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15574\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34623\,
            ce => \N__15660\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI1QV41_2_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15727\,
            in1 => \N__15549\,
            in2 => \_gnd_net_\,
            in3 => \N__15704\,
            lcout => \b2v_inst200.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIC03N_0_0_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15606\,
            in2 => \_gnd_net_\,
            in3 => \N__33585\,
            lcout => \b2v_inst200.count_1_0\,
            ltout => OPEN,
            carryin => \bfn_2_6_0_\,
            carryout => \b2v_inst200.un2_count_1_cry_1_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIC03N_5_0_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15585\,
            in2 => \_gnd_net_\,
            in3 => \N__15565\,
            lcout => \b2v_inst200.count_RNIC03N_5Z0Z_0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_1_cy\,
            carryout => \b2v_inst200.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15561\,
            in2 => \_gnd_net_\,
            in3 => \N__15535\,
            lcout => \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_1\,
            carryout => \b2v_inst200.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15531\,
            in2 => \_gnd_net_\,
            in3 => \N__15511\,
            lcout => \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_2\,
            carryout => \b2v_inst200.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15504\,
            in2 => \_gnd_net_\,
            in3 => \N__15484\,
            lcout => \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_3\,
            carryout => \b2v_inst200.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15480\,
            in2 => \_gnd_net_\,
            in3 => \N__15460\,
            lcout => \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_4\,
            carryout => \b2v_inst200.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15952\,
            in3 => \N__15925\,
            lcout => \b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_5\,
            carryout => \b2v_inst200.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15921\,
            in2 => \_gnd_net_\,
            in3 => \N__15895\,
            lcout => \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_6\,
            carryout => \b2v_inst200.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15892\,
            in2 => \_gnd_net_\,
            in3 => \N__15868\,
            lcout => \b2v_inst200.un2_count_1_cry_7_c_RNIP33EZ0\,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => \b2v_inst200.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15865\,
            in2 => \_gnd_net_\,
            in3 => \N__15850\,
            lcout => \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_8\,
            carryout => \b2v_inst200.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15847\,
            in2 => \_gnd_net_\,
            in3 => \N__15817\,
            lcout => \b2v_inst200.un2_count_1_cry_9_c_RNIR75EZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_9\,
            carryout => \b2v_inst200.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15814\,
            in2 => \_gnd_net_\,
            in3 => \N__15784\,
            lcout => \b2v_inst200.un2_count_1_cry_10_c_RNI3AZ0Z29\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_10\,
            carryout => \b2v_inst200.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15780\,
            in2 => \_gnd_net_\,
            in3 => \N__15760\,
            lcout => \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_11\,
            carryout => \b2v_inst200.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15756\,
            in2 => \_gnd_net_\,
            in3 => \N__15736\,
            lcout => \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_12\,
            carryout => \b2v_inst200.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16086\,
            in2 => \_gnd_net_\,
            in3 => \N__16066\,
            lcout => \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_13\,
            carryout => \b2v_inst200.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_14_c_RNI7I69_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16062\,
            in2 => \_gnd_net_\,
            in3 => \N__16036\,
            lcout => \b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_14\,
            carryout => \b2v_inst200.un2_count_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__33608\,
            in1 => \N__16033\,
            in2 => \_gnd_net_\,
            in3 => \N__16003\,
            lcout => \b2v_inst200.count_1_16\,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => \b2v_inst200.un2_count_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__16000\,
            in1 => \N__33609\,
            in2 => \_gnd_net_\,
            in3 => \N__15985\,
            lcout => \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIQRSE5_11_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__15961\,
            in1 => \N__16610\,
            in2 => \N__17499\,
            in3 => \N__15969\,
            lcout => \b2v_inst11.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_10_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__16613\,
            in1 => \N__16201\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34608\,
            ce => \N__17511\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_11_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16612\,
            in2 => \_gnd_net_\,
            in3 => \N__15970\,
            lcout => \b2v_inst11.count_clk_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34608\,
            ce => \N__17511\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIS1M95_0_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16450\,
            in1 => \N__16213\,
            in2 => \_gnd_net_\,
            in3 => \N__17466\,
            lcout => \b2v_inst11.count_clkZ0Z_0\,
            ltout => \b2v_inst11.count_clkZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_0_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15955\,
            in3 => \N__16611\,
            lcout => \b2v_inst11.count_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34608\,
            ce => \N__17511\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIHFHA5_10_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__16207\,
            in1 => \N__17467\,
            in2 => \N__16617\,
            in3 => \N__16200\,
            lcout => \b2v_inst11.count_clkZ0Z_10\,
            ltout => \b2v_inst11.count_clkZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_15_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16488\,
            in1 => \N__16182\,
            in2 => \N__16168\,
            in3 => \N__16165\,
            lcout => OPEN,
            ltout => \b2v_inst11.un2_count_clk_17_0_o2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_13_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16431\,
            in1 => \N__16146\,
            in2 => \N__16150\,
            in3 => \N__16116\,
            lcout => \b2v_inst11.N_172\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI050F5_14_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17485\,
            in1 => \N__16093\,
            in2 => \_gnd_net_\,
            in3 => \N__16101\,
            lcout => \b2v_inst11.count_clkZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_13_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16126\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34612\,
            ce => \N__17527\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIU1VE5_13_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17484\,
            in1 => \N__16132\,
            in2 => \_gnd_net_\,
            in3 => \N__16125\,
            lcout => \b2v_inst11.count_clkZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_14_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16102\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34612\,
            ce => \N__17527\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIR4RV4_1_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__22846\,
            in1 => \N__27587\,
            in2 => \N__16498\,
            in3 => \N__17929\,
            lcout => \b2v_inst11.count_clk_en\,
            ltout => \b2v_inst11.count_clk_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIQ9CF5_2_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__16366\,
            in1 => \_gnd_net_\,
            in2 => \N__16369\,
            in3 => \N__16357\,
            lcout => \b2v_inst11.count_clkZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_2_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16365\,
            lcout => \b2v_inst11.count_clk_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34612\,
            ce => \N__17527\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNISCDF5_3_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17554\,
            in2 => \N__17500\,
            in3 => \N__17565\,
            lcout => \b2v_inst11.count_clkZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_7_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__16233\,
            in1 => \N__16348\,
            in2 => \_gnd_net_\,
            in3 => \N__16377\,
            lcout => \b2v_inst11.N_421\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_3_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16313\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16255\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_2_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__16334\,
            in1 => \N__16289\,
            in2 => \N__16351\,
            in3 => \N__16269\,
            lcout => \b2v_inst11.N_373\,
            ltout => \b2v_inst11.N_373_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_5_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16397\,
            in2 => \N__16342\,
            in3 => \N__16232\,
            lcout => \b2v_inst11.count_clk_RNIZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_2_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__16335\,
            in1 => \N__16314\,
            in2 => \N__16296\,
            in3 => \N__16268\,
            lcout => OPEN,
            ltout => \b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_3_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__16378\,
            in1 => \N__16254\,
            in2 => \N__16240\,
            in3 => \N__16231\,
            lcout => \b2v_inst11.count_clk_RNIZ0Z_3\,
            ltout => \b2v_inst11.count_clk_RNIZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNINJ641_3_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27318\,
            in2 => \N__16501\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un1_clk_100khz_32_and_i_o2_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIOEM52_1_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100011111100"
        )
    port map (
            in0 => \N__27317\,
            in1 => \N__29672\,
            in2 => \N__28751\,
            in3 => \N__22238\,
            lcout => \b2v_inst11.count_clk_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNISUTE5_12_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__17495\,
            in1 => \N__16456\,
            in2 => \N__16599\,
            in3 => \N__16467\,
            lcout => \b2v_inst11.count_clkZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_12_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16471\,
            in3 => \N__16565\,
            lcout => \b2v_inst11.count_clk_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34618\,
            ce => \N__17538\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_1_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__16691\,
            in1 => \N__16440\,
            in2 => \_gnd_net_\,
            in3 => \N__16543\,
            lcout => \b2v_inst11.count_clk_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34618\,
            ce => \N__17538\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_0_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__16439\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16564\,
            lcout => \b2v_inst11.count_clk_RNI_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__16692\,
            in1 => \N__16441\,
            in2 => \_gnd_net_\,
            in3 => \N__16542\,
            lcout => OPEN,
            ltout => \b2v_inst11.count_clk_RNIZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIT2M95_1_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16414\,
            in2 => \N__16408\,
            in3 => \N__17494\,
            lcout => \b2v_inst11.count_clkZ0Z_1\,
            ltout => \b2v_inst11.count_clkZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_1_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__16663\,
            in1 => \N__16713\,
            in2 => \N__16405\,
            in3 => \N__16398\,
            lcout => \b2v_inst11.N_187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_1_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__16712\,
            in1 => \N__16690\,
            in2 => \N__16672\,
            in3 => \N__16662\,
            lcout => \b2v_inst11.count_clk_RNI_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIF6NL_0_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29365\,
            in1 => \N__28459\,
            in2 => \N__23131\,
            in3 => \N__23342\,
            lcout => \b2v_inst11.N_328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIF6NL_0_0_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__23341\,
            in1 => \N__29364\,
            in2 => \N__16651\,
            in3 => \N__23127\,
            lcout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIVU5C_1_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24868\,
            in1 => \N__28572\,
            in2 => \N__19637\,
            in3 => \N__23340\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIE5T11_1_1_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__21597\,
            in1 => \N__29363\,
            in2 => \N__16630\,
            in3 => \N__28096\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNICC5V2_1_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__16627\,
            in1 => \N__22929\,
            in2 => \N__16621\,
            in3 => \N__28457\,
            lcout => \b2v_inst11.func_state_RNICC5V2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIF0H71_1_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__28458\,
            in1 => \_gnd_net_\,
            in2 => \N__22933\,
            in3 => \N__23343\,
            lcout => \b2v_inst11.N_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_10_c_RNI2O8H2_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19568\,
            in2 => \_gnd_net_\,
            in3 => \N__16824\,
            lcout => \b2v_inst11.count_off_1_11\,
            ltout => \b2v_inst11.count_off_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI4P25A_11_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16770\,
            in2 => \N__16513\,
            in3 => \N__18100\,
            lcout => \b2v_inst11.un3_count_off_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_11_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19571\,
            in2 => \_gnd_net_\,
            in3 => \N__16825\,
            lcout => \b2v_inst11.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34627\,
            ce => \N__18151\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIIP81A_0_9_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000111"
        )
    port map (
            in0 => \N__16723\,
            in1 => \N__18102\,
            in2 => \N__16963\,
            in3 => \N__17799\,
            lcout => OPEN,
            ltout => \b2v_inst11.un34_clk_100khz_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIQ1RAS1_9_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16816\,
            in1 => \N__16759\,
            in2 => \N__16810\,
            in3 => \N__16834\,
            lcout => \b2v_inst11.count_off_RNIQ1RAS1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_12_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__19570\,
            in1 => \_gnd_net_\,
            in2 => \N__16798\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34627\,
            ce => \N__18151\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI6S35A_12_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__18101\,
            in1 => \N__19569\,
            in2 => \N__16807\,
            in3 => \N__16794\,
            lcout => \b2v_inst11.count_offZ0Z_12\,
            ltout => \b2v_inst11.count_offZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI4P25A_0_11_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__16777\,
            in1 => \N__16771\,
            in2 => \N__16762\,
            in3 => \N__18152\,
            lcout => \b2v_inst11.un34_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_6_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19519\,
            in2 => \_gnd_net_\,
            in3 => \N__16939\,
            lcout => \b2v_inst11.count_offZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34631\,
            ce => \N__18156\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_9_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__19518\,
            in1 => \_gnd_net_\,
            in2 => \N__16735\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_offZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34631\,
            ce => \N__18156\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_8_c_RNIP80E2_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19517\,
            in2 => \_gnd_net_\,
            in3 => \N__16731\,
            lcout => \b2v_inst11.count_off_1_9\,
            ltout => \b2v_inst11.count_off_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIIP81A_9_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18143\,
            in1 => \_gnd_net_\,
            in2 => \N__16966\,
            in3 => \N__16962\,
            lcout => \b2v_inst11.un3_count_off_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_5_c_RNIM2TD2_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19515\,
            in2 => \_gnd_net_\,
            in3 => \N__16938\,
            lcout => \b2v_inst11.count_off_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_7_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19563\,
            in3 => \N__16906\,
            lcout => \b2v_inst11.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34631\,
            ce => \N__18156\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_6_c_RNIN4UD2_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19516\,
            in2 => \_gnd_net_\,
            in3 => \N__16905\,
            lcout => \b2v_inst11.count_off_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI01TT1_7_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__27034\,
            in1 => \N__26234\,
            in2 => \_gnd_net_\,
            in3 => \N__26253\,
            lcout => \b2v_inst11.dutycycle_RNI01TT1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_15_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19566\,
            in2 => \_gnd_net_\,
            in3 => \N__16887\,
            lcout => \b2v_inst11.count_off_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34639\,
            ce => \N__18158\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIC575A_15_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__19567\,
            in1 => \N__16894\,
            in2 => \N__18163\,
            in3 => \N__16888\,
            lcout => \b2v_inst11.count_offZ0Z_15\,
            ltout => \b2v_inst11.count_offZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_15_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16869\,
            in1 => \N__16855\,
            in2 => \N__16837\,
            in3 => \N__17862\,
            lcout => \b2v_inst11.un34_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_8_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__19565\,
            in1 => \_gnd_net_\,
            in2 => \N__17053\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34639\,
            ce => \N__18158\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIGM71A_8_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__17059\,
            in1 => \N__19564\,
            in2 => \N__18157\,
            in3 => \N__17049\,
            lcout => \b2v_inst11.count_offZ0Z_8\,
            ltout => \b2v_inst11.count_offZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIEJ61A_0_7_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000111"
        )
    port map (
            in0 => \N__18162\,
            in1 => \N__17002\,
            in2 => \N__17026\,
            in3 => \N__17011\,
            lcout => \b2v_inst11.un34_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIEJ61A_7_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17010\,
            in1 => \N__18139\,
            in2 => \_gnd_net_\,
            in3 => \N__17001\,
            lcout => \b2v_inst11.un3_count_off_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18790\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_1_0_\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18327\,
            in2 => \N__20191\,
            in3 => \N__16978\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17110\,
            in2 => \N__18331\,
            in3 => \N__16975\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17954\,
            in2 => \N__17101\,
            in3 => \N__16972\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17089\,
            in2 => \N__17959\,
            in3 => \N__16969\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__19999\,
            in1 => \N__18326\,
            in2 => \N__17080\,
            in3 => \N__17119\,
            lcout => \b2v_inst11.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17068\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17116\,
            lcout => \b2v_inst11.mult1_un96_sum_s_8\,
            ltout => \b2v_inst11.mult1_un96_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17113\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20212\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_2_0_\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17183\,
            in2 => \N__18385\,
            in3 => \N__17104\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17173\,
            in2 => \N__17188\,
            in3 => \N__17092\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21824\,
            in2 => \N__17164\,
            in3 => \N__17083\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17152\,
            in2 => \N__21831\,
            in3 => \N__17071\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17952\,
            in1 => \N__17187\,
            in2 => \N__17143\,
            in3 => \N__17062\,
            lcout => \b2v_inst11.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17131\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17191\,
            lcout => \b2v_inst11.mult1_un89_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21823\,
            lcout => \b2v_inst11.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18766\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_3_0_\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17201\,
            in2 => \N__18376\,
            in3 => \N__17167\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17263\,
            in2 => \N__17206\,
            in3 => \N__17155\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20069\,
            in2 => \N__17254\,
            in3 => \N__17146\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17242\,
            in2 => \N__20076\,
            in3 => \N__17134\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__21822\,
            in1 => \N__17205\,
            in2 => \N__17233\,
            in3 => \N__17125\,
            lcout => \b2v_inst11.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__17221\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17122\,
            lcout => \b2v_inst11.mult1_un82_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17953\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un85_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18745\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_4_0_\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18404\,
            in2 => \N__19897\,
            in3 => \N__17257\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18466\,
            in2 => \N__18409\,
            in3 => \N__17245\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20384\,
            in2 => \N__18457\,
            in3 => \N__17236\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18445\,
            in2 => \N__20389\,
            in3 => \N__17224\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20068\,
            in1 => \N__18408\,
            in2 => \N__18436\,
            in3 => \N__17215\,
            lcout => \b2v_inst11.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18424\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17212\,
            lcout => \b2v_inst11.mult1_un75_sum_s_8\,
            ltout => \b2v_inst11.mult1_un75_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17209\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18934\,
            in2 => \N__18865\,
            in3 => \N__18898\,
            lcout => \b2v_inst11.mult1_un40_sum_i_5\,
            ltout => \b2v_inst11.mult1_un40_sum_i_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17323\,
            in3 => \N__18633\,
            lcout => \b2v_inst11.mult1_un47_sum_s_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI4M8F1_10_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17281\,
            in1 => \N__17295\,
            in2 => \_gnd_net_\,
            in3 => \N__30567\,
            lcout => \b2v_inst16.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_10_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17296\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34634\,
            ce => \N__30605\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18955\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_6_0_\,
            carryout => \b2v_inst11.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17350\,
            in3 => \N__17275\,
            lcout => \b2v_inst11.mult1_un47_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un47_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17332\,
            in3 => \N__17272\,
            lcout => \b2v_inst11.mult1_un47_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un47_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20118\,
            in2 => \N__17341\,
            in3 => \N__17269\,
            lcout => \b2v_inst11.mult1_un47_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un47_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17266\,
            lcout => \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__18500\,
            in1 => \N__18501\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un47_sum_l_fx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__18671\,
            in1 => \N__18672\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un47_sum_l_fx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_en_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33717\,
            in2 => \_gnd_net_\,
            in3 => \N__33082\,
            lcout => \b2v_inst200.count_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18925\,
            lcout => \b2v_inst11.un1_dutycycle_53_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000101"
        )
    port map (
            in0 => \N__18927\,
            in1 => \_gnd_net_\,
            in2 => \N__18897\,
            in3 => \N__18858\,
            lcout => \b2v_inst11.mult1_un40_sum_i_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18951\,
            lcout => \b2v_inst11.mult1_un47_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__18926\,
            in1 => \_gnd_net_\,
            in2 => \N__18896\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un47_sum_s_4_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18783\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNI_0_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30403\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.N_2925_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_3_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17572\,
            lcout => \b2v_inst11.count_clk_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34620\,
            ce => \N__17526\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI3JFN6_13_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100000000"
        )
    port map (
            in0 => \N__27759\,
            in1 => \N__22253\,
            in2 => \N__17401\,
            in3 => \N__27596\,
            lcout => \b2v_inst11.dutycycle_en_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIAI7C4_13_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__21313\,
            in1 => \N__22586\,
            in2 => \_gnd_net_\,
            in3 => \N__22396\,
            lcout => \b2v_inst11.N_150_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIAI7C4_14_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__22587\,
            in1 => \_gnd_net_\,
            in2 => \N__22402\,
            in3 => \N__21244\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_152_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI3JFN6_14_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010101010"
        )
    port map (
            in0 => \N__27597\,
            in1 => \N__22255\,
            in2 => \N__17392\,
            in3 => \N__27760\,
            lcout => \b2v_inst11.dutycycle_en_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI4UUA8_15_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__27292\,
            in1 => \N__17373\,
            in2 => \N__21106\,
            in3 => \N__17383\,
            lcout => \b2v_inst11.dutycycleZ0Z_12\,
            ltout => \b2v_inst11.dutycycleZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIAI7C4_15_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22588\,
            in2 => \N__17389\,
            in3 => \N__22400\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_155_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI3JFN6_15_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100000000"
        )
    port map (
            in0 => \N__27758\,
            in1 => \N__22254\,
            in2 => \N__17386\,
            in3 => \N__27595\,
            lcout => \b2v_inst11.dutycycle_en_12\,
            ltout => \b2v_inst11.dutycycle_en_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_15_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__21105\,
            in1 => \N__17374\,
            in2 => \N__17377\,
            in3 => \N__27316\,
            lcout => \b2v_inst11.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34613\,
            ce => 'H',
            sr => \N__24232\
        );

    \b2v_inst11.dutycycle_13_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__17605\,
            in1 => \N__21265\,
            in2 => \N__17596\,
            in3 => \N__27315\,
            lcout => \b2v_inst11.dutycycleZ1Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34619\,
            ce => 'H',
            sr => \N__24227\
        );

    \b2v_inst11.dutycycle_RNI_2_12_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__21434\,
            in1 => \N__19339\,
            in2 => \_gnd_net_\,
            in3 => \N__22359\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_2Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_10_9_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__19340\,
            in1 => \N__19011\,
            in2 => \N__17611\,
            in3 => \N__21014\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_10Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_13_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21246\,
            in2 => \N__17608\,
            in3 => \N__21306\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI0OSA8_13_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__17604\,
            in1 => \N__21264\,
            in2 => \N__17595\,
            in3 => \N__27314\,
            lcout => \b2v_inst11.dutycycleZ0Z_9\,
            ltout => \b2v_inst11.dutycycleZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_13_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__21433\,
            in1 => \_gnd_net_\,
            in2 => \N__17581\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_0Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_10_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001011"
        )
    port map (
            in0 => \N__22360\,
            in1 => \N__19345\,
            in2 => \N__17578\,
            in3 => \N__19177\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_10\,
            ltout => \b2v_inst11.dutycycle_RNI_1Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_14_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17575\,
            in3 => \N__21245\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIHTFQ_8_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__17672\,
            in1 => \N__26954\,
            in2 => \_gnd_net_\,
            in3 => \N__26879\,
            lcout => \b2v_inst11.dutycycle_RNIHTFQZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIJU083_8_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001100"
        )
    port map (
            in0 => \N__22593\,
            in1 => \N__28117\,
            in2 => \N__22783\,
            in3 => \N__22240\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNIJU083Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNITG8K7_8_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__27312\,
            in1 => \_gnd_net_\,
            in2 => \N__17695\,
            in3 => \N__17647\,
            lcout => \b2v_inst11.N_108_f0\,
            ltout => \b2v_inst11.N_108_f0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_8_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__17680\,
            in1 => \N__27780\,
            in2 => \N__17692\,
            in3 => \N__17674\,
            lcout => \b2v_inst11.dutycycleZ1Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34624\,
            ce => 'H',
            sr => \N__24231\
        );

    \b2v_inst11.dutycycle_RNI2NK31_8_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__17673\,
            in1 => \N__26955\,
            in2 => \N__21034\,
            in3 => \N__26880\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI2NK31Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIA8B23_8_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17689\,
            in2 => \N__17683\,
            in3 => \N__27313\,
            lcout => \b2v_inst11.dutycycle_e_1_8\,
            ltout => \b2v_inst11.dutycycle_e_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI9QKHC_8_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__17671\,
            in1 => \N__17659\,
            in2 => \N__17653\,
            in3 => \N__27778\,
            lcout => \b2v_inst11.dutycycleZ0Z_1\,
            ltout => \b2v_inst11.dutycycleZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIJU083_0_8_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22592\,
            in2 => \N__17650\,
            in3 => \N__22239\,
            lcout => \b2v_inst11.dutycycle_RNIJU083_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_RNIM6F44_0_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33778\,
            lcout => \delayed_vccin_vccinaux_ok_RNIM6F44_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_9_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21013\,
            in2 => \_gnd_net_\,
            in3 => \N__22361\,
            lcout => \b2v_inst11.un1_dutycycle_53_41_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_12_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21417\,
            in1 => \N__19337\,
            in2 => \N__24382\,
            in3 => \N__19432\,
            lcout => \b2v_inst11.g0_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_1_1_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28455\,
            lcout => \b2v_inst11.func_state_RNI_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIT4D71_1_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__28456\,
            in1 => \N__17986\,
            in2 => \N__29362\,
            in3 => \N__26964\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_289_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIFIVO1_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__28292\,
            in1 => \N__20776\,
            in2 => \N__17707\,
            in3 => \N__21591\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_1_0_iv_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI666T2_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111111"
        )
    port map (
            in0 => \N__28291\,
            in1 => \N__28708\,
            in2 => \N__17704\,
            in3 => \N__29099\,
            lcout => \b2v_inst11.N_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_12_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__19431\,
            in1 => \N__18580\,
            in2 => \N__19344\,
            in3 => \N__21416\,
            lcout => \b2v_inst11.m15_e_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_12_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__27296\,
            in1 => \N__17761\,
            in2 => \N__17755\,
            in3 => \N__21355\,
            lcout => \b2v_inst11.dutycycleZ1Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34633\,
            ce => 'H',
            sr => \N__24238\
        );

    \b2v_inst11.dutycycle_RNINJ641_11_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19318\,
            in2 => \_gnd_net_\,
            in3 => \N__27294\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_302_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIGKEF3_11_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100000000"
        )
    port map (
            in0 => \N__27779\,
            in1 => \N__17734\,
            in2 => \N__17701\,
            in3 => \N__27599\,
            lcout => \b2v_inst11.dutycycle_RNIGKEF3Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNINJ641_12_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27295\,
            in2 => \_gnd_net_\,
            in3 => \N__21415\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIGKEF3_12_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101010"
        )
    port map (
            in0 => \N__27598\,
            in1 => \N__27777\,
            in2 => \N__17698\,
            in3 => \N__17733\,
            lcout => \b2v_inst11.dutycycle_RNIGKEF3Z0Z_12\,
            ltout => \b2v_inst11.dutycycle_RNIGKEF3Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIBMQ25_12_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__21354\,
            in1 => \N__17751\,
            in2 => \N__17743\,
            in3 => \N__27293\,
            lcout => \b2v_inst11.dutycycleZ0Z_10\,
            ltout => \b2v_inst11.dutycycleZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_12_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__19319\,
            in1 => \_gnd_net_\,
            in2 => \N__17740\,
            in3 => \N__19015\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_56_a0_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_13_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010000"
        )
    port map (
            in0 => \N__19084\,
            in1 => \N__21335\,
            in2 => \N__17737\,
            in3 => \N__19246\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIAI7C4_2_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110001111"
        )
    port map (
            in0 => \N__19357\,
            in1 => \N__27304\,
            in2 => \N__22603\,
            in3 => \N__19402\,
            lcout => \b2v_inst11.N_232_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_1_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23375\,
            in1 => \N__29112\,
            in2 => \N__23286\,
            in3 => \N__29236\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_func_state25_6_0_o_N_325_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__17719\,
            in1 => \N__28462\,
            in2 => \N__17725\,
            in3 => \N__19605\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_func_state25_6_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_en_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__27619\,
            in1 => \N__21505\,
            in2 => \N__17722\,
            in3 => \N__17713\,
            lcout => \b2v_inst11.count_off_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__25086\,
            in1 => \N__28461\,
            in2 => \N__19396\,
            in3 => \N__23374\,
            lcout => \b2v_inst11.un1_func_state25_6_0_o_N_323_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_0_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22875\,
            in1 => \N__29111\,
            in2 => \N__23285\,
            in3 => \N__19641\,
            lcout => \b2v_inst11.un1_func_state25_6_0_o_N_324_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINJ641_1_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__23054\,
            in1 => \N__28460\,
            in2 => \N__23382\,
            in3 => \N__24313\,
            lcout => \b2v_inst11.N_322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI51SU9_1_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__17869\,
            in1 => \N__19468\,
            in2 => \N__18077\,
            in3 => \N__17878\,
            lcout => \b2v_inst11.count_offZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI40SU9_0_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__19467\,
            in1 => \N__17827\,
            in2 => \N__17852\,
            in3 => \N__18033\,
            lcout => \b2v_inst11.count_offZ0Z_0\,
            ltout => \b2v_inst11.count_offZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_1_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17914\,
            in3 => \N__17897\,
            lcout => \b2v_inst11.count_off_RNIZ0Z_1\,
            ltout => \b2v_inst11.count_off_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_1_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__19471\,
            in1 => \_gnd_net_\,
            in2 => \N__17872\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34648\,
            ce => \N__18037\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_0_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17845\,
            in2 => \_gnd_net_\,
            in3 => \N__19472\,
            lcout => \b2v_inst11.count_off_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34648\,
            ce => \N__18037\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_10_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17811\,
            lcout => \b2v_inst11.count_off_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34648\,
            ce => \N__18037\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIRAR1A_10_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__18038\,
            in1 => \N__17821\,
            in2 => \N__17815\,
            in3 => \N__19466\,
            lcout => \b2v_inst11.count_offZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_13_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19470\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17776\,
            lcout => \b2v_inst11.count_off_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34648\,
            ce => \N__18037\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIVU5C_0_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28488\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24316\,
            lcout => \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18826\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_1_0_\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18185\,
            in2 => \N__18367\,
            in3 => \N__17977\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18298\,
            in2 => \N__18190\,
            in3 => \N__17974\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18351\,
            in2 => \N__18283\,
            in3 => \N__17971\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18262\,
            in2 => \N__18355\,
            in3 => \N__17968\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20148\,
            in1 => \N__18189\,
            in2 => \N__18247\,
            in3 => \N__17965\,
            lcout => \b2v_inst11.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18211\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17962\,
            lcout => \b2v_inst11.mult1_un110_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17958\,
            lcout => \b2v_inst11.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18808\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_2_0_\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18230\,
            in2 => \N__18316\,
            in3 => \N__18292\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18289\,
            in2 => \N__18235\,
            in3 => \N__18274\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20000\,
            in2 => \N__18271\,
            in3 => \N__18256\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18253\,
            in2 => \N__20007\,
            in3 => \N__18238\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18349\,
            in1 => \N__18234\,
            in2 => \N__18220\,
            in3 => \N__18205\,
            lcout => \b2v_inst11.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18202\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18196\,
            lcout => \b2v_inst11.mult1_un103_sum_s_8\,
            ltout => \b2v_inst11.mult1_un103_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18193\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19728\,
            in2 => \_gnd_net_\,
            in3 => \N__20272\,
            lcout => \b2v_inst11.mult1_un131_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18825\,
            lcout => \b2v_inst11.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20271\,
            lcout => \b2v_inst11.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20273\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19944\,
            lcout => \b2v_inst11.mult1_un131_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18762\,
            lcout => \b2v_inst11.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18741\,
            lcout => \b2v_inst11.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18807\,
            lcout => \b2v_inst11.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18350\,
            lcout => \b2v_inst11.un85_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19914\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_4_0_\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_2_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20171\,
            in2 => \N__20398\,
            in3 => \N__18460\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_2_c\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_3_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18394\,
            in2 => \N__20176\,
            in3 => \N__18448\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_3_c\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_4_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18562\,
            in2 => \N__20050\,
            in3 => \N__18439\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_4_c\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_5_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18553\,
            in2 => \N__20049\,
            in3 => \N__18427\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_5_c\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_6_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20383\,
            in1 => \N__20175\,
            in2 => \N__18544\,
            in3 => \N__18418\,
            lcout => \b2v_inst11.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_6_c\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18532\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18415\,
            lcout => \b2v_inst11.mult1_un68_sum_s_8\,
            ltout => \b2v_inst11.mult1_un68_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18412\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20415\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_5_0_\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20422\,
            in2 => \N__18597\,
            in3 => \N__18388\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18593\,
            in2 => \N__18514\,
            in3 => \N__18556\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18475\,
            in2 => \N__18619\,
            in3 => \N__18547\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18618\,
            in2 => \N__18712\,
            in3 => \N__18535\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20038\,
            in1 => \N__18691\,
            in2 => \N__18598\,
            in3 => \N__18526\,
            lcout => \b2v_inst11.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18655\,
            in3 => \N__18523\,
            lcout => \b2v_inst11.mult1_un61_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20443\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_6_0_\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18520\,
            in2 => \_gnd_net_\,
            in3 => \N__18505\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18502\,
            in2 => \N__18484\,
            in3 => \N__18469\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20096\,
            in2 => \N__18721\,
            in3 => \N__18703\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20114\,
            in2 => \N__18700\,
            in3 => \N__18685\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18614\,
            in1 => \N__18682\,
            in2 => \N__18676\,
            in3 => \N__18646\,
            lcout => \b2v_inst11.mult1_un61_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18643\,
            in2 => \N__18637\,
            in3 => \N__18622\,
            lcout => \b2v_inst11.mult1_un54_sum_s_8\,
            ltout => \b2v_inst11.mult1_un54_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18601\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24819\,
            in2 => \N__25597\,
            in3 => \N__25385\,
            lcout => \b2v_inst11.m15_e_2\,
            ltout => OPEN,
            carryin => \bfn_5_7_0_\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_0_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25594\,
            in2 => \N__20521\,
            in3 => \N__18568\,
            lcout => \b2v_inst11.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_0_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27428\,
            in2 => \N__20464\,
            in3 => \N__18565\,
            lcout => \b2v_inst11.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_1_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23992\,
            in2 => \N__27435\,
            in3 => \N__18832\,
            lcout => \b2v_inst11.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_2_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22465\,
            in2 => \N__22453\,
            in3 => \N__18829\,
            lcout => \b2v_inst11.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_3_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_4_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26766\,
            in2 => \N__22483\,
            in3 => \N__18811\,
            lcout => \b2v_inst11.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_4_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20449\,
            in2 => \N__26779\,
            in3 => \N__18793\,
            lcout => \b2v_inst11.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_5_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20455\,
            in2 => \N__22363\,
            in3 => \N__18772\,
            lcout => \b2v_inst11.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_6_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20892\,
            in2 => \N__19096\,
            in3 => \N__18769\,
            lcout => \b2v_inst11.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21442\,
            in2 => \N__19192\,
            in3 => \N__18748\,
            lcout => \b2v_inst11.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_8_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_9_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21324\,
            in2 => \N__19060\,
            in3 => \N__18727\,
            lcout => \b2v_inst11.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_9_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21224\,
            in2 => \N__19036\,
            in3 => \N__18724\,
            lcout => \b2v_inst11.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_10\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21140\,
            in2 => \N__19027\,
            in3 => \N__18985\,
            lcout => \b2v_inst11.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_11\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21325\,
            in2 => \N__18982\,
            in3 => \N__18967\,
            lcout => \b2v_inst11.mult1_un54_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_12\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18964\,
            in2 => \N__21240\,
            in3 => \N__18937\,
            lcout => \b2v_inst11.mult1_un47_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_13\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18838\,
            in2 => \N__21154\,
            in3 => \N__18910\,
            lcout => \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_14\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21155\,
            in2 => \N__18907\,
            in3 => \N__18871\,
            lcout => \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \b2v_inst11.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.CO2_THRU_LUT4_0_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18868\,
            lcout => \b2v_inst11.CO2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_15_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__21149\,
            in1 => \N__21223\,
            in2 => \_gnd_net_\,
            in3 => \N__18844\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_9_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__26232\,
            in1 => \N__22779\,
            in2 => \N__22362\,
            in3 => \N__21011\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_44_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_9_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__21012\,
            in1 => \N__18991\,
            in2 => \N__19042\,
            in3 => \N__20659\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_6Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_11_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22354\,
            in1 => \N__21231\,
            in2 => \N__19039\,
            in3 => \N__20891\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_10_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22778\,
            in1 => \N__28972\,
            in2 => \N__28036\,
            in3 => \N__22350\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_15_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011001100"
        )
    port map (
            in0 => \N__21156\,
            in1 => \N__18997\,
            in2 => \N__19213\,
            in3 => \N__20647\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_7_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__26213\,
            in1 => \N__22728\,
            in2 => \_gnd_net_\,
            in3 => \N__19142\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_m7_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_4_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010110110101"
        )
    port map (
            in0 => \N__22729\,
            in1 => \N__28014\,
            in2 => \N__19018\,
            in3 => \N__28934\,
            lcout => \b2v_inst11.un1_i3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_11_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20890\,
            in2 => \_gnd_net_\,
            in3 => \N__21436\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_4_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__28016\,
            in1 => \N__28936\,
            in2 => \N__19154\,
            in3 => \N__19338\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_4_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__26215\,
            in1 => \N__22734\,
            in2 => \N__28973\,
            in3 => \N__28018\,
            lcout => \b2v_inst11.un1_dutycycle_53_44_0_2_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_4_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110101011"
        )
    port map (
            in0 => \N__19143\,
            in1 => \N__28935\,
            in2 => \N__22771\,
            in3 => \N__26214\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_39_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_9_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000001110"
        )
    port map (
            in0 => \N__20996\,
            in1 => \N__22733\,
            in2 => \N__19078\,
            in3 => \N__28017\,
            lcout => \b2v_inst11.un1_dutycycle_53_39_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__22414\,
            in1 => \N__22761\,
            in2 => \N__19155\,
            in3 => \N__20674\,
            lcout => \b2v_inst11.N_357\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_9_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111001111"
        )
    port map (
            in0 => \N__20592\,
            in1 => \N__22645\,
            in2 => \N__28032\,
            in3 => \N__20957\,
            lcout => \b2v_inst11.dutycycle_RNI_8Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNINJ641_9_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011111"
        )
    port map (
            in0 => \N__27305\,
            in1 => \N__28107\,
            in2 => \N__19156\,
            in3 => \N__22241\,
            lcout => \b2v_inst11.dutycycle_eena_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__22776\,
            in1 => \N__26189\,
            in2 => \N__28974\,
            in3 => \N__19150\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_39_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_13_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111000000"
        )
    port map (
            in0 => \N__21314\,
            in1 => \N__19075\,
            in2 => \N__19069\,
            in3 => \N__19066\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_9_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20956\,
            lcout => \b2v_inst11.dutycycle_RNI_5Z0Z_9\,
            ltout => \b2v_inst11.dutycycle_RNI_5Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_9_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110111"
        )
    port map (
            in0 => \N__20958\,
            in1 => \N__28940\,
            in2 => \N__19048\,
            in3 => \N__22775\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_10_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111010001100"
        )
    port map (
            in0 => \N__28024\,
            in1 => \N__26188\,
            in2 => \N__19045\,
            in3 => \N__22764\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNIZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_12_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__20959\,
            in1 => \N__22777\,
            in2 => \N__19195\,
            in3 => \N__21440\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_4_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28971\,
            in1 => \N__19162\,
            in2 => \_gnd_net_\,
            in3 => \N__19111\,
            lcout => OPEN,
            ltout => \b2v_inst11.m18_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_11_9_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__19168\,
            in1 => \N__20994\,
            in2 => \N__19180\,
            in3 => \N__28011\,
            lcout => \b2v_inst11.dutycycle_RNI_11Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_7_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__19141\,
            in1 => \N__26203\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_7_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101011101"
        )
    port map (
            in0 => \N__22725\,
            in1 => \N__19140\,
            in2 => \N__26230\,
            in3 => \N__28010\,
            lcout => \b2v_inst11.dutycycle_RNI_5Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_7_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__19139\,
            in1 => \N__26199\,
            in2 => \_gnd_net_\,
            in3 => \N__22726\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_7_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100101101010"
        )
    port map (
            in0 => \N__19201\,
            in1 => \N__19105\,
            in2 => \N__26231\,
            in3 => \N__28012\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_11_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19099\,
            in3 => \N__20880\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_9_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__22727\,
            in1 => \N__20995\,
            in2 => \N__22615\,
            in3 => \N__22348\,
            lcout => \b2v_inst11.un1_dutycycle_53_13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_11_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__20876\,
            in1 => \N__21409\,
            in2 => \_gnd_net_\,
            in3 => \N__22345\,
            lcout => \b2v_inst11.G_6_i_a4_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_11_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__19228\,
            in1 => \N__19239\,
            in2 => \N__21457\,
            in3 => \N__27303\,
            lcout => \b2v_inst11.dutycycleZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34641\,
            ce => 'H',
            sr => \N__24237\
        );

    \b2v_inst11.dutycycle_RNI_0_11_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100110101"
        )
    port map (
            in0 => \N__20875\,
            in1 => \N__19328\,
            in2 => \N__21441\,
            in3 => \N__22346\,
            lcout => OPEN,
            ltout => \b2v_inst11.G_6_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_9_9_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001111"
        )
    port map (
            in0 => \N__20998\,
            in1 => \N__19270\,
            in2 => \N__19255\,
            in3 => \N__19252\,
            lcout => \b2v_inst11.un1_dutycycle_53_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI9JP25_11_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__27302\,
            in1 => \N__21453\,
            in2 => \N__19240\,
            in3 => \N__19227\,
            lcout => \b2v_inst11.dutycycleZ0Z_7\,
            ltout => \b2v_inst11.dutycycleZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_11_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19219\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_11\,
            ltout => \b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_9_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100001100"
        )
    port map (
            in0 => \N__22774\,
            in1 => \N__20997\,
            in2 => \N__19216\,
            in3 => \N__22347\,
            lcout => \b2v_inst11.un1_dutycycle_53_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_11_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22773\,
            in2 => \_gnd_net_\,
            in3 => \N__20874\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_0_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__25571\,
            in1 => \N__25364\,
            in2 => \N__28028\,
            in3 => \N__24512\,
            lcout => \b2v_inst11.g2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_12_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__19333\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21394\,
            lcout => \b2v_inst11.N_354\,
            ltout => \b2v_inst11.N_354_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_2_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__27417\,
            in1 => \_gnd_net_\,
            in2 => \N__19348\,
            in3 => \N__19429\,
            lcout => \b2v_inst11.N_360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_2_1_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24511\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_3046_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_12_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__21395\,
            in1 => \N__19332\,
            in2 => \_gnd_net_\,
            in3 => \N__19430\,
            lcout => OPEN,
            ltout => \b2v_inst11.g3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_0_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111101"
        )
    port map (
            in0 => \N__19279\,
            in1 => \N__28832\,
            in2 => \N__19273\,
            in3 => \N__28141\,
            lcout => \b2v_inst11.g2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_4_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010011"
        )
    port map (
            in0 => \N__26219\,
            in1 => \N__22772\,
            in2 => \N__28996\,
            in3 => \N__27999\,
            lcout => \b2v_inst11.N_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNINJ641_0_5_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111111"
        )
    port map (
            in0 => \N__28829\,
            in1 => \N__19264\,
            in2 => \N__27322\,
            in3 => \N__24314\,
            lcout => \b2v_inst11.dutycycle_RNINJ641_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_5_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21492\,
            in2 => \_gnd_net_\,
            in3 => \N__23176\,
            lcout => \b2v_inst11.dutycycle_RNI_6Z0Z_5\,
            ltout => \b2v_inst11.dutycycle_RNI_6Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINJ641_2_1_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__29239\,
            in1 => \N__21073\,
            in2 => \N__19258\,
            in3 => \N__21600\,
            lcout => \b2v_inst11.func_state_1_m2s2_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_3_1_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21601\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24317\,
            lcout => \b2v_inst11.func_state_RNI_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIT4D71_1_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__28559\,
            in1 => \N__24092\,
            in2 => \N__23428\,
            in3 => \N__19642\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIKOJB2_0_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__22882\,
            in1 => \N__23242\,
            in2 => \N__19609\,
            in3 => \N__19606\,
            lcout => \b2v_inst11.N_122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__28668\,
            in1 => \N__28253\,
            in2 => \_gnd_net_\,
            in3 => \N__28560\,
            lcout => \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__21082\,
            in1 => \N__28142\,
            in2 => \N__27427\,
            in3 => \N__19428\,
            lcout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_0_0_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__28219\,
            in1 => \N__28549\,
            in2 => \_gnd_net_\,
            in3 => \N__24301\,
            lcout => \b2v_inst11.un1_func_state25_6_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIC5UE2_1_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101010"
        )
    port map (
            in0 => \N__19384\,
            in1 => \N__28548\,
            in2 => \N__24097\,
            in3 => \N__23376\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_1_m0_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIIVR84_0_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__23377\,
            in1 => \N__19372\,
            in2 => \N__19360\,
            in3 => \N__21475\,
            lcout => \b2v_inst11.func_state_1_m0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19858\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_1_0_\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19757\,
            in2 => \N__19714\,
            in3 => \N__19702\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19699\,
            in2 => \N__19762\,
            in3 => \N__19693\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20149\,
            in2 => \N__19690\,
            in3 => \N__19681\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19678\,
            in2 => \N__20157\,
            in3 => \N__19672\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__19876\,
            in1 => \N__19761\,
            in2 => \N__19669\,
            in3 => \N__19660\,
            lcout => \b2v_inst11.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19657\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19651\,
            lcout => \b2v_inst11.mult1_un117_sum_s_8\,
            ltout => \b2v_inst11.mult1_un117_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19648\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20236\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_2_0_\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19793\,
            in2 => \N__19840\,
            in3 => \N__19645\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19828\,
            in2 => \N__19798\,
            in3 => \N__19822\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19877\,
            in2 => \N__19819\,
            in3 => \N__19810\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19807\,
            in2 => \N__19884\,
            in3 => \N__19801\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20263\,
            in1 => \N__19797\,
            in2 => \N__19783\,
            in3 => \N__19774\,
            lcout => \b2v_inst11.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__19771\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19765\,
            lcout => \b2v_inst11.mult1_un124_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20153\,
            lcout => \b2v_inst11.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21744\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20218\,
            in2 => \N__19747\,
            in3 => \N__19738\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19735\,
            in2 => \N__19729\,
            in3 => \N__19981\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20264\,
            in2 => \N__19978\,
            in3 => \N__19966\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19963\,
            in2 => \N__20274\,
            in3 => \N__19957\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__21796\,
            in1 => \N__19954\,
            in2 => \N__19948\,
            in3 => \N__19930\,
            lcout => \b2v_inst11.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19927\,
            in2 => \_gnd_net_\,
            in3 => \N__19921\,
            lcout => \b2v_inst11.mult1_un131_sum_s_8\,
            ltout => \b2v_inst11.mult1_un131_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19918\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19915\,
            lcout => \b2v_inst11.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19885\,
            lcout => \b2v_inst11.un85_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19854\,
            lcout => \b2v_inst11.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20275\,
            lcout => \b2v_inst11.un85_clk_100khz_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20232\,
            lcout => \b2v_inst11.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20208\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20045\,
            lcout => \b2v_inst11.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20161\,
            lcout => \b2v_inst11.un85_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20080\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un85_clk_100khz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20037\,
            lcout => \b2v_inst11.mult1_un61_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20011\,
            lcout => \b2v_inst11.un85_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20442\,
            lcout => \b2v_inst11.mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20416\,
            lcout => \b2v_inst11.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20388\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un85_clk_100khz_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.delayed_vddq_pwrgd_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__20629\,
            in1 => \N__20543\,
            in2 => \_gnd_net_\,
            in3 => \N__25077\,
            lcout => \b2v_inst16.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34643\,
            ce => \N__33684\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIPRCE_1_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20540\,
            in1 => \N__20358\,
            in2 => \N__20305\,
            in3 => \N__34058\,
            lcout => \b2v_inst16.curr_stateZ0Z_1\,
            ltout => \b2v_inst16.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNI7SG01_1_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__20628\,
            in1 => \_gnd_net_\,
            in2 => \N__20365\,
            in3 => \N__25073\,
            lcout => OPEN,
            ltout => \b2v_inst16.curr_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_1_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__20542\,
            in1 => \N__20554\,
            in2 => \N__20362\,
            in3 => \N__20359\,
            lcout => \b2v_inst16.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34643\,
            ce => \N__33684\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.delayed_vddq_pwrgd_RNIJ10L1_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011111111"
        )
    port map (
            in0 => \N__33715\,
            in1 => \N__20296\,
            in2 => \N__20548\,
            in3 => \N__25078\,
            lcout => b2v_inst16_un2_vpp_en_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_0_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__20541\,
            in1 => \_gnd_net_\,
            in2 => \N__25085\,
            in3 => \N__20627\,
            lcout => \b2v_inst16.curr_state_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34643\,
            ce => \N__33684\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNO_0_1_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__34059\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20560\,
            lcout => \b2v_inst16.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIKEBL_1_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20544\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33714\,
            lcout => \b2v_inst16.count_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_0_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__28990\,
            in1 => \N__25595\,
            in2 => \_gnd_net_\,
            in3 => \N__25389\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33081\,
            in2 => \_gnd_net_\,
            in3 => \N__20509\,
            lcout => \b2v_inst200.m11_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.DSW_PWROK_RNIUDI9_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34060\,
            in1 => \N__22156\,
            in2 => \_gnd_net_\,
            in3 => \N__29998\,
            lcout => \V105A_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__25390\,
            in1 => \N__26765\,
            in2 => \N__27436\,
            in3 => \N__28991\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_10_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20572\,
            in3 => \N__22355\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_5_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20596\,
            in1 => \N__21015\,
            in2 => \N__26782\,
            in3 => \N__28019\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_14_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__27307\,
            in1 => \N__20701\,
            in2 => \N__21186\,
            in3 => \N__20692\,
            lcout => \b2v_inst11.dutycycleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34621\,
            ce => 'H',
            sr => \N__24163\
        );

    \b2v_inst11.dutycycle_RNI2RTA8_14_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__20700\,
            in1 => \N__20691\,
            in2 => \N__21187\,
            in3 => \N__27306\,
            lcout => \b2v_inst11.dutycycleZ0Z_13\,
            ltout => \b2v_inst11.dutycycleZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_15_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21336\,
            in1 => \N__22309\,
            in2 => \N__20677\,
            in3 => \N__21153\,
            lcout => \b2v_inst11.un2_count_clk_17_0_a2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_10_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22786\,
            in2 => \_gnd_net_\,
            in3 => \N__22308\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_50_a4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_7_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101011"
        )
    port map (
            in0 => \N__26223\,
            in1 => \N__20668\,
            in2 => \N__20662\,
            in3 => \N__20658\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_1_sqmuxa_0_o2_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__28747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28307\,
            lcout => \b2v_inst11.N_158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst17.un4_vccio_en_0_a3_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__20641\,
            in1 => \N__20626\,
            in2 => \_gnd_net_\,
            in3 => \N__29652\,
            lcout => \VCCIO_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_10_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26212\,
            in2 => \_gnd_net_\,
            in3 => \N__22287\,
            lcout => \b2v_inst11.un1_dutycycle_53_axb_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011100000"
        )
    port map (
            in0 => \N__26211\,
            in1 => \N__22784\,
            in2 => \N__28962\,
            in3 => \N__24779\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_3\,
            ltout => \b2v_inst11.dutycycle_RNIZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_9_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110101000010"
        )
    port map (
            in0 => \N__28015\,
            in1 => \N__20976\,
            in2 => \N__20581\,
            in3 => \N__20578\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI03R98_4_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__27231\,
            in1 => \N__21064\,
            in2 => \N__20733\,
            in3 => \N__20742\,
            lcout => \b2v_inst11.dutycycleZ0Z_8\,
            ltout => \b2v_inst11.dutycycleZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIAI7C4_4_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001100"
        )
    port map (
            in0 => \N__22585\,
            in1 => \N__27234\,
            in2 => \N__20761\,
            in3 => \N__28118\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNIAI7C4Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI3JFN6_4_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101010"
        )
    port map (
            in0 => \N__27618\,
            in1 => \N__27751\,
            in2 => \N__20758\,
            in3 => \N__22242\,
            lcout => \b2v_inst11.dutycycle_RNI3JFN6Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI3JFN6_0_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001100000000"
        )
    port map (
            in0 => \N__22584\,
            in1 => \N__27750\,
            in2 => \N__20755\,
            in3 => \N__27617\,
            lcout => \b2v_inst11.func_state_RNI3JFN6Z0Z_0\,
            ltout => \b2v_inst11.func_state_RNI3JFN6Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_9_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__27233\,
            in1 => \N__20910\,
            in2 => \N__20746\,
            in3 => \N__20719\,
            lcout => \b2v_inst11.dutycycleZ1Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34635\,
            ce => 'H',
            sr => \N__24162\
        );

    \b2v_inst11.dutycycle_4_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__27232\,
            in1 => \N__21063\,
            in2 => \N__20734\,
            in3 => \N__20743\,
            lcout => \b2v_inst11.dutycycleZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34635\,
            ce => 'H',
            sr => \N__24162\
        );

    \b2v_inst11.dutycycle_RNIAI0A8_9_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__20718\,
            in1 => \N__20710\,
            in2 => \N__20914\,
            in3 => \N__27230\,
            lcout => \b2v_inst11.dutycycleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI0KJ31_7_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010101010101"
        )
    port map (
            in0 => \N__20799\,
            in1 => \N__21043\,
            in2 => \N__26881\,
            in3 => \N__26960\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI0KJ31Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI74A23_7_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__27275\,
            in1 => \_gnd_net_\,
            in2 => \N__20704\,
            in3 => \N__20785\,
            lcout => \b2v_inst11.dutycycle_RNI74A23Z0Z_7\,
            ltout => \b2v_inst11.dutycycle_RNI74A23Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIF271B_7_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000001111"
        )
    port map (
            in0 => \N__20797\,
            in1 => \N__20839\,
            in2 => \N__20842\,
            in3 => \N__27752\,
            lcout => \b2v_inst11.dutycycleZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI7UR36_0_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011111"
        )
    port map (
            in0 => \N__27274\,
            in1 => \N__28140\,
            in2 => \N__20809\,
            in3 => \N__22227\,
            lcout => \b2v_inst11.dutycycle_e_1_7\,
            ltout => \b2v_inst11.dutycycle_e_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_7_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101000110011"
        )
    port map (
            in0 => \N__20800\,
            in1 => \N__20833\,
            in2 => \N__20827\,
            in3 => \N__27753\,
            lcout => \b2v_inst11.dutycycleZ1Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34642\,
            ce => 'H',
            sr => \N__24210\
        );

    \b2v_inst11.dutycycle_RNI25OT3_7_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__24484\,
            in1 => \N__20824\,
            in2 => \_gnd_net_\,
            in3 => \N__26680\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI25OT3Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIGALV4_0_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__23290\,
            in1 => \N__26210\,
            in2 => \N__20812\,
            in3 => \N__23121\,
            lcout => \b2v_inst11.func_state_RNIGALV4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIGSFQ_7_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__26959\,
            in1 => \N__20798\,
            in2 => \_gnd_net_\,
            in3 => \N__26873\,
            lcout => \b2v_inst11.dutycycle_RNIGSFQZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_0_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25548\,
            in2 => \_gnd_net_\,
            in3 => \N__25383\,
            lcout => \b2v_inst11.g0_2_3\,
            ltout => OPEN,
            carryin => \bfn_6_13_0_\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_0_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29217\,
            in2 => \N__25392\,
            in3 => \N__20779\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_0_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDU8_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29237\,
            in2 => \N__27413\,
            in3 => \N__20764\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDUZ0Z8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_1\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29216\,
            in2 => \N__24816\,
            in3 => \N__21067\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_2\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29238\,
            in2 => \N__28992\,
            in3 => \N__21052\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_3\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_4_c_RNI578D1_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__27235\,
            in1 => \N__29222\,
            in2 => \N__26781\,
            in3 => \N__21049\,
            lcout => \b2v_inst11.g1_4_0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_4\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_5_c_RNI_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27956\,
            in2 => \N__29250\,
            in3 => \N__21046\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_5_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29221\,
            in2 => \N__26224\,
            in3 => \N__21037\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_6_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHP49_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22785\,
            in2 => \N__29247\,
            in3 => \N__21019\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHPZ0Z49\,
            ltout => OPEN,
            carryin => \bfn_6_14_0_\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIR59_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29214\,
            in2 => \N__21016\,
            in3 => \N__20899\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_8_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_9_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJT69_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22349\,
            in2 => \N__29248\,
            in3 => \N__20896\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJTZ0Z69\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_9_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNP5_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29200\,
            in2 => \N__20893\,
            in3 => \N__21445\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNPZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_10\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQ5_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21435\,
            in2 => \N__29246\,
            in3 => \N__21340\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_11\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29201\,
            in2 => \N__21337\,
            in3 => \N__21250\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_12\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21247\,
            in2 => \N__29249\,
            in3 => \N__21166\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_13\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__21163\,
            in1 => \N__29215\,
            in2 => \_gnd_net_\,
            in3 => \N__21109\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_5_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__25346\,
            in1 => \N__26780\,
            in2 => \N__25570\,
            in3 => \N__27912\,
            lcout => \b2v_inst11.dutycycle_RNI_5Z0Z_5\,
            ltout => \b2v_inst11.dutycycle_RNI_5Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_0_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__23110\,
            in1 => \N__24279\,
            in2 => \N__21085\,
            in3 => \N__23204\,
            lcout => \b2v_inst11.N_156\,
            ltout => \b2v_inst11.N_156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_2_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21076\,
            in3 => \N__23174\,
            lcout => \b2v_inst11.N_418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINJ641_1_1_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__24722\,
            in1 => \N__23238\,
            in2 => \_gnd_net_\,
            in3 => \N__24278\,
            lcout => \b2v_inst11.N_331\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23205\,
            in1 => \N__29235\,
            in2 => \N__23056\,
            in3 => \N__23175\,
            lcout => \b2v_inst11.un1_func_state25_6_0_o_N_307_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_1_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28454\,
            in2 => \_gnd_net_\,
            in3 => \N__24277\,
            lcout => \b2v_inst11.N_169\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIQQRO_5_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21493\,
            in1 => \N__24854\,
            in2 => \N__23184\,
            in3 => \N__25065\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI8PGM6_5_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101011101"
        )
    port map (
            in0 => \N__27776\,
            in1 => \N__29023\,
            in2 => \N__21481\,
            in3 => \N__23455\,
            lcout => \b2v_inst11.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_0_0_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23109\,
            in2 => \N__23206\,
            in3 => \N__23183\,
            lcout => \b2v_inst11.func_state_RNI_0Z0Z_0\,
            ltout => \b2v_inst11.func_state_RNI_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINJ641_0_0_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21478\,
            in3 => \N__24723\,
            lcout => \b2v_inst11.func_state_RNINJ641_0Z0Z_0\,
            ltout => \b2v_inst11.func_state_RNINJ641_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIQCBN4_9_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__21463\,
            in1 => \N__27772\,
            in2 => \N__21469\,
            in3 => \N__23308\,
            lcout => \b2v_inst11.count_off_RNIQCBN4Z0Z_9\,
            ltout => \b2v_inst11.count_off_RNIQCBN4Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDINH9_0_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__21547\,
            in1 => \N__21526\,
            in2 => \N__21466\,
            in3 => \N__25066\,
            lcout => \b2v_inst11.func_state_RNIDINH9Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI7J1P_1_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__28674\,
            in1 => \N__34006\,
            in2 => \N__28308\,
            in3 => \N__21598\,
            lcout => \b2v_inst11.N_333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIQBAL3_1_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111101111"
        )
    port map (
            in0 => \N__21599\,
            in1 => \N__21553\,
            in2 => \N__27781\,
            in3 => \N__24096\,
            lcout => \b2v_inst11.N_73\,
            ltout => \b2v_inst11.N_73_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI673P9_0_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001010100"
        )
    port map (
            in0 => \N__25067\,
            in1 => \N__21541\,
            in2 => \N__21535\,
            in3 => \N__21532\,
            lcout => \b2v_inst11.func_state_RNI673P9Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIPAG14_0_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__23467\,
            in1 => \N__23212\,
            in2 => \N__23427\,
            in3 => \N__24724\,
            lcout => \b2v_inst11.func_state_1_m0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23953\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_2_0_\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21713\,
            in2 => \N__21757\,
            in3 => \N__21520\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21703\,
            in2 => \N__21718\,
            in3 => \N__21517\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21855\,
            in2 => \N__21685\,
            in3 => \N__21514\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21661\,
            in2 => \N__21859\,
            in3 => \N__21511\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__23709\,
            in1 => \N__21717\,
            in2 => \N__21646\,
            in3 => \N__21508\,
            lcout => \b2v_inst11.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21610\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21721\,
            lcout => \b2v_inst11.mult1_un145_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21854\,
            lcout => \b2v_inst11.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21778\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_3_0_\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21994\,
            in2 => \N__21627\,
            in3 => \N__21697\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21623\,
            in2 => \N__21694\,
            in3 => \N__21676\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21797\,
            in2 => \N__21673\,
            in3 => \N__21655\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21652\,
            in2 => \N__21802\,
            in3 => \N__21637\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__21853\,
            in1 => \N__21634\,
            in2 => \N__21628\,
            in3 => \N__21604\,
            lcout => \b2v_inst11.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__21868\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21862\,
            lcout => \b2v_inst11.mult1_un138_sum_s_8\,
            ltout => \b2v_inst11.mult1_un138_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21838\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un85_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23718\,
            lcout => \b2v_inst11.un85_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23619\,
            lcout => \b2v_inst11.un85_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23949\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25465\,
            lcout => \b2v_inst11.un85_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21835\,
            lcout => \b2v_inst11.un85_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21801\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un85_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21774\,
            lcout => \b2v_inst11.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21745\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26536\,
            in1 => \N__25408\,
            in2 => \N__21988\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un1_count_cry_0_i\,
            ltout => OPEN,
            carryin => \bfn_7_5_0_\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21964\,
            in2 => \N__21973\,
            in3 => \N__26563\,
            lcout => \b2v_inst11.N_5647_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_0\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25920\,
            in1 => \N__21958\,
            in2 => \N__21952\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5648_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_1\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25624\,
            in1 => \N__21943\,
            in2 => \N__21937\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5649_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_2\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21913\,
            in2 => \N__21925\,
            in3 => \N__26029\,
            lcout => \b2v_inst11.N_5650_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_3\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21898\,
            in2 => \N__21907\,
            in3 => \N__25987\,
            lcout => \b2v_inst11.N_5651_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_4\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25758\,
            in1 => \N__21892\,
            in2 => \N__21886\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5652_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_5\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22120\,
            in2 => \N__21877\,
            in3 => \N__25894\,
            lcout => \b2v_inst11.N_5653_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_6\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26407\,
            in1 => \N__22105\,
            in2 => \N__22114\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5654_i\,
            ltout => OPEN,
            carryin => \bfn_7_6_0_\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26364\,
            in1 => \N__22099\,
            in2 => \N__22087\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5655_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_8\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22069\,
            in2 => \N__22078\,
            in3 => \N__25819\,
            lcout => \b2v_inst11.N_5656_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_9\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25846\,
            in1 => \N__22063\,
            in2 => \N__22051\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5657_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_10\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22030\,
            in2 => \N__22042\,
            in3 => \N__25787\,
            lcout => \b2v_inst11.N_5658_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_11\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26071\,
            in1 => \N__22024\,
            in2 => \N__22018\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5659_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_12\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22000\,
            in2 => \N__22009\,
            in3 => \N__25731\,
            lcout => \b2v_inst11.N_5660_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_13\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22165\,
            in2 => \N__22174\,
            in3 => \N__25866\,
            lcout => \b2v_inst11.N_5661_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_14\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_15_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22159\,
            lcout => \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_0_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26531\,
            in2 => \_gnd_net_\,
            in3 => \N__26440\,
            lcout => \b2v_inst11.count_RNI_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__25701\,
            in1 => \N__25656\,
            in2 => \_gnd_net_\,
            in3 => \N__26638\,
            lcout => \b2v_inst11.curr_state_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNI8TT2_0_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__30402\,
            in1 => \N__30306\,
            in2 => \_gnd_net_\,
            in3 => \N__30358\,
            lcout => \b2v_inst36.curr_state_RNI8TT2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_15_c_RNICRLO_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__25655\,
            in1 => \N__22126\,
            in2 => \N__26649\,
            in3 => \N__33718\,
            lcout => OPEN,
            ltout => \b2v_inst11.pwm_out_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.pwm_out_RNIEV5S_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26611\,
            in2 => \N__22147\,
            in3 => \N__25654\,
            lcout => \PWRBTN_LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNIOCA3_0_0_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__25653\,
            in1 => \_gnd_net_\,
            in2 => \N__34085\,
            in3 => \N__25700\,
            lcout => \b2v_inst11.pwm_out_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_0_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26642\,
            in2 => \N__25702\,
            in3 => \N__25652\,
            lcout => \b2v_inst11.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34637\,
            ce => \N__33679\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNIJK34_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22432\,
            in1 => \N__34036\,
            in2 => \_gnd_net_\,
            in3 => \N__22426\,
            lcout => \b2v_inst11.curr_stateZ0Z_0\,
            ltout => \b2v_inst11.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNIOCA3_0_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__34037\,
            in1 => \_gnd_net_\,
            in2 => \N__22420\,
            in3 => \N__25696\,
            lcout => \b2v_inst11.count_0_sqmuxa_i\,
            ltout => \b2v_inst11.count_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_0_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22417\,
            in3 => \N__26535\,
            lcout => \b2v_inst11.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34637\,
            ce => \N__33679\,
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_4_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__31005\,
            in1 => \N__30985\,
            in2 => \_gnd_net_\,
            in3 => \N__26878\,
            lcout => \b2v_inst20.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34625\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_3_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26236\,
            in1 => \N__24818\,
            in2 => \N__25596\,
            in3 => \N__25391\,
            lcout => \b2v_inst11.g0_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIJU083_0_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010111111"
        )
    port map (
            in0 => \N__23251\,
            in1 => \N__24464\,
            in2 => \N__27090\,
            in3 => \N__27021\,
            lcout => \b2v_inst11.func_state_RNIJU083Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_3_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__24817\,
            in1 => \N__28994\,
            in2 => \_gnd_net_\,
            in3 => \N__26235\,
            lcout => \b2v_inst11.N_349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIAI7C4_10_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__22244\,
            in1 => \N__22310\,
            in2 => \N__22577\,
            in3 => \N__22401\,
            lcout => \b2v_inst11.dutycycle_RNIAI7C4Z0Z_10\,
            ltout => \b2v_inst11.dutycycle_RNIAI7C4Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIP8IN8_10_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100110001"
        )
    port map (
            in0 => \N__27693\,
            in1 => \N__22513\,
            in2 => \N__22366\,
            in3 => \N__22493\,
            lcout => \b2v_inst11.dutycycleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNINJ641_3_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001110"
        )
    port map (
            in0 => \N__27257\,
            in1 => \N__28153\,
            in2 => \N__24812\,
            in3 => \N__22243\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_clk_100khz_43_and_i_o2_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI3JFN6_3_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000000"
        )
    port map (
            in0 => \N__22553\,
            in1 => \N__27692\,
            in2 => \N__22528\,
            in3 => \N__27535\,
            lcout => \b2v_inst11.dutycycle_e_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.N_221_i_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__29071\,
            in1 => \N__29314\,
            in2 => \N__34091\,
            in3 => \N__28591\,
            lcout => \b2v_inst11.N_221_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI4I3C2_10_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001111"
        )
    port map (
            in0 => \N__22525\,
            in1 => \N__27258\,
            in2 => \N__22498\,
            in3 => \N__27536\,
            lcout => \b2v_inst11.dutycycle_RNI4I3C2Z0Z_10\,
            ltout => \b2v_inst11.dutycycle_RNI4I3C2Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_10_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111110001101"
        )
    port map (
            in0 => \N__27694\,
            in1 => \N__22497\,
            in2 => \N__22507\,
            in3 => \N__22504\,
            lcout => \b2v_inst11.dutycycleZ1Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34636\,
            ce => 'H',
            sr => \N__24160\
        );

    \b2v_inst11.dutycycle_RNI_1_5_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22763\,
            in1 => \N__22831\,
            in2 => \N__26757\,
            in3 => \N__28956\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_3_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__27229\,
            in1 => \N__22800\,
            in2 => \N__22813\,
            in3 => \N__22825\,
            lcout => \b2v_inst11.dutycycleZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34644\,
            ce => 'H',
            sr => \N__24161\
        );

    \b2v_inst11.dutycycle_RNI_4_3_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25379\,
            in2 => \N__24807\,
            in3 => \N__27987\,
            lcout => OPEN,
            ltout => \b2v_inst11.d_i3_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_5_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__23977\,
            in1 => \N__22446\,
            in2 => \N__22468\,
            in3 => \N__26732\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_3_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__26180\,
            in1 => \_gnd_net_\,
            in2 => \N__24808\,
            in3 => \N__28955\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_3_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__28954\,
            in1 => \N__24782\,
            in2 => \_gnd_net_\,
            in3 => \N__26179\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIUVP98_3_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__22824\,
            in1 => \N__22809\,
            in2 => \N__22801\,
            in3 => \N__27228\,
            lcout => \b2v_inst11.dutycycleZ0Z_6\,
            ltout => \b2v_inst11.dutycycleZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_3_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010111"
        )
    port map (
            in0 => \N__28953\,
            in1 => \N__26178\,
            in2 => \N__22789\,
            in3 => \N__22762\,
            lcout => \b2v_inst11.dutycycle_RNI_5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINJ641_0_1_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011101"
        )
    port map (
            in0 => \N__27029\,
            in1 => \N__24482\,
            in2 => \N__27109\,
            in3 => \N__22912\,
            lcout => \b2v_inst11.func_state_RNINJ641_0Z0Z_1\,
            ltout => \b2v_inst11.func_state_RNINJ641_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNINJ641_2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__27389\,
            in1 => \N__24393\,
            in2 => \N__22636\,
            in3 => \N__24315\,
            lcout => \b2v_inst11.g0_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_0_o3_1_1_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28739\,
            in2 => \_gnd_net_\,
            in3 => \N__28322\,
            lcout => \b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1\,
            ltout => \b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111101111111"
        )
    port map (
            in0 => \N__24483\,
            in1 => \N__27103\,
            in2 => \N__22633\,
            in3 => \N__27030\,
            lcout => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_6_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22630\,
            in1 => \N__22624\,
            in2 => \N__28013\,
            in3 => \N__28168\,
            lcout => \b2v_inst11.un1_dutycycle_164_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_4_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__28930\,
            in1 => \N__26187\,
            in2 => \_gnd_net_\,
            in3 => \N__27965\,
            lcout => \b2v_inst11.g0_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010111111111"
        )
    port map (
            in0 => \N__28746\,
            in1 => \N__33994\,
            in2 => \N__28345\,
            in3 => \N__29085\,
            lcout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIF6NL_1_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__28740\,
            in1 => \_gnd_net_\,
            in2 => \N__28343\,
            in3 => \N__28395\,
            lcout => \b2v_inst11.un1_clk_100khz_2_i_o3_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__27547\,
            in1 => \N__22900\,
            in2 => \N__24544\,
            in3 => \N__22894\,
            lcout => \b2v_inst11.dutycycleZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34653\,
            ce => 'H',
            sr => \N__24187\
        );

    \b2v_inst11.un1_dutycycle_94_cry_0_c_RNI1V3D1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110011"
        )
    port map (
            in0 => \N__23113\,
            in1 => \N__22906\,
            in2 => \N__23053\,
            in3 => \N__28405\,
            lcout => \b2v_inst11.dutycycle_1_0_1\,
            ltout => \b2v_inst11.dutycycle_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIP4GA6_1_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__27546\,
            in1 => \N__22893\,
            in2 => \N__22885\,
            in3 => \N__24537\,
            lcout => \b2v_inst11.dutycycle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_1_0_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__23112\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28404\,
            lcout => \b2v_inst11.func_state_RNI_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_0_1_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28403\,
            in2 => \_gnd_net_\,
            in3 => \N__23422\,
            lcout => \b2v_inst11.func_state_RNI_0Z0Z_1\,
            ltout => \b2v_inst11.func_state_RNI_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_3_0_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001111"
        )
    port map (
            in0 => \N__23423\,
            in1 => \N__28429\,
            in2 => \N__22852\,
            in3 => \N__23111\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_func_state25_4_i_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIOJI01_0_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__28577\,
            in1 => \_gnd_net_\,
            in2 => \N__22849\,
            in3 => \N__29660\,
            lcout => \b2v_inst11.N_321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_6_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__22984\,
            in1 => \N__22990\,
            in2 => \N__27620\,
            in3 => \N__22972\,
            lcout => \b2v_inst11.dutycycle_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34659\,
            ce => 'H',
            sr => \N__24214\
        );

    \b2v_inst11.func_state_RNINJ641_0_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__25549\,
            in1 => \N__28413\,
            in2 => \N__23055\,
            in3 => \N__23114\,
            lcout => \b2v_inst11.dutycycle_1_0_0\,
            ltout => \b2v_inst11.dutycycle_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIEOI16_0_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100001000"
        )
    port map (
            in0 => \N__27606\,
            in1 => \N__22960\,
            in2 => \N__23005\,
            in3 => \N__22941\,
            lcout => \b2v_inst11.dutycycleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIKOJB2_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__24109\,
            in1 => \N__27262\,
            in2 => \N__26965\,
            in3 => \N__23002\,
            lcout => \b2v_inst11.g1\,
            ltout => \b2v_inst11.g1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIBDKS9_6_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__27603\,
            in1 => \N__22983\,
            in2 => \N__22975\,
            in3 => \N__22971\,
            lcout => \b2v_inst11.dutycycleZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIEFS24_0_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111101"
        )
    port map (
            in0 => \N__27770\,
            in1 => \N__25550\,
            in2 => \N__29678\,
            in3 => \N__24835\,
            lcout => \b2v_inst11.dutycycle_eena\,
            ltout => \b2v_inst11.dutycycle_eena_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_0_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__22942\,
            in1 => \N__22951\,
            in2 => \N__22945\,
            in3 => \N__27610\,
            lcout => \b2v_inst11.dutycycleZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34659\,
            ce => 'H',
            sr => \N__24214\
        );

    \b2v_inst11.count_clk_RNI_2_3_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__29277\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28158\,
            lcout => \N_19_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_9_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23383\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_RNIZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNITBKN1_1_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001111"
        )
    port map (
            in0 => \N__28678\,
            in1 => \N__24493\,
            in2 => \N__28290\,
            in3 => \N__28157\,
            lcout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1\,
            ltout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIBHHP2_0_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__23284\,
            in1 => \_gnd_net_\,
            in2 => \N__23254\,
            in3 => \N__23108\,
            lcout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI2N9T2_1_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__27771\,
            in1 => \N__23231\,
            in2 => \_gnd_net_\,
            in3 => \N__23062\,
            lcout => \b2v_inst11.func_state_1_m0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_0_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27957\,
            in1 => \N__25551\,
            in2 => \N__24378\,
            in3 => \N__25318\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_0\,
            ltout => \b2v_inst11.dutycycle_RNI_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIF6NL_2_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101111111"
        )
    port map (
            in0 => \N__23188\,
            in1 => \N__23143\,
            in2 => \N__23134\,
            in3 => \N__28159\,
            lcout => \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIS50RB_0_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__27604\,
            in1 => \N__24690\,
            in2 => \N__23440\,
            in3 => \N__23448\,
            lcout => \b2v_inst11.func_stateZ0Z_0\,
            ltout => \b2v_inst11.func_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_2_0_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23068\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_3013_i\,
            ltout => \b2v_inst11.N_3013_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIT4D71_9_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__23414\,
            in1 => \N__28576\,
            in2 => \N__23065\,
            in3 => \N__24082\,
            lcout => \b2v_inst11.N_330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI70K8_0_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28276\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23466\,
            lcout => \b2v_inst11.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_0_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__23449\,
            in1 => \N__23439\,
            in2 => \N__24694\,
            in3 => \N__27605\,
            lcout => \b2v_inst11.func_stateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34669\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_0_9_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23415\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29284\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_335_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNINJ641_9_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__24291\,
            in1 => \N__24716\,
            in2 => \N__23386\,
            in3 => \N__23378\,
            lcout => \b2v_inst11.func_state_1_ss0_i_0_o2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI_2_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29968\,
            in1 => \N__24918\,
            in2 => \N__25179\,
            in3 => \N__29909\,
            lcout => \b2v_inst36.un12_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_2_c_RNIBSB8_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__29883\,
            in1 => \N__32205\,
            in2 => \N__29914\,
            in3 => \N__32080\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIH5D01_3_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__31932\,
            in1 => \N__29872\,
            in2 => \N__23302\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIPHH01_7_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23296\,
            in1 => \N__31934\,
            in2 => \_gnd_net_\,
            in3 => \N__23488\,
            lcout => \b2v_inst36.countZ0Z_7\,
            ltout => \b2v_inst36.countZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_7_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__32082\,
            in1 => \N__32208\,
            in2 => \N__23299\,
            in3 => \N__25156\,
            lcout => \b2v_inst36.count_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34682\,
            ce => \N__31935\,
            sr => \N__31827\
        );

    \b2v_inst36.un2_count_1_cry_4_c_RNID0E8_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__24903\,
            in1 => \N__32206\,
            in2 => \N__24922\,
            in3 => \N__32081\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNILBF01_5_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31933\,
            in1 => \_gnd_net_\,
            in2 => \N__23500\,
            in3 => \N__23494\,
            lcout => \b2v_inst36.countZ0Z_5\,
            ltout => \b2v_inst36.countZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_5_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__24904\,
            in1 => \N__32207\,
            in2 => \N__23497\,
            in3 => \N__32083\,
            lcout => \b2v_inst36.count_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34682\,
            ce => \N__31935\,
            sr => \N__31827\
        );

    \b2v_inst36.un2_count_1_cry_10_c_RNIQ3J1_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__32086\,
            in1 => \N__30084\,
            in2 => \N__29749\,
            in3 => \N__32197\,
            lcout => \b2v_inst36.count_rst_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_6_c_RNIF4G8_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__25180\,
            in1 => \N__32193\,
            in2 => \N__32089\,
            in3 => \N__25152\,
            lcout => \b2v_inst36.count_rst_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_7_c_RNIG6H8_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__32084\,
            in1 => \N__29859\,
            in2 => \N__25138\,
            in3 => \N__32196\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIRKI01_8_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23476\,
            in2 => \N__23482\,
            in3 => \N__31907\,
            lcout => \b2v_inst36.countZ0Z_8\,
            ltout => \b2v_inst36.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_8_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__32087\,
            in1 => \N__25137\,
            in2 => \N__23479\,
            in3 => \N__32198\,
            lcout => \b2v_inst36.count_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34675\,
            ce => \N__31976\,
            sr => \N__31840\
        );

    \b2v_inst36.un2_count_1_cry_9_c_RNIIAJ8_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__25116\,
            in1 => \N__32194\,
            in2 => \N__29841\,
            in3 => \N__32085\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI6MB61_10_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31908\,
            in1 => \_gnd_net_\,
            in2 => \N__23470\,
            in3 => \N__23575\,
            lcout => \b2v_inst36.countZ0Z_10\,
            ltout => \b2v_inst36.countZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_10_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__25117\,
            in1 => \N__32195\,
            in2 => \N__23578\,
            in3 => \N__32088\,
            lcout => \b2v_inst36.count_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34675\,
            ce => \N__31976\,
            sr => \N__31840\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27426\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23684\,
            in2 => \N__23569\,
            in3 => \N__23557\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23554\,
            in2 => \N__23689\,
            in3 => \N__23548\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23714\,
            in2 => \N__23545\,
            in3 => \N__23536\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23533\,
            in2 => \N__23719\,
            in3 => \N__23527\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__23613\,
            in1 => \N__23688\,
            in2 => \N__23524\,
            in3 => \N__23512\,
            lcout => \b2v_inst11.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__23509\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23503\,
            lcout => \b2v_inst11.mult1_un152_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23713\,
            lcout => \b2v_inst11.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25384\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23588\,
            in2 => \N__24343\,
            in3 => \N__23674\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_1\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23671\,
            in2 => \N__23593\,
            in3 => \N__23665\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23615\,
            in2 => \N__23662\,
            in3 => \N__23653\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23650\,
            in2 => \N__23620\,
            in3 => \N__23644\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__25464\,
            in1 => \N__23592\,
            in2 => \N__23641\,
            in3 => \N__23632\,
            lcout => \b2v_inst11.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__23629\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23623\,
            lcout => \b2v_inst11.mult1_un159_sum_s_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23614\,
            lcout => \b2v_inst11.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIQF4M_14_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23743\,
            in1 => \N__34055\,
            in2 => \_gnd_net_\,
            in3 => \N__23847\,
            lcout => \b2v_inst11.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_14_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23851\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34661\,
            ce => \N__33687\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIS3FN_6_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23737\,
            in1 => \N__34053\,
            in2 => \_gnd_net_\,
            in3 => \N__23775\,
            lcout => \b2v_inst11.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_6_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23776\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34661\,
            ce => \N__33687\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNISI5M_15_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23731\,
            in1 => \N__34056\,
            in2 => \_gnd_net_\,
            in3 => \N__23826\,
            lcout => \b2v_inst11.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_15_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23830\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34661\,
            ce => \N__33687\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIU6GN_7_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23725\,
            in1 => \N__34054\,
            in2 => \_gnd_net_\,
            in3 => \N__23763\,
            lcout => \b2v_inst11.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_7_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23764\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34661\,
            ce => \N__33687\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_1_c_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26517\,
            in2 => \N__26559\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \b2v_inst11.un1_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__26479\,
            in1 => \_gnd_net_\,
            in2 => \N__25921\,
            in3 => \N__23788\,
            lcout => \b2v_inst11.un1_count_cry_1_c_RNIIIQDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_1\,
            carryout => \b2v_inst11.un1_count_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__26483\,
            in1 => \_gnd_net_\,
            in2 => \N__25620\,
            in3 => \N__23785\,
            lcout => \b2v_inst11.un1_count_cry_2_c_RNIJKRDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_2\,
            carryout => \b2v_inst11.un1_count_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__26480\,
            in1 => \_gnd_net_\,
            in2 => \N__26025\,
            in3 => \N__23782\,
            lcout => \b2v_inst11.un1_count_cry_3_c_RNIKMSDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_3\,
            carryout => \b2v_inst11.un1_count_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__26484\,
            in1 => \_gnd_net_\,
            in2 => \N__25983\,
            in3 => \N__23779\,
            lcout => \b2v_inst11.un1_count_cry_4_c_RNILOTDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_4\,
            carryout => \b2v_inst11.un1_count_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__26481\,
            in1 => \_gnd_net_\,
            in2 => \N__25759\,
            in3 => \N__23767\,
            lcout => \b2v_inst11.un1_count_cry_5_c_RNIMQUDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_5\,
            carryout => \b2v_inst11.un1_count_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__26485\,
            in1 => \_gnd_net_\,
            in2 => \N__25893\,
            in3 => \N__23755\,
            lcout => \b2v_inst11.un1_count_cry_6_c_RNINSVDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_6\,
            carryout => \b2v_inst11.un1_count_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26482\,
            in1 => \N__26396\,
            in2 => \_gnd_net_\,
            in3 => \N__23752\,
            lcout => \b2v_inst11.un1_count_cry_7_c_RNIOU0EZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_7\,
            carryout => \b2v_inst11.un1_count_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__26488\,
            in1 => \_gnd_net_\,
            in2 => \N__26354\,
            in3 => \N__23749\,
            lcout => \b2v_inst11.un1_count_cry_8_c_RNIP02EZ0\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \b2v_inst11.un1_count_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__26462\,
            in1 => \_gnd_net_\,
            in2 => \N__25814\,
            in3 => \N__23746\,
            lcout => \b2v_inst11.un1_count_cry_9_c_RNIQ23EZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_9\,
            carryout => \b2v_inst11.un1_count_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26489\,
            in1 => \N__25835\,
            in2 => \_gnd_net_\,
            in3 => \N__23860\,
            lcout => \b2v_inst11.un1_count_cry_10_c_RNI24RZ0Z6\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_10\,
            carryout => \b2v_inst11.un1_count_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__26463\,
            in1 => \_gnd_net_\,
            in2 => \N__25788\,
            in3 => \N__23857\,
            lcout => \b2v_inst11.un1_count_cry_11_c_RNI36SZ0Z6\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_11\,
            carryout => \b2v_inst11.un1_count_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__26490\,
            in1 => \_gnd_net_\,
            in2 => \N__26070\,
            in3 => \N__23854\,
            lcout => \b2v_inst11.un1_count_cry_12_c_RNI48TZ0Z6\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_12\,
            carryout => \b2v_inst11.un1_count_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__26464\,
            in1 => \_gnd_net_\,
            in2 => \N__25735\,
            in3 => \N__23836\,
            lcout => \b2v_inst11.un1_count_cry_13_c_RNI5AUZ0Z6\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_13\,
            carryout => \b2v_inst11.un1_count_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__26491\,
            in1 => \N__25870\,
            in2 => \_gnd_net_\,
            in3 => \N__23833\,
            lcout => \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIM92M_12_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23893\,
            in1 => \N__34057\,
            in2 => \_gnd_net_\,
            in3 => \N__23904\,
            lcout => \b2v_inst11.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIB49T_10_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23803\,
            in2 => \N__23815\,
            in3 => \N__34051\,
            lcout => \b2v_inst11.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_10_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23814\,
            lcout => \b2v_inst11.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34646\,
            ce => \N__33682\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIK61M_11_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23929\,
            in1 => \N__34052\,
            in2 => \_gnd_net_\,
            in3 => \N__23796\,
            lcout => \b2v_inst11.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_11_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23797\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34646\,
            ce => \N__33682\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIKNAN_2_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23911\,
            in1 => \N__34050\,
            in2 => \_gnd_net_\,
            in3 => \N__23922\,
            lcout => \b2v_inst11.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_2_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23923\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34646\,
            ce => \N__33682\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_12_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23905\,
            lcout => \b2v_inst11.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34646\,
            ce => \N__33682\,
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_7_1_0__m6_i_a2_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23874\,
            in2 => \_gnd_net_\,
            in3 => \N__32959\,
            lcout => \G_2727\,
            ltout => \G_2727_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_1_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23887\,
            in3 => \N__26668\,
            lcout => \b2v_inst5.curr_state_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34629\,
            ce => \N__33680\,
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__34753\,
            in1 => \N__26306\,
            in2 => \_gnd_net_\,
            in3 => \N__23875\,
            lcout => \RSMRSTn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34629\,
            ce => \N__33680\,
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNITB7B1_1_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__23873\,
            in1 => \N__34065\,
            in2 => \N__26308\,
            in3 => \N__34756\,
            lcout => \b2v_inst5.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_7_1_0__m6_i_o3_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__34754\,
            in1 => \N__26301\,
            in2 => \_gnd_net_\,
            in3 => \N__23872\,
            lcout => \N_229\,
            ltout => \N_229_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNI76HI_1_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__26282\,
            in1 => \N__23884\,
            in2 => \N__23878\,
            in3 => \N__34064\,
            lcout => \b2v_inst5.curr_stateZ0Z_1\,
            ltout => \b2v_inst5.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNI5VS71_1_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__34755\,
            in1 => \_gnd_net_\,
            in2 => \N__23959\,
            in3 => \N__26305\,
            lcout => \curr_state_RNI5VS71_0_1\,
            ltout => \curr_state_RNI5VS71_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_0_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011110010"
        )
    port map (
            in0 => \N__26283\,
            in1 => \N__26307\,
            in2 => \N__23956\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.curr_state_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34629\,
            ce => \N__33680\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_3_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25589\,
            in2 => \_gnd_net_\,
            in3 => \N__24795\,
            lcout => \b2v_inst11.mult1_un145_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_fast_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24455\,
            in2 => \_gnd_net_\,
            in3 => \N__26866\,
            lcout => \SYNTHESIZED_WIRE_47keep_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34645\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_0_c_RNO_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31079\,
            in1 => \N__31001\,
            in2 => \N__31044\,
            in3 => \N__31108\,
            lcout => \b2v_inst20.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.G_146_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26925\,
            in2 => \_gnd_net_\,
            in3 => \N__26827\,
            lcout => b2v_inst16_delayed_vddq_pwrgd_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_RNI8DFE_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27071\,
            in2 => \N__24468\,
            in3 => \N__27004\,
            lcout => \RSMRSTn_RNI8DFE\,
            ltout => \RSMRSTn_RNI8DFE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_0_sqmuxa_0_o2_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__29328\,
            in1 => \N__28597\,
            in2 => \N__23932\,
            in3 => \N__26924\,
            lcout => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_0_sqmuxa_0_o2_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__26926\,
            in1 => \N__27070\,
            in2 => \N__28753\,
            in3 => \N__28347\,
            lcout => \b2v_inst11.N_182\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIE5T11_2_1_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__28573\,
            in1 => \N__27091\,
            in2 => \N__29353\,
            in3 => \N__29273\,
            lcout => \b2v_inst11.g0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_5_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011111100"
        )
    port map (
            in0 => \N__24028\,
            in1 => \N__24018\,
            in2 => \N__24037\,
            in3 => \N__27451\,
            lcout => \b2v_inst11.dutycycle_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34649\,
            ce => 'H',
            sr => \N__24164\
        );

    \b2v_inst11.func_state_RNIT4D71_0_1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__24058\,
            in1 => \N__28574\,
            in2 => \_gnd_net_\,
            in3 => \N__29272\,
            lcout => \b2v_inst11.func_state_RNIT4D71_0Z0Z_1\,
            ltout => \b2v_inst11.func_state_RNIT4D71_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIIOE3D_5_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111100"
        )
    port map (
            in0 => \N__24027\,
            in1 => \N__24019\,
            in2 => \N__24004\,
            in3 => \N__27450\,
            lcout => \dutycycle_RNIIOE3D_0_5\,
            ltout => \dutycycle_RNIIOE3D_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_5_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24001\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_5\,
            ltout => \b2v_inst11.dutycycle_RNI_4Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110101"
        )
    port map (
            in0 => \N__25333\,
            in1 => \_gnd_net_\,
            in2 => \N__23998\,
            in3 => \N__28958\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_axb_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_2_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100101101001"
        )
    port map (
            in0 => \N__27986\,
            in1 => \N__24781\,
            in2 => \N__23995\,
            in3 => \N__27409\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_3_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__24780\,
            in1 => \N__27985\,
            in2 => \N__25360\,
            in3 => \N__28957\,
            lcout => \b2v_inst11.un1_i3_mux_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_4_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__28163\,
            in1 => \N__23971\,
            in2 => \_gnd_net_\,
            in3 => \N__28993\,
            lcout => \b2v_inst11.un1_dutycycle_inv_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__24526\,
            in1 => \N__24421\,
            in2 => \N__28020\,
            in3 => \N__28164\,
            lcout => \b2v_inst11.N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNINJ641_5_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__28744\,
            in1 => \N__29092\,
            in2 => \N__28344\,
            in3 => \N__24364\,
            lcout => OPEN,
            ltout => \b2v_inst11.g1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIE7D82_2_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001110010"
        )
    port map (
            in0 => \N__24412\,
            in1 => \N__24406\,
            in2 => \N__24397\,
            in3 => \N__24394\,
            lcout => \b2v_inst11.un1_dutycycle_172_m4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.SYNTHESIZED_WIRE_49_i_0_o3_0_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101111111"
        )
    port map (
            in0 => \N__27092\,
            in1 => \N__26927\,
            in2 => \N__28752\,
            in3 => \N__27028\,
            lcout => \SYNTHESIZED_WIRE_49_i_0_o3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_5_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__24365\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28828\,
            lcout => \G_26_0_a5_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27408\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINJ641_1_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__24324\,
            in1 => \N__27236\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => b2v_inst11_count_off_1_sqmuxa_0_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_2_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0111111100001000"
        )
    port map (
            in0 => \N__27550\,
            in1 => \N__24586\,
            in2 => \N__24580\,
            in3 => \N__24553\,
            lcout => \b2v_inst11.dutycycleZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34660\,
            ce => 'H',
            sr => \N__24236\
        );

    \b2v_inst11.func_state_RNI4IKJB_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__24676\,
            in1 => \N__27548\,
            in2 => \N__24628\,
            in3 => \N__24651\,
            lcout => \b2v_inst11.func_state\,
            ltout => \b2v_inst11.func_state_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIPKCK_2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010001"
        )
    port map (
            in0 => \N__29634\,
            in1 => \N__29286\,
            in2 => \N__24592\,
            in3 => \N__27382\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_303_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNILQFE3_2_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100110011"
        )
    port map (
            in0 => \N__24677\,
            in1 => \N__27754\,
            in2 => \N__24589\,
            in3 => \N__24874\,
            lcout => \b2v_inst11.dutycycle_eena_1\,
            ltout => \b2v_inst11.dutycycle_eena_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI6O567_2_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__27549\,
            in1 => \N__24579\,
            in2 => \N__24556\,
            in3 => \N__24552\,
            lcout => \b2v_inst11.dutycycleZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIEFS24_1_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111101111"
        )
    port map (
            in0 => \N__25308\,
            in1 => \N__29633\,
            in2 => \N__27741\,
            in3 => \N__24831\,
            lcout => \b2v_inst11.dutycycle_eena_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIOJI01_1_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100110101"
        )
    port map (
            in0 => \N__28582\,
            in1 => \N__28798\,
            in2 => \N__29671\,
            in3 => \N__24525\,
            lcout => \b2v_inst11.un1_clk_100khz_26_and_i_o2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIE5T11_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100000000"
        )
    port map (
            in0 => \N__28581\,
            in1 => \N__28731\,
            in2 => \N__28346\,
            in3 => \N__28412\,
            lcout => \b2v_inst11.N_375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_sx_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__28732\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28336\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_sxZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__27026\,
            in1 => \N__27108\,
            in2 => \N__24487\,
            in3 => \N__24469\,
            lcout => \b2v_inst11.un1_clk_100khz_52_and_i_a2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNINJ641_0_2_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__27107\,
            in1 => \N__27027\,
            in2 => \N__24481\,
            in3 => \N__24427\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIVFCT3_1_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111010101010"
        )
    port map (
            in0 => \N__24892\,
            in1 => \N__24886\,
            in2 => \N__24877\,
            in3 => \N__29653\,
            lcout => \b2v_inst11.N_183\,
            ltout => \b2v_inst11.N_183_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIG8JO1_1_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001111"
        )
    port map (
            in0 => \N__29654\,
            in1 => \N__24867\,
            in2 => \N__24838\,
            in3 => \N__24675\,
            lcout => \b2v_inst11.N_114_f0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_3_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__29268\,
            in1 => \N__25552\,
            in2 => \N__25337\,
            in3 => \N__24820\,
            lcout => \b2v_inst11.g1_4_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_1_ss0_i_0_a2_3_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__28707\,
            in1 => \N__28252\,
            in2 => \_gnd_net_\,
            in3 => \N__29095\,
            lcout => \b2v_inst11.N_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst31.un8_output_0_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__29659\,
            in1 => \N__34743\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst31.un8_outputZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNI8OKQ2_0_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__29510\,
            in1 => \N__27843\,
            in2 => \_gnd_net_\,
            in3 => \N__33713\,
            lcout => \b2v_inst6.curr_state_RNI8OKQ2Z0Z_0\,
            ltout => \b2v_inst6.curr_state_RNI8OKQ2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_RNITH2G3_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__24600\,
            in1 => \N__29511\,
            in2 => \N__24697\,
            in3 => \N__29475\,
            lcout => \b2v_inst6.delayed_vccin_vccinaux_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_1_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__24624\,
            in1 => \N__27624\,
            in2 => \N__24689\,
            in3 => \N__24652\,
            lcout => \b2v_inst11.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34670\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__24610\,
            in1 => \N__29513\,
            in2 => \N__24604\,
            in3 => \N__29476\,
            lcout => \b2v_inst6.delayed_vccin_vccinaux_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34670\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33929\,
            in2 => \_gnd_net_\,
            in3 => \N__26877\,
            lcout => \SYNTHESIZED_WIRE_47keep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34670\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNI7OBF3_0_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100000"
        )
    port map (
            in0 => \N__33712\,
            in1 => \N__29512\,
            in2 => \N__27844\,
            in3 => \N__35178\,
            lcout => \b2v_inst6.count_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un1_vddq_en_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25055\,
            in2 => \_gnd_net_\,
            in3 => \N__25006\,
            lcout => \VDDQ_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst31.un8_output_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24982\,
            in1 => \N__24976\,
            in2 => \N__24970\,
            in3 => \N__24961\,
            lcout => \VCCIN_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_1_c_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32245\,
            in2 => \N__29818\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_1_0_\,
            carryout => \b2v_inst36.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29967\,
            in2 => \_gnd_net_\,
            in3 => \N__24931\,
            lcout => \b2v_inst36.un2_count_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_1\,
            carryout => \b2v_inst36.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29905\,
            in2 => \_gnd_net_\,
            in3 => \N__24928\,
            lcout => \b2v_inst36.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_2\,
            carryout => \b2v_inst36.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_3_c_RNICUC8_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__32214\,
            in1 => \N__30442\,
            in2 => \_gnd_net_\,
            in3 => \N__24925\,
            lcout => \b2v_inst36.count_rst_10\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_3\,
            carryout => \b2v_inst36.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24917\,
            in2 => \_gnd_net_\,
            in3 => \N__24895\,
            lcout => \b2v_inst36.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_4\,
            carryout => \b2v_inst36.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_5_c_RNINEG01_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__32215\,
            in1 => \N__29770\,
            in2 => \_gnd_net_\,
            in3 => \N__25183\,
            lcout => \b2v_inst36.count_rst_8\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_5\,
            carryout => \b2v_inst36.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25172\,
            in2 => \_gnd_net_\,
            in3 => \N__25141\,
            lcout => \b2v_inst36.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_6\,
            carryout => \b2v_inst36.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29858\,
            in2 => \_gnd_net_\,
            in3 => \N__25123\,
            lcout => \b2v_inst36.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_7\,
            carryout => \b2v_inst36.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_8_c_RNIH8I8_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31552\,
            in3 => \N__25120\,
            lcout => \b2v_inst36.un2_count_1_cry_8_c_RNIH8IZ0Z8\,
            ltout => OPEN,
            carryin => \bfn_9_2_0_\,
            carryout => \b2v_inst36.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29834\,
            in2 => \_gnd_net_\,
            in3 => \N__25108\,
            lcout => \b2v_inst36.un2_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_9\,
            carryout => \b2v_inst36.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29745\,
            in2 => \_gnd_net_\,
            in3 => \N__25105\,
            lcout => \b2v_inst36.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_10\,
            carryout => \b2v_inst36.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_11_c_RNIR5K1_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__32199\,
            in1 => \N__30027\,
            in2 => \_gnd_net_\,
            in3 => \N__25102\,
            lcout => \b2v_inst36.count_rst_2\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_11\,
            carryout => \b2v_inst36.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_12_c_RNIS7L1_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31569\,
            in2 => \_gnd_net_\,
            in3 => \N__25099\,
            lcout => \b2v_inst36.un2_count_1_cry_12_c_RNIS7LZ0Z1\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_12\,
            carryout => \b2v_inst36.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_13_c_RNIT9M1_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__32200\,
            in1 => \N__29430\,
            in2 => \_gnd_net_\,
            in3 => \N__25246\,
            lcout => \b2v_inst36.count_rst_0\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_13\,
            carryout => \b2v_inst36.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_14_c_RNIUBN1_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__29415\,
            in1 => \N__32201\,
            in2 => \_gnd_net_\,
            in3 => \N__25243\,
            lcout => \b2v_inst36.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNILPEV_14_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25210\,
            in1 => \N__31915\,
            in2 => \_gnd_net_\,
            in3 => \N__25221\,
            lcout => \b2v_inst36.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_12_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25231\,
            lcout => \b2v_inst36.count_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34677\,
            ce => \N__31958\,
            sr => \N__31835\
        );

    \b2v_inst36.curr_state_RNIKEBL_1_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__31800\,
            in1 => \N__30259\,
            in2 => \N__30357\,
            in3 => \N__33716\,
            lcout => \b2v_inst36.count_en\,
            ltout => \b2v_inst36.count_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIHJCV_12_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25240\,
            in2 => \N__25234\,
            in3 => \N__25230\,
            lcout => \b2v_inst36.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_14_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25222\,
            lcout => \b2v_inst36.count_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34677\,
            ce => \N__31958\,
            sr => \N__31835\
        );

    \b2v_inst36.count_15_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25197\,
            lcout => \b2v_inst36.count_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34677\,
            ce => \N__31958\,
            sr => \N__31835\
        );

    \b2v_inst36.count_RNINSFV_15_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31959\,
            in1 => \_gnd_net_\,
            in2 => \N__25201\,
            in3 => \N__25189\,
            lcout => \b2v_inst36.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_4_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30462\,
            lcout => \b2v_inst36.count_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34677\,
            ce => \N__31958\,
            sr => \N__31835\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25590\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_4_0_\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25439\,
            in2 => \N__25255\,
            in3 => \N__25466\,
            lcout => \G_2890\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_0\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25492\,
            in2 => \N__25444\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_1\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25467\,
            in2 => \N__25486\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25477\,
            in2 => \N__25471\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25443\,
            in2 => \N__25429\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__25417\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25411\,
            lcout => \b2v_inst11.un85_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__25396\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.pwm_out_RNO_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__25663\,
            in1 => \N__34092\,
            in2 => \_gnd_net_\,
            in3 => \N__25679\,
            lcout => \b2v_inst11.pwm_out_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_2_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__25919\,
            in1 => \N__25616\,
            in2 => \_gnd_net_\,
            in3 => \N__26021\,
            lcout => \b2v_inst11.un79_clk_100khzlt6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_15_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__25889\,
            in1 => \N__26403\,
            in2 => \_gnd_net_\,
            in3 => \N__25862\,
            lcout => \b2v_inst11.un79_clk_100khzlto15_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_9_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25842\,
            in1 => \N__25815\,
            in2 => \N__26365\,
            in3 => \N__25789\,
            lcout => OPEN,
            ltout => \b2v_inst11.un79_clk_100khzlto15_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_5_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__25765\,
            in1 => \N__25757\,
            in2 => \N__25738\,
            in3 => \N__25979\,
            lcout => OPEN,
            ltout => \b2v_inst11.un79_clk_100khzlto15_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_13_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__25730\,
            in1 => \N__26066\,
            in2 => \N__25711\,
            in3 => \N__25708\,
            lcout => \b2v_inst11.count_RNIZ0Z_13\,
            ltout => \b2v_inst11.count_RNIZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.pwm_out_RNO_1_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100010001"
        )
    port map (
            in0 => \N__25662\,
            in1 => \N__26610\,
            in2 => \N__25627\,
            in3 => \N__34093\,
            lcout => \b2v_inst11.g0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIMQBN_3_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34076\,
            in1 => \N__26077\,
            in2 => \_gnd_net_\,
            in3 => \N__26085\,
            lcout => \b2v_inst11.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_3_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26086\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34662\,
            ce => \N__33688\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIOC3M_13_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34079\,
            in1 => \N__26035\,
            in2 => \_gnd_net_\,
            in3 => \N__26043\,
            lcout => \b2v_inst11.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_13_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26047\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34662\,
            ce => \N__33688\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIOTCN_4_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34077\,
            in1 => \N__25993\,
            in2 => \_gnd_net_\,
            in3 => \N__26001\,
            lcout => \b2v_inst11.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_4_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26002\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34662\,
            ce => \N__33688\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIQ0EN_5_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34078\,
            in1 => \N__25951\,
            in2 => \_gnd_net_\,
            in3 => \N__25959\,
            lcout => \b2v_inst11.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_5_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25960\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34662\,
            ce => \N__33688\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI03G9_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25945\,
            in1 => \N__34086\,
            in2 => \_gnd_net_\,
            in3 => \N__25933\,
            lcout => \b2v_inst11.countZ0Z_0\,
            ltout => \b2v_inst11.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__26555\,
            in1 => \_gnd_net_\,
            in2 => \N__25924\,
            in3 => \N__26486\,
            lcout => OPEN,
            ltout => \b2v_inst11.count_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI14G9_1_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26413\,
            in2 => \N__26566\,
            in3 => \N__34087\,
            lcout => \b2v_inst11.countZ0Z_1\,
            ltout => \b2v_inst11.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_1_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26518\,
            in2 => \N__26494\,
            in3 => \N__26487\,
            lcout => \b2v_inst11.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34655\,
            ce => \N__33685\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI0AHN_8_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26371\,
            in1 => \N__34088\,
            in2 => \_gnd_net_\,
            in3 => \N__26379\,
            lcout => \b2v_inst11.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_8_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26380\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34655\,
            ce => \N__33685\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI2DIN_9_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26320\,
            in1 => \N__34089\,
            in2 => \_gnd_net_\,
            in3 => \N__26328\,
            lcout => \b2v_inst11.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_9_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26329\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34655\,
            ce => \N__33685\,
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNI65HI_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26266\,
            in1 => \N__26314\,
            in2 => \_gnd_net_\,
            in3 => \N__34090\,
            lcout => \b2v_inst5.curr_stateZ0Z_0\,
            ltout => \b2v_inst5.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_7_1_0__m4_0_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001010"
        )
    port map (
            in0 => \N__26284\,
            in1 => \_gnd_net_\,
            in2 => \N__26269\,
            in3 => \N__27089\,
            lcout => \b2v_inst5.m4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNITBKN1_7_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__27088\,
            in1 => \N__26260\,
            in2 => \_gnd_net_\,
            in3 => \N__26233\,
            lcout => \b2v_inst11.dutycycle_RNITBKN1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_en_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26667\,
            in2 => \_gnd_net_\,
            in3 => \N__27593\,
            lcout => \b2v_inst5.count_enZ0\,
            ltout => \b2v_inst5.count_enZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNICVEB2_6_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__30676\,
            in1 => \N__30745\,
            in2 => \N__26656\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.un2_count_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.pwm_out_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101010"
        )
    port map (
            in0 => \N__26606\,
            in1 => \N__27594\,
            in2 => \N__26653\,
            in3 => \N__26620\,
            lcout => \b2v_inst11.pwm_outZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34651\,
            ce => 'H',
            sr => \N__26587\
        );

    \b2v_inst5.count_RNIE2GB2_7_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30214\,
            in1 => \N__32546\,
            in2 => \_gnd_net_\,
            in3 => \N__30868\,
            lcout => \b2v_inst5.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIA2IH2_14_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32547\,
            in1 => \N__30229\,
            in2 => \_gnd_net_\,
            in3 => \N__30774\,
            lcout => \b2v_inst5.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_0_c_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26575\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \b2v_inst20.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_1_c_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26689\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_0\,
            carryout => \b2v_inst20.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_2_c_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33370\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_1\,
            carryout => \b2v_inst20.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_3_c_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33304\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_2\,
            carryout => \b2v_inst20.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_4_c_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33241\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_3\,
            carryout => \b2v_inst20.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_5_c_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33175\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_4\,
            carryout => \b2v_inst20.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_6_c_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33100\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_5\,
            carryout => \b2v_inst20.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_7_c_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33433\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_6\,
            carryout => b2v_inst20_un4_counter_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26692\,
            lcout => \b2v_inst20_un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_6_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26848\,
            in1 => \N__30929\,
            in2 => \_gnd_net_\,
            in3 => \N__30913\,
            lcout => \b2v_inst20.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_2_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__31063\,
            in1 => \N__31083\,
            in2 => \_gnd_net_\,
            in3 => \N__26849\,
            lcout => \b2v_inst20.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_5_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30966\,
            in2 => \N__26867\,
            in3 => \N__30952\,
            lcout => \b2v_inst20.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_1_c_RNO_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__30965\,
            in1 => \N__31136\,
            in2 => \N__30933\,
            in3 => \N__31231\,
            lcout => \b2v_inst20.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.SYNTHESIZED_WIRE_48_i_0_o3_2_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101011111"
        )
    port map (
            in0 => \N__28348\,
            in1 => \N__27087\,
            in2 => \N__27025\,
            in3 => \N__26923\,
            lcout => \SYNTHESIZED_WIRE_48_i_0_o3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__31140\,
            in1 => \N__26844\,
            in2 => \_gnd_net_\,
            in3 => \N__31112\,
            lcout => \b2v_inst20.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_3_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26843\,
            in1 => \N__31021\,
            in2 => \_gnd_net_\,
            in3 => \N__31043\,
            lcout => \b2v_inst20.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_5_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28434\,
            in1 => \N__26742\,
            in2 => \_gnd_net_\,
            in3 => \N__29285\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_234_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIG8JO1_5_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001111"
        )
    port map (
            in0 => \N__29072\,
            in1 => \N__27442\,
            in2 => \N__26971\,
            in3 => \N__29639\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_clk_100khz_52_and_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI8S5P2_5_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29615\,
            in2 => \N__26968\,
            in3 => \N__28575\,
            lcout => \b2v_inst11.g2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_rep1_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26851\,
            in2 => \_gnd_net_\,
            in3 => \N__26942\,
            lcout => \SYNTHESIZED_WIRE_47keep_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26850\,
            in2 => \_gnd_net_\,
            in3 => \N__31113\,
            lcout => \b2v_inst20.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_S4n_ibuf_RNINJ641_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__27118\,
            in1 => \N__29093\,
            in2 => \N__26764\,
            in3 => \N__28830\,
            lcout => \G_26_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_9_4_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__28831\,
            in1 => \N__28762\,
            in2 => \_gnd_net_\,
            in3 => \N__27331\,
            lcout => OPEN,
            ltout => \G_26_0_a5_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_S4n_ibuf_RNIE7D82_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100100"
        )
    port map (
            in0 => \N__27832\,
            in1 => \N__27826\,
            in2 => \N__27820\,
            in3 => \N__27817\,
            lcout => OPEN,
            ltout => \b2v_inst11_un1_dutycycle_172_m3_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIL3755_0_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101111111111"
        )
    port map (
            in0 => \N__27811\,
            in1 => \N__27799\,
            in2 => \N__27793\,
            in3 => \N__29619\,
            lcout => OPEN,
            ltout => \b2v_inst11.g4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIM0L9A_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011111111"
        )
    port map (
            in0 => \N__27790\,
            in1 => \N__27695\,
            in2 => \N__27628\,
            in3 => \N__27545\,
            lcout => \b2v_inst11.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_x_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28745\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28332\,
            lcout => \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_xZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_2_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__27390\,
            in1 => \N__28761\,
            in2 => \_gnd_net_\,
            in3 => \N__27330\,
            lcout => \N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNINJ641_6_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__28031\,
            in1 => \N__27311\,
            in2 => \_gnd_net_\,
            in3 => \N__28165\,
            lcout => \b2v_inst11.g3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_S4n_ibuf_RNIF6NL_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__28309\,
            in1 => \N__28705\,
            in2 => \N__28837\,
            in3 => \N__27124\,
            lcout => \G_26_0_a5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIE5T11_6_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000101"
        )
    port map (
            in0 => \N__28029\,
            in1 => \N__29354\,
            in2 => \N__29293\,
            in3 => \N__28592\,
            lcout => OPEN,
            ltout => \b2v_inst11.g2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI2C4V3_6_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__29128\,
            in1 => \N__27862\,
            in2 => \N__29122\,
            in3 => \N__29094\,
            lcout => \b2v_inst11.N_228_N_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_RNIM6F44_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29011\,
            in2 => \_gnd_net_\,
            in3 => \N__29638\,
            lcout => \N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_4_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__28166\,
            in1 => \N__29002\,
            in2 => \N__28995\,
            in3 => \N__28836\,
            lcout => \b2v_inst11.g0_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIE5T11_0_1_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000001010"
        )
    port map (
            in0 => \N__28706\,
            in1 => \N__28593\,
            in2 => \N__28433\,
            in3 => \N__28311\,
            lcout => OPEN,
            ltout => \b2v_inst11.g1_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIL5HA1_6_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010111111111"
        )
    port map (
            in0 => \N__28310\,
            in1 => \N__28167\,
            in2 => \N__28039\,
            in3 => \N__28030\,
            lcout => \b2v_inst11.g1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIRLUM4_11_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34346\,
            in1 => \N__27850\,
            in2 => \_gnd_net_\,
            in3 => \N__29395\,
            lcout => \b2v_inst6.countZ0Z_11\,
            ltout => \b2v_inst6.countZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_11_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__35203\,
            in1 => \N__34939\,
            in2 => \N__27853\,
            in3 => \N__31297\,
            lcout => \b2v_inst6.count_3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34671\,
            ce => \N__34429\,
            sr => \N__35270\
        );

    \b2v_inst6.curr_state_RNIDMSJ1_1_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__29706\,
            in1 => \N__29536\,
            in2 => \N__29670\,
            in3 => \N__29722\,
            lcout => \b2v_inst6.curr_state_RNIDMSJ1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_10_c_RNI6P001_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__35202\,
            in1 => \N__34937\,
            in2 => \N__31488\,
            in3 => \N__31296\,
            lcout => \b2v_inst6.count_rst_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_3_c_RNIO6IO_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__34936\,
            in1 => \N__31332\,
            in2 => \N__35054\,
            in3 => \N__35201\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIVJVD4_4_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29383\,
            in2 => \N__29389\,
            in3 => \N__34345\,
            lcout => \b2v_inst6.countZ0Z_4\,
            ltout => \b2v_inst6.countZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_4_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__34938\,
            in1 => \N__31333\,
            in2 => \N__29386\,
            in3 => \N__35205\,
            lcout => \b2v_inst6.count_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34671\,
            ce => \N__34429\,
            sr => \N__35270\
        );

    \b2v_inst6.count_5_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__35204\,
            in1 => \N__34940\,
            in2 => \N__31378\,
            in3 => \N__35131\,
            lcout => \b2v_inst6.count_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34671\,
            ce => \N__34429\,
            sr => \N__35270\
        );

    \b2v_inst6.curr_state_RNIVVMK_0_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__29472\,
            in1 => \N__29505\,
            in2 => \_gnd_net_\,
            in3 => \N__33906\,
            lcout => \b2v_inst6.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_7_1_0__m4_0_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000001000"
        )
    port map (
            in0 => \N__29533\,
            in1 => \N__34960\,
            in2 => \N__29515\,
            in3 => \N__29471\,
            lcout => OPEN,
            ltout => \G_2746_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNI7JCH_0_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29371\,
            in2 => \N__29377\,
            in3 => \N__33905\,
            lcout => \b2v_inst6.curr_stateZ0Z_0\,
            ltout => \b2v_inst6.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_0_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000001000"
        )
    port map (
            in0 => \N__29534\,
            in1 => \N__34959\,
            in2 => \N__29374\,
            in3 => \N__29473\,
            lcout => \b2v_inst6.curr_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34676\,
            ce => \N__33678\,
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIDMSJ1_0_1_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__29721\,
            in1 => \N__29532\,
            in2 => \N__29707\,
            in3 => \N__29658\,
            lcout => \b2v_inst6.N_413\,
            ltout => \b2v_inst6.N_413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_7_1_0__m6_0_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__29535\,
            in1 => \N__34942\,
            in2 => \N__29542\,
            in3 => \N__29514\,
            lcout => OPEN,
            ltout => \b2v_inst6.curr_state_7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIF7P21_1_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29452\,
            in2 => \N__29539\,
            in3 => \N__33904\,
            lcout => \b2v_inst6.curr_stateZ0Z_1\,
            ltout => \b2v_inst6.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_1_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101000000"
        )
    port map (
            in0 => \N__29506\,
            in1 => \N__34941\,
            in2 => \N__29479\,
            in3 => \N__29474\,
            lcout => \b2v_inst6.curr_state_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34676\,
            ce => \N__33678\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI471O_1_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29401\,
            in1 => \N__31960\,
            in2 => \_gnd_net_\,
            in3 => \N__29443\,
            lcout => \b2v_inst36.countZ0Z_1\,
            ltout => \b2v_inst36.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI_1_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__32236\,
            in1 => \_gnd_net_\,
            in2 => \N__29446\,
            in3 => \N__32143\,
            lcout => \b2v_inst36.count_rst_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI_15_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29437\,
            in1 => \N__32235\,
            in2 => \N__31570\,
            in3 => \N__29419\,
            lcout => \b2v_inst36.un12_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_1_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__32237\,
            in1 => \N__29810\,
            in2 => \_gnd_net_\,
            in3 => \N__32146\,
            lcout => \b2v_inst36.count_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34689\,
            ce => \N__31962\,
            sr => \N__31828\
        );

    \b2v_inst36.un2_count_1_cry_1_c_RNIAQA8_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__32144\,
            in1 => \N__32038\,
            in2 => \N__29941\,
            in3 => \N__29963\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIF2C01_2_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31961\,
            in1 => \_gnd_net_\,
            in2 => \N__29971\,
            in3 => \N__29920\,
            lcout => \b2v_inst36.countZ0Z_2\,
            ltout => \b2v_inst36.countZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_2_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__32145\,
            in1 => \N__32042\,
            in2 => \N__29944\,
            in3 => \N__29940\,
            lcout => \b2v_inst36.count_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34689\,
            ce => \N__31962\,
            sr => \N__31828\
        );

    \b2v_inst36.count_3_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000000000"
        )
    port map (
            in0 => \N__29913\,
            in1 => \N__29887\,
            in2 => \N__32056\,
            in3 => \N__32147\,
            lcout => \b2v_inst36.count_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34689\,
            ce => \N__31962\,
            sr => \N__31828\
        );

    \b2v_inst36.count_RNI_0_1_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__29863\,
            in1 => \N__29842\,
            in2 => \N__29817\,
            in3 => \N__29741\,
            lcout => OPEN,
            ltout => \b2v_inst36.un12_clk_100khz_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI9C1O_2_6_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29791\,
            in1 => \N__30013\,
            in2 => \N__29779\,
            in3 => \N__29776\,
            lcout => \b2v_inst36.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_6_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30060\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.count_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34687\,
            ce => \N__31977\,
            sr => \N__31815\
        );

    \b2v_inst36.count_RNI9C1O_6_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30042\,
            in1 => \N__31964\,
            in2 => \_gnd_net_\,
            in3 => \N__30059\,
            lcout => \b2v_inst36.un2_count_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIFGBV_11_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31965\,
            in1 => \N__30070\,
            in2 => \_gnd_net_\,
            in3 => \N__29758\,
            lcout => \b2v_inst36.countZ0Z_11\,
            ltout => \b2v_inst36.countZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_11_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__30091\,
            in1 => \N__32182\,
            in2 => \N__30073\,
            in3 => \N__32054\,
            lcout => \b2v_inst36.count_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34687\,
            ce => \N__31977\,
            sr => \N__31815\
        );

    \b2v_inst36.count_RNI9C1O_0_6_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31966\,
            in1 => \_gnd_net_\,
            in2 => \N__30064\,
            in3 => \N__30043\,
            lcout => OPEN,
            ltout => \b2v_inst36.countZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI9C1O_1_6_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30034\,
            in1 => \N__31548\,
            in2 => \N__30016\,
            in3 => \N__30441\,
            lcout => \b2v_inst36.un12_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNI3NTL_1_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29983\,
            in1 => \N__29977\,
            in2 => \_gnd_net_\,
            in3 => \N__34073\,
            lcout => \b2v_inst36.curr_stateZ0Z_1\,
            ltout => \b2v_inst36.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_7_1_0__m4_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100000001000"
        )
    port map (
            in0 => \N__30301\,
            in1 => \N__30389\,
            in2 => \N__30007\,
            in3 => \N__32034\,
            lcout => OPEN,
            ltout => \b2v_inst36.curr_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNI2MTL_0_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30364\,
            in2 => \N__30004\,
            in3 => \N__34074\,
            lcout => \b2v_inst36.curr_stateZ0Z_0\,
            ltout => \b2v_inst36.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.DSW_PWROK_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000100000"
        )
    port map (
            in0 => \N__30298\,
            in1 => \N__30336\,
            in2 => \N__30001\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.DSW_PWROK_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34684\,
            ce => \N__33689\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_1_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101000100000"
        )
    port map (
            in0 => \N__30257\,
            in1 => \N__32052\,
            in2 => \N__30349\,
            in3 => \N__30300\,
            lcout => \b2v_inst36.curr_state_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34684\,
            ce => \N__33689\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_7_1_0__m6_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001000"
        )
    port map (
            in0 => \N__30302\,
            in1 => \N__30258\,
            in2 => \N__30353\,
            in3 => \N__32033\,
            lcout => \b2v_inst36.curr_state_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_0_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__30335\,
            in1 => \N__30299\,
            in2 => \N__32055\,
            in3 => \N__30388\,
            lcout => \b2v_inst36.curr_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34684\,
            ce => \N__33689\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNI0A86_1_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__34075\,
            in1 => \N__30334\,
            in2 => \N__30307\,
            in3 => \N__30256\,
            lcout => \b2v_inst36.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_14_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30775\,
            lcout => \b2v_inst5.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34679\,
            ce => \N__32686\,
            sr => \N__32867\
        );

    \b2v_inst5.count_6_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30669\,
            lcout => \b2v_inst5.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34679\,
            ce => \N__32686\,
            sr => \N__32867\
        );

    \b2v_inst5.count_7_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30867\,
            lcout => \b2v_inst5.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34679\,
            ce => \N__32686\,
            sr => \N__32867\
        );

    \b2v_inst16.count_RNIPM3K1_8_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30174\,
            in1 => \N__30157\,
            in2 => \_gnd_net_\,
            in3 => \N__30603\,
            lcout => \b2v_inst16.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_8_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30175\,
            lcout => \b2v_inst16.count_4_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34672\,
            ce => \N__30604\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIRP4K1_9_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30118\,
            in1 => \N__30097\,
            in2 => \_gnd_net_\,
            in3 => \N__30602\,
            lcout => \b2v_inst16.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_9_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30117\,
            lcout => \b2v_inst16.count_4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34672\,
            ce => \N__30604\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIJ8E01_4_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30475\,
            in1 => \N__31963\,
            in2 => \_gnd_net_\,
            in3 => \N__30463\,
            lcout => \b2v_inst36.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI_0_0_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32332\,
            lcout => \b2v_inst5.N_2906_i\,
            ltout => \b2v_inst5.N_2906_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIU55SG_2_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__32443\,
            in1 => \_gnd_net_\,
            in2 => \N__30424\,
            in3 => \N__32302\,
            lcout => \b2v_inst5.N_390\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIC5JH2_15_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32642\,
            in1 => \N__31153\,
            in2 => \_gnd_net_\,
            in3 => \N__31168\,
            lcout => \b2v_inst5.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_12_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30820\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34666\,
            ce => \N__32680\,
            sr => \N__32893\
        );

    \b2v_inst5.count_RNI6SFH2_12_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30417\,
            in1 => \N__32637\,
            in2 => \_gnd_net_\,
            in3 => \N__30818\,
            lcout => \b2v_inst5.un2_count_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIASDB2_0_5_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__32681\,
            in1 => \N__30754\,
            in2 => \N__30799\,
            in3 => \N__30703\,
            lcout => OPEN,
            ltout => \b2v_inst5.count_1_i_a2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNISNC87_5_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30724\,
            in1 => \N__32509\,
            in2 => \N__30421\,
            in3 => \N__30409\,
            lcout => \b2v_inst5.count_1_i_a2_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI6SFH2_0_12_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010011"
        )
    port map (
            in0 => \N__30819\,
            in1 => \N__30418\,
            in2 => \N__32664\,
            in3 => \N__31182\,
            lcout => \b2v_inst5.count_1_i_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_5_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30702\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34666\,
            ce => \N__32680\,
            sr => \N__32893\
        );

    \b2v_inst5.count_RNIASDB2_5_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32641\,
            in1 => \N__30753\,
            in2 => \_gnd_net_\,
            in3 => \N__30701\,
            lcout => \b2v_inst5.un2_count_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNICVEB2_0_6_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001101"
        )
    port map (
            in0 => \N__30744\,
            in1 => \N__32682\,
            in2 => \N__30895\,
            in3 => \N__30665\,
            lcout => \b2v_inst5.count_1_i_a2_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_1_c_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32331\,
            in2 => \N__32398\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \b2v_inst5.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_1_c_RNIJQ1L1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32808\,
            in1 => \N__32404\,
            in2 => \_gnd_net_\,
            in3 => \N__30718\,
            lcout => \b2v_inst5.count_rst_12\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_1\,
            carryout => \b2v_inst5.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32469\,
            in2 => \_gnd_net_\,
            in3 => \N__30715\,
            lcout => \b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_2\,
            carryout => \b2v_inst5.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32997\,
            in2 => \_gnd_net_\,
            in3 => \N__30712\,
            lcout => \b2v_inst5.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_3\,
            carryout => \b2v_inst5.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_4_c_RNIM05L1_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32803\,
            in1 => \N__30709\,
            in2 => \_gnd_net_\,
            in3 => \N__30691\,
            lcout => \b2v_inst5.count_rst_9\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_4\,
            carryout => \b2v_inst5.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_5_c_RNIN26L1_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32809\,
            in1 => \N__30688\,
            in2 => \_gnd_net_\,
            in3 => \N__30646\,
            lcout => \b2v_inst5.count_rst_8\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_5\,
            carryout => \b2v_inst5.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_6_c_RNIO47L1_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32802\,
            in1 => \N__30891\,
            in2 => \_gnd_net_\,
            in3 => \N__30847\,
            lcout => \b2v_inst5.count_rst_7\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_6\,
            carryout => \b2v_inst5.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33046\,
            in2 => \_gnd_net_\,
            in3 => \N__30844\,
            lcout => \b2v_inst5.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_7\,
            carryout => \b2v_inst5.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31750\,
            in2 => \_gnd_net_\,
            in3 => \N__30841\,
            lcout => \b2v_inst5.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \b2v_inst5.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31705\,
            in2 => \_gnd_net_\,
            in3 => \N__30838\,
            lcout => \b2v_inst5.un2_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_9\,
            carryout => \b2v_inst5.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_10_c_RNI3GUD1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32804\,
            in1 => \N__32347\,
            in2 => \_gnd_net_\,
            in3 => \N__30835\,
            lcout => \b2v_inst5.count_rst_3\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_10\,
            carryout => \b2v_inst5.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_11_c_RNI4IVD1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__32806\,
            in1 => \_gnd_net_\,
            in2 => \N__30832\,
            in3 => \N__30805\,
            lcout => \b2v_inst5.count_rst_2\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_11\,
            carryout => \b2v_inst5.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32500\,
            in2 => \_gnd_net_\,
            in3 => \N__30802\,
            lcout => \b2v_inst5.un2_count_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_12\,
            carryout => \b2v_inst5.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_13_c_RNI6M1E1_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32807\,
            in1 => \N__30792\,
            in2 => \_gnd_net_\,
            in3 => \N__30757\,
            lcout => \b2v_inst5.count_rst_0\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_13\,
            carryout => \b2v_inst5.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_14_c_RNI7O2E1_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32805\,
            in1 => \N__31186\,
            in2 => \_gnd_net_\,
            in3 => \N__31171\,
            lcout => \b2v_inst5.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_15_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31167\,
            lcout => \b2v_inst5.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34658\,
            ce => \N__32679\,
            sr => \N__32880\
        );

    \b2v_inst20.counter_1_cry_1_c_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31144\,
            in2 => \N__31120\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \b2v_inst20.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31087\,
            in2 => \_gnd_net_\,
            in3 => \N__31051\,
            lcout => \b2v_inst20.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_1\,
            carryout => \b2v_inst20.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31048\,
            in2 => \_gnd_net_\,
            in3 => \N__31009\,
            lcout => \b2v_inst20.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_2\,
            carryout => \b2v_inst20.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31006\,
            in2 => \_gnd_net_\,
            in3 => \N__30976\,
            lcout => \b2v_inst20.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_3\,
            carryout => \b2v_inst20.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30973\,
            in2 => \_gnd_net_\,
            in3 => \N__30940\,
            lcout => \b2v_inst20.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_4\,
            carryout => \b2v_inst20.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30937\,
            in2 => \_gnd_net_\,
            in3 => \N__30898\,
            lcout => \b2v_inst20.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_5\,
            carryout => \b2v_inst20.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_7_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31227\,
            in2 => \_gnd_net_\,
            in3 => \N__31213\,
            lcout => \b2v_inst20.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_6\,
            carryout => \b2v_inst20.counter_1_cry_7\,
            clk => \N__34652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_8_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33409\,
            in2 => \_gnd_net_\,
            in3 => \N__31210\,
            lcout => \b2v_inst20.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_7\,
            carryout => \b2v_inst20.counter_1_cry_8\,
            clk => \N__34652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_9_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33382\,
            in2 => \_gnd_net_\,
            in3 => \N__31207\,
            lcout => \b2v_inst20.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \b2v_inst20.counter_1_cry_9\,
            clk => \N__34657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_10_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33396\,
            in2 => \_gnd_net_\,
            in3 => \N__31204\,
            lcout => \b2v_inst20.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_9\,
            carryout => \b2v_inst20.counter_1_cry_10\,
            clk => \N__34657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_11_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33421\,
            in2 => \_gnd_net_\,
            in3 => \N__31201\,
            lcout => \b2v_inst20.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_10\,
            carryout => \b2v_inst20.counter_1_cry_11\,
            clk => \N__34657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_12_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33355\,
            in2 => \_gnd_net_\,
            in3 => \N__31198\,
            lcout => \b2v_inst20.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_11\,
            carryout => \b2v_inst20.counter_1_cry_12\,
            clk => \N__34657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_13_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33316\,
            in2 => \_gnd_net_\,
            in3 => \N__31195\,
            lcout => \b2v_inst20.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_12\,
            carryout => \b2v_inst20.counter_1_cry_13\,
            clk => \N__34657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_14_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33343\,
            in2 => \_gnd_net_\,
            in3 => \N__31192\,
            lcout => \b2v_inst20.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_13\,
            carryout => \b2v_inst20.counter_1_cry_14\,
            clk => \N__34657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_15_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33330\,
            in2 => \_gnd_net_\,
            in3 => \N__31189\,
            lcout => \b2v_inst20.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_14\,
            carryout => \b2v_inst20.counter_1_cry_15\,
            clk => \N__34657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_16_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33280\,
            in2 => \_gnd_net_\,
            in3 => \N__31258\,
            lcout => \b2v_inst20.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_15\,
            carryout => \b2v_inst20.counter_1_cry_16\,
            clk => \N__34657\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_17_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33267\,
            in2 => \_gnd_net_\,
            in3 => \N__31255\,
            lcout => \b2v_inst20.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \b2v_inst20.counter_1_cry_17\,
            clk => \N__34663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_18_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33253\,
            in2 => \_gnd_net_\,
            in3 => \N__31252\,
            lcout => \b2v_inst20.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_17\,
            carryout => \b2v_inst20.counter_1_cry_18\,
            clk => \N__34663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_19_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33292\,
            in2 => \_gnd_net_\,
            in3 => \N__31249\,
            lcout => \b2v_inst20.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_18\,
            carryout => \b2v_inst20.counter_1_cry_19\,
            clk => \N__34663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_20_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33187\,
            in2 => \_gnd_net_\,
            in3 => \N__31246\,
            lcout => \b2v_inst20.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_19\,
            carryout => \b2v_inst20.counter_1_cry_20\,
            clk => \N__34663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_21_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33201\,
            in2 => \_gnd_net_\,
            in3 => \N__31243\,
            lcout => \b2v_inst20.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_20\,
            carryout => \b2v_inst20.counter_1_cry_21\,
            clk => \N__34663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_22_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33214\,
            in2 => \_gnd_net_\,
            in3 => \N__31240\,
            lcout => \b2v_inst20.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_21\,
            carryout => \b2v_inst20.counter_1_cry_22\,
            clk => \N__34663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_23_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33226\,
            in2 => \_gnd_net_\,
            in3 => \N__31237\,
            lcout => \b2v_inst20.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_22\,
            carryout => \b2v_inst20.counter_1_cry_23\,
            clk => \N__34663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_24_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33160\,
            in2 => \_gnd_net_\,
            in3 => \N__31234\,
            lcout => \b2v_inst20.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_23\,
            carryout => \b2v_inst20.counter_1_cry_24\,
            clk => \N__34663\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_25_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33129\,
            in2 => \_gnd_net_\,
            in3 => \N__31282\,
            lcout => \b2v_inst20.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \b2v_inst20.counter_1_cry_25\,
            clk => \N__34665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_26_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33114\,
            in2 => \_gnd_net_\,
            in3 => \N__31279\,
            lcout => \b2v_inst20.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_25\,
            carryout => \b2v_inst20.counter_1_cry_26\,
            clk => \N__34665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_27_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33147\,
            in2 => \_gnd_net_\,
            in3 => \N__31276\,
            lcout => \b2v_inst20.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_26\,
            carryout => \b2v_inst20.counter_1_cry_27\,
            clk => \N__34665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_28_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33472\,
            in2 => \_gnd_net_\,
            in3 => \N__31273\,
            lcout => \b2v_inst20.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_27\,
            carryout => \b2v_inst20.counter_1_cry_28\,
            clk => \N__34665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_29_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33484\,
            in2 => \_gnd_net_\,
            in3 => \N__31270\,
            lcout => \b2v_inst20.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_28\,
            carryout => \b2v_inst20.counter_1_cry_29\,
            clk => \N__34665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_30_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33445\,
            in2 => \_gnd_net_\,
            in3 => \N__31267\,
            lcout => \b2v_inst20.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_29\,
            carryout => \b2v_inst20.counter_1_cry_30\,
            clk => \N__34665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_31_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33459\,
            in2 => \_gnd_net_\,
            in3 => \N__31264\,
            lcout => \b2v_inst20.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34665\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_1_c_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34214\,
            in2 => \N__35026\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \b2v_inst6.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_1_c_RNIM2GO_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35273\,
            in1 => \N__34230\,
            in2 => \_gnd_net_\,
            in3 => \N__31261\,
            lcout => \b2v_inst6.count_rst_1\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_1\,
            carryout => \b2v_inst6.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35093\,
            in2 => \_gnd_net_\,
            in3 => \N__31336\,
            lcout => \b2v_inst6.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_2\,
            carryout => \b2v_inst6.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35058\,
            in2 => \_gnd_net_\,
            in3 => \N__31318\,
            lcout => \b2v_inst6.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_3\,
            carryout => \b2v_inst6.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35126\,
            in2 => \_gnd_net_\,
            in3 => \N__31315\,
            lcout => \b2v_inst6.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_4\,
            carryout => \b2v_inst6.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_5_c_RNIQAKO_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35274\,
            in1 => \N__34255\,
            in2 => \_gnd_net_\,
            in3 => \N__31312\,
            lcout => \b2v_inst6.count_rst_5\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_5\,
            carryout => \b2v_inst6.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31455\,
            in2 => \_gnd_net_\,
            in3 => \N__31309\,
            lcout => \b2v_inst6.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_6\,
            carryout => \b2v_inst6.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31410\,
            in2 => \_gnd_net_\,
            in3 => \N__31306\,
            lcout => \b2v_inst6.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_7\,
            carryout => \b2v_inst6.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31633\,
            in2 => \_gnd_net_\,
            in3 => \N__31303\,
            lcout => \b2v_inst6.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \b2v_inst6.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_9_c_RNIUIOO_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35290\,
            in1 => \N__34242\,
            in2 => \_gnd_net_\,
            in3 => \N__31300\,
            lcout => \b2v_inst6.count_rst_9\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_9\,
            carryout => \b2v_inst6.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31484\,
            in2 => \_gnd_net_\,
            in3 => \N__31285\,
            lcout => \b2v_inst6.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_10\,
            carryout => \b2v_inst6.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_11_c_RNI7R101_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35291\,
            in1 => \N__34200\,
            in2 => \_gnd_net_\,
            in3 => \N__31390\,
            lcout => \b2v_inst6.count_rst_11\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_11\,
            carryout => \b2v_inst6.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_12_c_RNI8T201_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35296\,
            in1 => \N__34173\,
            in2 => \_gnd_net_\,
            in3 => \N__31387\,
            lcout => \b2v_inst6.count_rst_12\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_12\,
            carryout => \b2v_inst6.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_13_c_RNI9V301_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35292\,
            in1 => \N__34848\,
            in2 => \_gnd_net_\,
            in3 => \N__31384\,
            lcout => \b2v_inst6.count_rst_13\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_13\,
            carryout => \b2v_inst6.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_14_c_RNIA1501_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__34803\,
            in1 => \N__35293\,
            in2 => \_gnd_net_\,
            in3 => \N__31381\,
            lcout => \b2v_inst6.count_rst_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_15_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34816\,
            lcout => \b2v_inst6.count_3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34678\,
            ce => \N__34430\,
            sr => \N__35297\
        );

    \b2v_inst6.un2_count_1_cry_4_c_RNIP8JO_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__34895\,
            in1 => \N__31371\,
            in2 => \N__35130\,
            in3 => \N__35226\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI1N0E4_5_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34370\,
            in1 => \_gnd_net_\,
            in2 => \N__31354\,
            in3 => \N__31351\,
            lcout => \b2v_inst6.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_2_c_RNIN4HO_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__34894\,
            in1 => \N__34716\,
            in2 => \N__35095\,
            in3 => \N__35225\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNITGUD4_3_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34369\,
            in1 => \_gnd_net_\,
            in2 => \N__31339\,
            in3 => \N__34699\,
            lcout => \b2v_inst6.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_8_c_RNITGNO_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__34896\,
            in1 => \N__31611\,
            in2 => \N__31639\,
            in3 => \N__35227\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI935E4_9_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34371\,
            in1 => \_gnd_net_\,
            in2 => \N__31510\,
            in3 => \N__31600\,
            lcout => \b2v_inst6.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIIEMF4_10_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31498\,
            in1 => \N__31506\,
            in2 => \_gnd_net_\,
            in3 => \N__34372\,
            lcout => \b2v_inst6.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_10_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31507\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.count_3_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34683\,
            ce => \N__34420\,
            sr => \N__35294\
        );

    \b2v_inst6.count_RNI_7_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31406\,
            in1 => \N__31634\,
            in2 => \N__31456\,
            in3 => \N__31489\,
            lcout => \b2v_inst6.un12_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_6_c_RNIRCLO_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__31434\,
            in1 => \N__31454\,
            in2 => \N__34928\,
            in3 => \N__35275\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI5T2E4_7_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31420\,
            in2 => \N__31459\,
            in3 => \N__34418\,
            lcout => \b2v_inst6.countZ0Z_7\,
            ltout => \b2v_inst6.countZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_7_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__31435\,
            in1 => \N__34935\,
            in2 => \N__31423\,
            in3 => \N__35278\,
            lcout => \b2v_inst6.count_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34686\,
            ce => \N__34434\,
            sr => \N__35307\
        );

    \b2v_inst6.un2_count_1_cry_7_c_RNISEMO_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__35276\,
            in1 => \N__31656\,
            in2 => \N__31411\,
            in3 => \N__34903\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI704E4_8_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34419\,
            in1 => \_gnd_net_\,
            in2 => \N__31414\,
            in3 => \N__31645\,
            lcout => \b2v_inst6.countZ0Z_8\,
            ltout => \b2v_inst6.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_8_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__35277\,
            in1 => \N__34904\,
            in2 => \N__31660\,
            in3 => \N__31657\,
            lcout => \b2v_inst6.count_3_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34686\,
            ce => \N__34434\,
            sr => \N__35307\
        );

    \b2v_inst6.count_9_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__31635\,
            in1 => \N__31615\,
            in2 => \N__34929\,
            in3 => \N__35279\,
            lcout => \b2v_inst6.count_3_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34686\,
            ce => \N__34434\,
            sr => \N__35307\
        );

    \b2v_inst36.count_RNI_0_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__32241\,
            in1 => \N__32181\,
            in2 => \_gnd_net_\,
            in3 => \N__32051\,
            lcout => \b2v_inst36.count_rst_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNI_1_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31785\,
            lcout => \b2v_inst36.N_2928_i\,
            ltout => \b2v_inst36.N_2928_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_13_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__31582\,
            in1 => \_gnd_net_\,
            in2 => \N__31591\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.count_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34690\,
            ce => \N__31975\,
            sr => \N__31836\
        );

    \b2v_inst36.count_RNIJMDV_13_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__32178\,
            in1 => \N__31588\,
            in2 => \N__31978\,
            in3 => \N__31581\,
            lcout => \b2v_inst36.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNITNJ01_9_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__31516\,
            in1 => \N__31970\,
            in2 => \N__31534\,
            in3 => \N__32177\,
            lcout => \b2v_inst36.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_9_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32179\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31530\,
            lcout => \b2v_inst36.count_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34690\,
            ce => \N__31975\,
            sr => \N__31836\
        );

    \b2v_inst36.count_RNI361O_0_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31974\,
            in1 => \N__32251\,
            in2 => \_gnd_net_\,
            in3 => \N__31984\,
            lcout => \b2v_inst36.countZ0Z_0\,
            ltout => \b2v_inst36.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_0_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32180\,
            in2 => \N__32092\,
            in3 => \N__32053\,
            lcout => \b2v_inst36.count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34690\,
            ce => \N__31975\,
            sr => \N__31836\
        );

    \b2v_inst5.count_RNII8IB2_0_9_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__31697\,
            in1 => \N__31759\,
            in2 => \N__32678\,
            in3 => \N__31717\,
            lcout => \b2v_inst5.count_1_i_a2_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_8_c_RNIQ89L1_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__31731\,
            in1 => \N__31743\,
            in2 => \N__32883\,
            in3 => \N__32946\,
            lcout => \b2v_inst5.count_rst_5\,
            ltout => \b2v_inst5.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNII8IB2_9_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32650\,
            in2 => \N__31753\,
            in3 => \N__31716\,
            lcout => \b2v_inst5.un2_count_1_axb_9\,
            ltout => \b2v_inst5.un2_count_1_axb_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_9_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__31732\,
            in1 => \N__32866\,
            in2 => \N__31720\,
            in3 => \N__32950\,
            lcout => \b2v_inst5.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34681\,
            ce => \N__32660\,
            sr => \N__32892\
        );

    \b2v_inst5.un2_count_1_cry_9_c_RNIRAAL1_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__32947\,
            in1 => \N__32861\,
            in2 => \N__31704\,
            in3 => \N__31680\,
            lcout => OPEN,
            ltout => \b2v_inst5.count_rst_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIRIQO2_10_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__32651\,
            in1 => \_gnd_net_\,
            in2 => \N__31708\,
            in3 => \N__31666\,
            lcout => \b2v_inst5.countZ0Z_10\,
            ltout => \b2v_inst5.countZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_10_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__32948\,
            in1 => \N__32865\,
            in2 => \N__31684\,
            in3 => \N__31681\,
            lcout => \b2v_inst5.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34681\,
            ce => \N__32660\,
            sr => \N__32892\
        );

    \b2v_inst5.count_13_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__32504\,
            in1 => \N__32908\,
            in2 => \N__32884\,
            in3 => \N__32949\,
            lcout => \b2v_inst5.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34681\,
            ce => \N__32660\,
            sr => \N__32892\
        );

    \b2v_inst5.count_RNIRHC7I_2_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__32297\,
            in1 => \N__32442\,
            in2 => \N__32868\,
            in3 => \N__32284\,
            lcout => OPEN,
            ltout => \b2v_inst5.count_RNIRHC7IZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIA8LTI_0_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32275\,
            in2 => \N__32335\,
            in3 => \N__32643\,
            lcout => \b2v_inst5.countZ0Z_0\,
            ltout => \b2v_inst5.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI_0_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32320\,
            in3 => \N__32397\,
            lcout => \b2v_inst5.count_RNIZ0Z_0\,
            ltout => \b2v_inst5.count_RNIZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNID3G12_1_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__32832\,
            in1 => \N__32308\,
            in2 => \N__32317\,
            in3 => \N__32644\,
            lcout => \b2v_inst5.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_1_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32314\,
            in2 => \_gnd_net_\,
            in3 => \N__32834\,
            lcout => \b2v_inst5.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34674\,
            ce => \N__32646\,
            sr => \N__32882\
        );

    \b2v_inst5.count_3_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32828\,
            in2 => \_gnd_net_\,
            in3 => \N__32260\,
            lcout => \b2v_inst5.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34674\,
            ce => \N__32646\,
            sr => \N__32882\
        );

    \b2v_inst5.count_0_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__32298\,
            in1 => \N__32283\,
            in2 => \N__32869\,
            in3 => \N__32441\,
            lcout => \b2v_inst5.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34674\,
            ce => \N__32646\,
            sr => \N__32882\
        );

    \b2v_inst5.count_RNI6MBB2_3_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__32833\,
            in1 => \N__32645\,
            in2 => \N__32269\,
            in3 => \N__32259\,
            lcout => \b2v_inst5.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_2_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32416\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34668\,
            ce => \N__32635\,
            sr => \N__32885\
        );

    \b2v_inst5.count_RNI4JAB2_0_2_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__32633\,
            in1 => \N__32425\,
            in2 => \N__32473\,
            in3 => \N__32415\,
            lcout => OPEN,
            ltout => \b2v_inst5.count_1_i_a2_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI2EOJ9_2_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32455\,
            in1 => \N__32341\,
            in2 => \N__32446\,
            in3 => \N__32377\,
            lcout => \b2v_inst5.count_1_i_a2_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI4JAB2_2_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__32632\,
            in1 => \N__32424\,
            in2 => \_gnd_net_\,
            in3 => \N__32414\,
            lcout => \b2v_inst5.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI4PEH2_0_11_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100111"
        )
    port map (
            in0 => \N__32634\,
            in1 => \N__32358\,
            in2 => \N__32371\,
            in3 => \N__32396\,
            lcout => \b2v_inst5.count_1_i_a2_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_11_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32359\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34668\,
            ce => \N__32635\,
            sr => \N__32885\
        );

    \b2v_inst5.count_RNI4PEH2_11_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__32367\,
            in1 => \N__32631\,
            in2 => \_gnd_net_\,
            in3 => \N__32357\,
            lcout => \b2v_inst5.un2_count_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI8PCB2_0_4_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__33045\,
            in1 => \N__33010\,
            in2 => \N__32974\,
            in3 => \N__32636\,
            lcout => \b2v_inst5.count_1_i_a2_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_7_c_RNIP68L1_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__32953\,
            in1 => \N__33027\,
            in2 => \N__32870\,
            in3 => \N__33044\,
            lcout => OPEN,
            ltout => \b2v_inst5.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIG5HB2_8_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__32649\,
            in1 => \_gnd_net_\,
            in2 => \N__33049\,
            in3 => \N__33016\,
            lcout => \b2v_inst5.countZ0Z_8\,
            ltout => \b2v_inst5.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_8_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__32955\,
            in1 => \N__33028\,
            in2 => \N__33019\,
            in3 => \N__32841\,
            lcout => \b2v_inst5.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34664\,
            ce => \N__32659\,
            sr => \N__32881\
        );

    \b2v_inst5.un2_count_1_cry_3_c_RNILU3L1_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__32985\,
            in1 => \N__32951\,
            in2 => \N__33001\,
            in3 => \N__32835\,
            lcout => \b2v_inst5.count_rst_10\,
            ltout => \b2v_inst5.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI8PCB2_4_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32970\,
            in2 => \N__33004\,
            in3 => \N__32647\,
            lcout => \b2v_inst5.un2_count_1_axb_4\,
            ltout => \b2v_inst5.un2_count_1_axb_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_4_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__32986\,
            in1 => \N__32954\,
            in2 => \N__32977\,
            in3 => \N__32839\,
            lcout => \b2v_inst5.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34664\,
            ce => \N__32659\,
            sr => \N__32881\
        );

    \b2v_inst5.un2_count_1_cry_12_c_RNI5K0E1_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__32952\,
            in1 => \N__32904\,
            in2 => \N__32505\,
            in3 => \N__32840\,
            lcout => OPEN,
            ltout => \b2v_inst5.count_rst_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI8VGH2_13_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__32648\,
            in1 => \_gnd_net_\,
            in2 => \N__32521\,
            in3 => \N__32518\,
            lcout => \b2v_inst5.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_2_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34114\,
            lcout => \b2v_inst200.curr_state_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34656\,
            ce => \N__33686\,
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_2_c_RNO_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33420\,
            in1 => \N__33408\,
            in2 => \N__33397\,
            in3 => \N__33381\,
            lcout => \b2v_inst20.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_3_c_RNO_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33354\,
            in1 => \N__33342\,
            in2 => \N__33331\,
            in3 => \N__33315\,
            lcout => \b2v_inst20.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_4_c_RNO_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33291\,
            in1 => \N__33279\,
            in2 => \N__33268\,
            in3 => \N__33252\,
            lcout => \b2v_inst20.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_5_c_RNO_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33225\,
            in1 => \N__33213\,
            in2 => \N__33202\,
            in3 => \N__33186\,
            lcout => \b2v_inst20.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_6_c_RNO_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33159\,
            in1 => \N__33148\,
            in2 => \N__33133\,
            in3 => \N__33115\,
            lcout => \b2v_inst20.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNIQ7EG4_1_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33514\,
            in1 => \N__33532\,
            in2 => \_gnd_net_\,
            in3 => \N__34069\,
            lcout => \b2v_inst200.curr_stateZ0Z_1\,
            ltout => \b2v_inst200.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33085\,
            in3 => \N__33821\,
            lcout => \N_405\,
            ltout => \N_405_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__33622\,
            in1 => \N__33616\,
            in2 => \N__33547\,
            in3 => \N__33522\,
            lcout => \b2v_inst200.m6_i_0\,
            ltout => \b2v_inst200.m6_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m6_i_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110001"
        )
    port map (
            in0 => \N__33768\,
            in1 => \N__33802\,
            in2 => \N__33544\,
            in3 => \N__33822\,
            lcout => OPEN,
            ltout => \b2v_inst200.N_57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNIKHBJ4_0_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33724\,
            in2 => \N__33541\,
            in3 => \N__34070\,
            lcout => \b2v_inst200.curr_stateZ0Z_0\,
            ltout => \b2v_inst200.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m8_i_a2_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33803\,
            in2 => \N__33538\,
            in3 => \_gnd_net_\,
            lcout => \N_406\,
            ltout => \N_406_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m8_i_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__33805\,
            in1 => \N__34147\,
            in2 => \N__33535\,
            in3 => \N__33767\,
            lcout => \b2v_inst200.N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_1_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__33769\,
            in1 => \N__33804\,
            in2 => \N__33526\,
            in3 => \N__34146\,
            lcout => \b2v_inst200.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34667\,
            ce => \N__33683\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNI_0_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33806\,
            in2 => \_gnd_net_\,
            in3 => \N__33830\,
            lcout => \b2v_inst200.N_202\,
            ltout => \b2v_inst200.N_202_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.HDA_SDO_FPGA_RNIJCSM_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001001110"
        )
    port map (
            in0 => \N__34072\,
            in1 => \N__33838\,
            in2 => \N__33508\,
            in3 => \N__33850\,
            lcout => \HDA_SDO_FPGA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_7_c_RNO_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33483\,
            in1 => \N__33471\,
            in2 => \N__33460\,
            in3 => \N__33444\,
            lcout => \b2v_inst20.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m11_0_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111101"
        )
    port map (
            in0 => \N__33770\,
            in1 => \N__34145\,
            in2 => \N__34123\,
            in3 => \N__33849\,
            lcout => \G_2788\,
            ltout => \G_2788_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNI52VB_2_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__34105\,
            in1 => \_gnd_net_\,
            in2 => \N__34096\,
            in3 => \N__34071\,
            lcout => \b2v_inst200.curr_stateZ0Z_2\,
            ltout => \b2v_inst200.curr_stateZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.HDA_SDO_FPGA_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011111000"
        )
    port map (
            in0 => \N__33831\,
            in1 => \N__33808\,
            in2 => \N__33841\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.HDA_SDO_FPGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34673\,
            ce => \N__33681\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_0_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001001"
        )
    port map (
            in0 => \N__33832\,
            in1 => \N__33807\,
            in2 => \N__33777\,
            in3 => \N__33730\,
            lcout => \b2v_inst200.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34673\,
            ce => \N__33681\,
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_6_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34264\,
            lcout => \b2v_inst6.count_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34680\,
            ce => \N__34417\,
            sr => \N__35295\
        );

    \b2v_inst6.count_RNIRDTD4_2_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34276\,
            in1 => \N__34284\,
            in2 => \_gnd_net_\,
            in3 => \N__34415\,
            lcout => \b2v_inst6.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIVVMK_1_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__34216\,
            in1 => \N__35020\,
            in2 => \_gnd_net_\,
            in3 => \N__35271\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI3A4A4_1_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34291\,
            in2 => \N__33625\,
            in3 => \N__34414\,
            lcout => \b2v_inst6.countZ0Z_1\,
            ltout => \b2v_inst6.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_1_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35021\,
            in2 => \N__34294\,
            in3 => \N__35272\,
            lcout => \b2v_inst6.count_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34680\,
            ce => \N__34417\,
            sr => \N__35295\
        );

    \b2v_inst6.count_2_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34285\,
            lcout => \b2v_inst6.count_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34680\,
            ce => \N__34417\,
            sr => \N__35295\
        );

    \b2v_inst6.count_RNI3Q1E4_6_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34416\,
            in1 => \N__34270\,
            in2 => \_gnd_net_\,
            in3 => \N__34263\,
            lcout => \b2v_inst6.countZ0Z_6\,
            ltout => \b2v_inst6.countZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI_1_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34249\,
            in1 => \N__34231\,
            in2 => \N__34219\,
            in3 => \N__34215\,
            lcout => \b2v_inst6.un12_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI_15_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34174\,
            in1 => \N__34201\,
            in2 => \N__34804\,
            in3 => \N__34849\,
            lcout => \b2v_inst6.un12_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNITOVM4_12_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34180\,
            in1 => \N__34188\,
            in2 => \_gnd_net_\,
            in3 => \N__34425\,
            lcout => \b2v_inst6.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_12_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34189\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.count_3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34685\,
            ce => \N__34435\,
            sr => \N__35308\
        );

    \b2v_inst6.count_RNIVR0N4_13_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34153\,
            in1 => \N__34426\,
            in2 => \_gnd_net_\,
            in3 => \N__34161\,
            lcout => \b2v_inst6.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_13_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34162\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.count_3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34685\,
            ce => \N__34435\,
            sr => \N__35308\
        );

    \b2v_inst6.count_RNI1V1N4_14_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34828\,
            in1 => \N__34836\,
            in2 => \_gnd_net_\,
            in3 => \N__34427\,
            lcout => \b2v_inst6.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_14_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.count_3_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34685\,
            ce => \N__34435\,
            sr => \N__35308\
        );

    \b2v_inst6.count_RNI323N4_15_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34822\,
            in1 => \N__34815\,
            in2 => \_gnd_net_\,
            in3 => \N__34428\,
            lcout => \b2v_inst6.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un8_rsmrst_pwrgd_4_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34789\,
            in1 => \N__34783\,
            in2 => \N__34777\,
            in3 => \N__34768\,
            lcout => \SYNTHESIZED_WIRE_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIVVMK_0_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__35025\,
            in1 => \N__34915\,
            in2 => \_gnd_net_\,
            in3 => \N__35222\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI294A4_0_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34723\,
            in2 => \N__34729\,
            in3 => \N__34368\,
            lcout => \b2v_inst6.countZ0Z_0\,
            ltout => \b2v_inst6.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_0_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34914\,
            in2 => \N__34726\,
            in3 => \N__35224\,
            lcout => \b2v_inst6.count_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34688\,
            ce => \N__34421\,
            sr => \N__35228\
        );

    \b2v_inst6.count_3_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__35223\,
            in1 => \N__34916\,
            in2 => \N__35094\,
            in3 => \N__34717\,
            lcout => \b2v_inst6.count_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34688\,
            ce => \N__34421\,
            sr => \N__35228\
        );

    \b2v_inst6.count_RNI_3_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__35125\,
            in1 => \N__35092\,
            in2 => \N__35062\,
            in3 => \N__35016\,
            lcout => OPEN,
            ltout => \b2v_inst6.un12_clk_100khz_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI_0_1_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34987\,
            in1 => \N__34981\,
            in2 => \N__34972\,
            in3 => \N__34969\,
            lcout => \b2v_inst6.N_1_i\,
            ltout => \b2v_inst6.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI_1_1_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34945\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.N_1_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
