// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Aug 28 2022 11:53:55

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VR_READY_VCCINAUX,
    V33A_ENn,
    V1P8A_EN,
    VDDQ_EN,
    VCCST_OVERRIDE_3V3,
    V5S_OK,
    SLP_S3n,
    SLP_S0n,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    GPIO_FPGA_SoC_2,
    VCCIN_VR_PROCHOT_FPGA,
    SLP_SUSn,
    CPU_C10_GATE_N,
    VCCST_EN,
    V33DSW_OK,
    TPM_GPIO,
    SUSWARN_N,
    PLTRSTn,
    GPIO_FPGA_SoC_4,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    FPGA_OSC,
    VCCST_PWRGD,
    SYS_PWROK,
    SPI_FP_IO2,
    SATAXPCIE1_FPGA,
    GPIO_FPGA_EXP_1,
    VCCINAUX_VR_PROCHOT_FPGA,
    VCCINAUX_VR_PE,
    HDA_SDO_ATP,
    GPIO_FPGA_EXP_2,
    VPP_EN,
    VDDQ_OK,
    SUSACK_N,
    SLP_S4n,
    VCCST_CPU_OK,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    GPIO_FPGA_SoC_1,
    DSW_PWROK,
    V5A_EN,
    GPIO_FPGA_SoC_3,
    VR_PROCHOT_FPGA_OUT_N,
    VPP_OK,
    VCCIN_VR_PE,
    VCCIN_EN,
    SOC_SPKR,
    SLP_S5n,
    V12_MAIN_MON,
    SPI_FP_IO3,
    SATAXPCIE0_FPGA,
    V33A_OK,
    PCH_PWROK,
    FPGA_SLP_WLAN_N);

    input VR_READY_VCCINAUX;
    output V33A_ENn;
    output V1P8A_EN;
    output VDDQ_EN;
    input VCCST_OVERRIDE_3V3;
    input V5S_OK;
    input SLP_S3n;
    input SLP_S0n;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input GPIO_FPGA_SoC_2;
    input VCCIN_VR_PROCHOT_FPGA;
    input SLP_SUSn;
    input CPU_C10_GATE_N;
    output VCCST_EN;
    input V33DSW_OK;
    input TPM_GPIO;
    output SUSWARN_N;
    input PLTRSTn;
    input GPIO_FPGA_SoC_4;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output SYS_PWROK;
    input SPI_FP_IO2;
    input SATAXPCIE1_FPGA;
    input GPIO_FPGA_EXP_1;
    input VCCINAUX_VR_PROCHOT_FPGA;
    output VCCINAUX_VR_PE;
    output HDA_SDO_ATP;
    input GPIO_FPGA_EXP_2;
    output VPP_EN;
    input VDDQ_OK;
    input SUSACK_N;
    input SLP_S4n;
    input VCCST_CPU_OK;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input GPIO_FPGA_SoC_1;
    output DSW_PWROK;
    output V5A_EN;
    input GPIO_FPGA_SoC_3;
    input VR_PROCHOT_FPGA_OUT_N;
    input VPP_OK;
    output VCCIN_VR_PE;
    output VCCIN_EN;
    input SOC_SPKR;
    input SLP_S5n;
    input V12_MAIN_MON;
    input SPI_FP_IO3;
    input SATAXPCIE0_FPGA;
    input V33A_OK;
    output PCH_PWROK;
    input FPGA_SLP_WLAN_N;

    wire N__21309;
    wire N__21308;
    wire N__21307;
    wire N__21300;
    wire N__21299;
    wire N__21298;
    wire N__21291;
    wire N__21290;
    wire N__21289;
    wire N__21282;
    wire N__21281;
    wire N__21280;
    wire N__21273;
    wire N__21272;
    wire N__21271;
    wire N__21264;
    wire N__21263;
    wire N__21262;
    wire N__21255;
    wire N__21254;
    wire N__21253;
    wire N__21246;
    wire N__21245;
    wire N__21244;
    wire N__21237;
    wire N__21236;
    wire N__21235;
    wire N__21228;
    wire N__21227;
    wire N__21226;
    wire N__21219;
    wire N__21218;
    wire N__21217;
    wire N__21210;
    wire N__21209;
    wire N__21208;
    wire N__21201;
    wire N__21200;
    wire N__21199;
    wire N__21192;
    wire N__21191;
    wire N__21190;
    wire N__21183;
    wire N__21182;
    wire N__21181;
    wire N__21174;
    wire N__21173;
    wire N__21172;
    wire N__21165;
    wire N__21164;
    wire N__21163;
    wire N__21156;
    wire N__21155;
    wire N__21154;
    wire N__21147;
    wire N__21146;
    wire N__21145;
    wire N__21138;
    wire N__21137;
    wire N__21136;
    wire N__21129;
    wire N__21128;
    wire N__21127;
    wire N__21120;
    wire N__21119;
    wire N__21118;
    wire N__21111;
    wire N__21110;
    wire N__21109;
    wire N__21102;
    wire N__21101;
    wire N__21100;
    wire N__21093;
    wire N__21092;
    wire N__21091;
    wire N__21084;
    wire N__21083;
    wire N__21082;
    wire N__21075;
    wire N__21074;
    wire N__21073;
    wire N__21066;
    wire N__21065;
    wire N__21064;
    wire N__21057;
    wire N__21056;
    wire N__21055;
    wire N__21048;
    wire N__21047;
    wire N__21046;
    wire N__21039;
    wire N__21038;
    wire N__21037;
    wire N__21030;
    wire N__21029;
    wire N__21028;
    wire N__21021;
    wire N__21020;
    wire N__21019;
    wire N__21012;
    wire N__21011;
    wire N__21010;
    wire N__21003;
    wire N__21002;
    wire N__21001;
    wire N__20994;
    wire N__20993;
    wire N__20992;
    wire N__20985;
    wire N__20984;
    wire N__20983;
    wire N__20976;
    wire N__20975;
    wire N__20974;
    wire N__20967;
    wire N__20966;
    wire N__20965;
    wire N__20958;
    wire N__20957;
    wire N__20956;
    wire N__20949;
    wire N__20948;
    wire N__20947;
    wire N__20940;
    wire N__20939;
    wire N__20938;
    wire N__20931;
    wire N__20930;
    wire N__20929;
    wire N__20922;
    wire N__20921;
    wire N__20920;
    wire N__20913;
    wire N__20912;
    wire N__20911;
    wire N__20904;
    wire N__20903;
    wire N__20902;
    wire N__20895;
    wire N__20894;
    wire N__20893;
    wire N__20886;
    wire N__20885;
    wire N__20884;
    wire N__20877;
    wire N__20876;
    wire N__20875;
    wire N__20868;
    wire N__20867;
    wire N__20866;
    wire N__20859;
    wire N__20858;
    wire N__20857;
    wire N__20850;
    wire N__20849;
    wire N__20848;
    wire N__20841;
    wire N__20840;
    wire N__20839;
    wire N__20832;
    wire N__20831;
    wire N__20830;
    wire N__20823;
    wire N__20822;
    wire N__20821;
    wire N__20814;
    wire N__20813;
    wire N__20812;
    wire N__20805;
    wire N__20804;
    wire N__20803;
    wire N__20796;
    wire N__20795;
    wire N__20794;
    wire N__20787;
    wire N__20786;
    wire N__20785;
    wire N__20768;
    wire N__20765;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20747;
    wire N__20746;
    wire N__20745;
    wire N__20744;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20729;
    wire N__20724;
    wire N__20717;
    wire N__20716;
    wire N__20715;
    wire N__20712;
    wire N__20709;
    wire N__20708;
    wire N__20705;
    wire N__20704;
    wire N__20703;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20663;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20651;
    wire N__20642;
    wire N__20641;
    wire N__20638;
    wire N__20637;
    wire N__20636;
    wire N__20635;
    wire N__20632;
    wire N__20631;
    wire N__20630;
    wire N__20629;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20615;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20605;
    wire N__20604;
    wire N__20601;
    wire N__20600;
    wire N__20597;
    wire N__20596;
    wire N__20595;
    wire N__20594;
    wire N__20593;
    wire N__20586;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20564;
    wire N__20561;
    wire N__20560;
    wire N__20559;
    wire N__20558;
    wire N__20557;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20547;
    wire N__20544;
    wire N__20543;
    wire N__20542;
    wire N__20539;
    wire N__20538;
    wire N__20535;
    wire N__20534;
    wire N__20533;
    wire N__20532;
    wire N__20529;
    wire N__20526;
    wire N__20521;
    wire N__20518;
    wire N__20511;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20499;
    wire N__20496;
    wire N__20495;
    wire N__20492;
    wire N__20491;
    wire N__20488;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20474;
    wire N__20473;
    wire N__20472;
    wire N__20471;
    wire N__20468;
    wire N__20467;
    wire N__20466;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20451;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20443;
    wire N__20438;
    wire N__20429;
    wire N__20428;
    wire N__20423;
    wire N__20418;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20408;
    wire N__20407;
    wire N__20404;
    wire N__20399;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20370;
    wire N__20365;
    wire N__20362;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20341;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20325;
    wire N__20320;
    wire N__20317;
    wire N__20314;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20296;
    wire N__20291;
    wire N__20288;
    wire N__20285;
    wire N__20282;
    wire N__20279;
    wire N__20274;
    wire N__20265;
    wire N__20260;
    wire N__20257;
    wire N__20254;
    wire N__20251;
    wire N__20248;
    wire N__20241;
    wire N__20238;
    wire N__20233;
    wire N__20228;
    wire N__20223;
    wire N__20216;
    wire N__20207;
    wire N__20206;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20192;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20159;
    wire N__20158;
    wire N__20157;
    wire N__20156;
    wire N__20155;
    wire N__20154;
    wire N__20153;
    wire N__20152;
    wire N__20151;
    wire N__20150;
    wire N__20149;
    wire N__20148;
    wire N__20147;
    wire N__20146;
    wire N__20145;
    wire N__20144;
    wire N__20143;
    wire N__20142;
    wire N__20141;
    wire N__20140;
    wire N__20139;
    wire N__20138;
    wire N__20137;
    wire N__20136;
    wire N__20135;
    wire N__20134;
    wire N__20133;
    wire N__20132;
    wire N__20131;
    wire N__20130;
    wire N__20129;
    wire N__20128;
    wire N__20127;
    wire N__20126;
    wire N__20125;
    wire N__20124;
    wire N__20123;
    wire N__20122;
    wire N__20121;
    wire N__20120;
    wire N__20119;
    wire N__20118;
    wire N__20117;
    wire N__20116;
    wire N__20115;
    wire N__20114;
    wire N__20113;
    wire N__20112;
    wire N__20111;
    wire N__20110;
    wire N__20109;
    wire N__20108;
    wire N__20107;
    wire N__20106;
    wire N__20105;
    wire N__20104;
    wire N__20103;
    wire N__20102;
    wire N__20101;
    wire N__20100;
    wire N__20099;
    wire N__20098;
    wire N__20097;
    wire N__20096;
    wire N__20095;
    wire N__20094;
    wire N__20093;
    wire N__20092;
    wire N__20091;
    wire N__20090;
    wire N__20089;
    wire N__20088;
    wire N__20087;
    wire N__20086;
    wire N__20085;
    wire N__20084;
    wire N__20083;
    wire N__20082;
    wire N__20081;
    wire N__20080;
    wire N__20079;
    wire N__20078;
    wire N__20077;
    wire N__20076;
    wire N__20075;
    wire N__20074;
    wire N__20073;
    wire N__20072;
    wire N__20071;
    wire N__20070;
    wire N__20069;
    wire N__20068;
    wire N__20067;
    wire N__20066;
    wire N__20065;
    wire N__20064;
    wire N__20063;
    wire N__20062;
    wire N__20061;
    wire N__20060;
    wire N__20059;
    wire N__20058;
    wire N__20057;
    wire N__20056;
    wire N__20047;
    wire N__20040;
    wire N__20033;
    wire N__20024;
    wire N__20015;
    wire N__20008;
    wire N__20001;
    wire N__19992;
    wire N__19983;
    wire N__19974;
    wire N__19969;
    wire N__19960;
    wire N__19951;
    wire N__19942;
    wire N__19935;
    wire N__19926;
    wire N__19919;
    wire N__19910;
    wire N__19901;
    wire N__19894;
    wire N__19885;
    wire N__19880;
    wire N__19871;
    wire N__19868;
    wire N__19859;
    wire N__19852;
    wire N__19843;
    wire N__19840;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19821;
    wire N__19816;
    wire N__19813;
    wire N__19812;
    wire N__19811;
    wire N__19810;
    wire N__19809;
    wire N__19808;
    wire N__19807;
    wire N__19806;
    wire N__19803;
    wire N__19802;
    wire N__19799;
    wire N__19798;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19787;
    wire N__19786;
    wire N__19785;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19774;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19763;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19742;
    wire N__19741;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19543;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19525;
    wire N__19524;
    wire N__19523;
    wire N__19520;
    wire N__19515;
    wire N__19512;
    wire N__19507;
    wire N__19504;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19471;
    wire N__19470;
    wire N__19467;
    wire N__19466;
    wire N__19465;
    wire N__19460;
    wire N__19453;
    wire N__19448;
    wire N__19445;
    wire N__19444;
    wire N__19443;
    wire N__19436;
    wire N__19435;
    wire N__19434;
    wire N__19433;
    wire N__19432;
    wire N__19431;
    wire N__19430;
    wire N__19427;
    wire N__19418;
    wire N__19413;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19388;
    wire N__19385;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19360;
    wire N__19357;
    wire N__19356;
    wire N__19353;
    wire N__19348;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19327;
    wire N__19326;
    wire N__19325;
    wire N__19324;
    wire N__19323;
    wire N__19310;
    wire N__19307;
    wire N__19306;
    wire N__19305;
    wire N__19304;
    wire N__19303;
    wire N__19302;
    wire N__19289;
    wire N__19286;
    wire N__19285;
    wire N__19284;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19237;
    wire N__19234;
    wire N__19229;
    wire N__19228;
    wire N__19227;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19196;
    wire N__19195;
    wire N__19190;
    wire N__19187;
    wire N__19186;
    wire N__19183;
    wire N__19180;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19085;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19070;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19058;
    wire N__19057;
    wire N__19054;
    wire N__19051;
    wire N__19046;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19034;
    wire N__19033;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19019;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19007;
    wire N__19006;
    wire N__19003;
    wire N__19000;
    wire N__18995;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18983;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18968;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18956;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18941;
    wire N__18940;
    wire N__18937;
    wire N__18934;
    wire N__18929;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18914;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18877;
    wire N__18874;
    wire N__18871;
    wire N__18868;
    wire N__18865;
    wire N__18860;
    wire N__18859;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18845;
    wire N__18844;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18830;
    wire N__18827;
    wire N__18826;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18812;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18797;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18782;
    wire N__18781;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18767;
    wire N__18766;
    wire N__18763;
    wire N__18760;
    wire N__18757;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18736;
    wire N__18731;
    wire N__18728;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18713;
    wire N__18710;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18674;
    wire N__18671;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18635;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18623;
    wire N__18622;
    wire N__18619;
    wire N__18616;
    wire N__18611;
    wire N__18608;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18589;
    wire N__18586;
    wire N__18583;
    wire N__18578;
    wire N__18577;
    wire N__18574;
    wire N__18571;
    wire N__18566;
    wire N__18565;
    wire N__18562;
    wire N__18559;
    wire N__18556;
    wire N__18551;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18529;
    wire N__18526;
    wire N__18523;
    wire N__18522;
    wire N__18519;
    wire N__18516;
    wire N__18513;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18490;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18458;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18446;
    wire N__18443;
    wire N__18442;
    wire N__18439;
    wire N__18436;
    wire N__18431;
    wire N__18428;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18413;
    wire N__18410;
    wire N__18409;
    wire N__18406;
    wire N__18403;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18388;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18377;
    wire N__18376;
    wire N__18375;
    wire N__18374;
    wire N__18371;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18357;
    wire N__18356;
    wire N__18353;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18337;
    wire N__18336;
    wire N__18333;
    wire N__18328;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18318;
    wire N__18315;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18301;
    wire N__18294;
    wire N__18289;
    wire N__18284;
    wire N__18281;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18266;
    wire N__18263;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18250;
    wire N__18247;
    wire N__18244;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18234;
    wire N__18233;
    wire N__18226;
    wire N__18223;
    wire N__18218;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18206;
    wire N__18205;
    wire N__18202;
    wire N__18199;
    wire N__18194;
    wire N__18193;
    wire N__18190;
    wire N__18187;
    wire N__18184;
    wire N__18179;
    wire N__18178;
    wire N__18175;
    wire N__18172;
    wire N__18167;
    wire N__18166;
    wire N__18163;
    wire N__18160;
    wire N__18155;
    wire N__18154;
    wire N__18151;
    wire N__18148;
    wire N__18143;
    wire N__18142;
    wire N__18139;
    wire N__18136;
    wire N__18133;
    wire N__18128;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18116;
    wire N__18115;
    wire N__18114;
    wire N__18111;
    wire N__18106;
    wire N__18101;
    wire N__18098;
    wire N__18097;
    wire N__18096;
    wire N__18093;
    wire N__18088;
    wire N__18083;
    wire N__18080;
    wire N__18079;
    wire N__18078;
    wire N__18077;
    wire N__18074;
    wire N__18069;
    wire N__18066;
    wire N__18059;
    wire N__18056;
    wire N__18055;
    wire N__18052;
    wire N__18051;
    wire N__18048;
    wire N__18045;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18023;
    wire N__18020;
    wire N__18019;
    wire N__18018;
    wire N__18017;
    wire N__18016;
    wire N__18013;
    wire N__18008;
    wire N__18007;
    wire N__18006;
    wire N__18001;
    wire N__18000;
    wire N__17997;
    wire N__17994;
    wire N__17991;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17973;
    wire N__17968;
    wire N__17965;
    wire N__17954;
    wire N__17951;
    wire N__17950;
    wire N__17949;
    wire N__17946;
    wire N__17941;
    wire N__17936;
    wire N__17933;
    wire N__17932;
    wire N__17931;
    wire N__17930;
    wire N__17927;
    wire N__17920;
    wire N__17915;
    wire N__17912;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17890;
    wire N__17887;
    wire N__17884;
    wire N__17883;
    wire N__17880;
    wire N__17877;
    wire N__17874;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17849;
    wire N__17848;
    wire N__17845;
    wire N__17842;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17832;
    wire N__17829;
    wire N__17824;
    wire N__17819;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17777;
    wire N__17776;
    wire N__17773;
    wire N__17770;
    wire N__17767;
    wire N__17764;
    wire N__17761;
    wire N__17758;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17746;
    wire N__17741;
    wire N__17738;
    wire N__17737;
    wire N__17734;
    wire N__17731;
    wire N__17728;
    wire N__17725;
    wire N__17722;
    wire N__17719;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17702;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17692;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17669;
    wire N__17668;
    wire N__17667;
    wire N__17666;
    wire N__17663;
    wire N__17656;
    wire N__17651;
    wire N__17648;
    wire N__17647;
    wire N__17644;
    wire N__17643;
    wire N__17640;
    wire N__17637;
    wire N__17634;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17611;
    wire N__17608;
    wire N__17607;
    wire N__17604;
    wire N__17601;
    wire N__17596;
    wire N__17591;
    wire N__17590;
    wire N__17587;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17577;
    wire N__17576;
    wire N__17571;
    wire N__17566;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17545;
    wire N__17544;
    wire N__17541;
    wire N__17536;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17521;
    wire N__17518;
    wire N__17515;
    wire N__17514;
    wire N__17511;
    wire N__17506;
    wire N__17501;
    wire N__17500;
    wire N__17497;
    wire N__17494;
    wire N__17489;
    wire N__17488;
    wire N__17485;
    wire N__17482;
    wire N__17477;
    wire N__17476;
    wire N__17473;
    wire N__17470;
    wire N__17467;
    wire N__17462;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17450;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17438;
    wire N__17437;
    wire N__17434;
    wire N__17431;
    wire N__17426;
    wire N__17425;
    wire N__17422;
    wire N__17419;
    wire N__17416;
    wire N__17411;
    wire N__17410;
    wire N__17407;
    wire N__17404;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17372;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17360;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17345;
    wire N__17344;
    wire N__17341;
    wire N__17338;
    wire N__17333;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17309;
    wire N__17308;
    wire N__17305;
    wire N__17302;
    wire N__17297;
    wire N__17296;
    wire N__17293;
    wire N__17290;
    wire N__17287;
    wire N__17282;
    wire N__17281;
    wire N__17278;
    wire N__17275;
    wire N__17270;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17258;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17246;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17236;
    wire N__17231;
    wire N__17230;
    wire N__17227;
    wire N__17224;
    wire N__17219;
    wire N__17218;
    wire N__17215;
    wire N__17212;
    wire N__17207;
    wire N__17206;
    wire N__17203;
    wire N__17200;
    wire N__17195;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17185;
    wire N__17180;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17165;
    wire N__17164;
    wire N__17161;
    wire N__17158;
    wire N__17153;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17141;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17126;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17096;
    wire N__17093;
    wire N__17090;
    wire N__17087;
    wire N__17084;
    wire N__17081;
    wire N__17078;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17063;
    wire N__17060;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17050;
    wire N__17049;
    wire N__17046;
    wire N__17041;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17026;
    wire N__17023;
    wire N__17022;
    wire N__17019;
    wire N__17014;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16999;
    wire N__16996;
    wire N__16993;
    wire N__16990;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16931;
    wire N__16930;
    wire N__16927;
    wire N__16924;
    wire N__16923;
    wire N__16918;
    wire N__16915;
    wire N__16910;
    wire N__16909;
    wire N__16908;
    wire N__16905;
    wire N__16900;
    wire N__16895;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16885;
    wire N__16882;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16826;
    wire N__16825;
    wire N__16822;
    wire N__16819;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16774;
    wire N__16773;
    wire N__16772;
    wire N__16771;
    wire N__16770;
    wire N__16769;
    wire N__16762;
    wire N__16761;
    wire N__16760;
    wire N__16759;
    wire N__16758;
    wire N__16757;
    wire N__16756;
    wire N__16753;
    wire N__16746;
    wire N__16743;
    wire N__16740;
    wire N__16739;
    wire N__16738;
    wire N__16737;
    wire N__16736;
    wire N__16735;
    wire N__16732;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16712;
    wire N__16709;
    wire N__16700;
    wire N__16697;
    wire N__16692;
    wire N__16687;
    wire N__16676;
    wire N__16673;
    wire N__16672;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16660;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16645;
    wire N__16642;
    wire N__16639;
    wire N__16634;
    wire N__16631;
    wire N__16630;
    wire N__16629;
    wire N__16624;
    wire N__16623;
    wire N__16620;
    wire N__16617;
    wire N__16614;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16591;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16583;
    wire N__16582;
    wire N__16581;
    wire N__16578;
    wire N__16577;
    wire N__16574;
    wire N__16567;
    wire N__16564;
    wire N__16561;
    wire N__16558;
    wire N__16557;
    wire N__16556;
    wire N__16553;
    wire N__16546;
    wire N__16543;
    wire N__16538;
    wire N__16537;
    wire N__16534;
    wire N__16531;
    wire N__16528;
    wire N__16525;
    wire N__16522;
    wire N__16517;
    wire N__16510;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16489;
    wire N__16486;
    wire N__16483;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16469;
    wire N__16468;
    wire N__16467;
    wire N__16466;
    wire N__16465;
    wire N__16462;
    wire N__16461;
    wire N__16460;
    wire N__16459;
    wire N__16458;
    wire N__16453;
    wire N__16452;
    wire N__16449;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16439;
    wire N__16434;
    wire N__16431;
    wire N__16428;
    wire N__16425;
    wire N__16420;
    wire N__16403;
    wire N__16402;
    wire N__16399;
    wire N__16398;
    wire N__16397;
    wire N__16396;
    wire N__16395;
    wire N__16394;
    wire N__16393;
    wire N__16390;
    wire N__16389;
    wire N__16388;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16372;
    wire N__16367;
    wire N__16362;
    wire N__16359;
    wire N__16346;
    wire N__16345;
    wire N__16344;
    wire N__16343;
    wire N__16340;
    wire N__16339;
    wire N__16336;
    wire N__16335;
    wire N__16334;
    wire N__16331;
    wire N__16330;
    wire N__16329;
    wire N__16326;
    wire N__16323;
    wire N__16318;
    wire N__16315;
    wire N__16312;
    wire N__16305;
    wire N__16292;
    wire N__16289;
    wire N__16288;
    wire N__16287;
    wire N__16286;
    wire N__16285;
    wire N__16284;
    wire N__16283;
    wire N__16282;
    wire N__16281;
    wire N__16276;
    wire N__16273;
    wire N__16268;
    wire N__16265;
    wire N__16258;
    wire N__16255;
    wire N__16244;
    wire N__16243;
    wire N__16242;
    wire N__16239;
    wire N__16238;
    wire N__16237;
    wire N__16236;
    wire N__16235;
    wire N__16232;
    wire N__16231;
    wire N__16228;
    wire N__16225;
    wire N__16222;
    wire N__16219;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16187;
    wire N__16186;
    wire N__16185;
    wire N__16184;
    wire N__16181;
    wire N__16180;
    wire N__16177;
    wire N__16174;
    wire N__16173;
    wire N__16172;
    wire N__16169;
    wire N__16168;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16156;
    wire N__16149;
    wire N__16146;
    wire N__16143;
    wire N__16130;
    wire N__16129;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16118;
    wire N__16117;
    wire N__16116;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16098;
    wire N__16095;
    wire N__16082;
    wire N__16081;
    wire N__16080;
    wire N__16077;
    wire N__16074;
    wire N__16073;
    wire N__16072;
    wire N__16069;
    wire N__16068;
    wire N__16067;
    wire N__16066;
    wire N__16065;
    wire N__16062;
    wire N__16059;
    wire N__16056;
    wire N__16053;
    wire N__16050;
    wire N__16043;
    wire N__16040;
    wire N__16035;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__16000;
    wire N__15999;
    wire N__15998;
    wire N__15997;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15981;
    wire N__15978;
    wire N__15975;
    wire N__15972;
    wire N__15969;
    wire N__15966;
    wire N__15963;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15944;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15916;
    wire N__15915;
    wire N__15914;
    wire N__15911;
    wire N__15908;
    wire N__15905;
    wire N__15904;
    wire N__15903;
    wire N__15902;
    wire N__15901;
    wire N__15900;
    wire N__15899;
    wire N__15896;
    wire N__15891;
    wire N__15886;
    wire N__15883;
    wire N__15880;
    wire N__15879;
    wire N__15876;
    wire N__15873;
    wire N__15872;
    wire N__15869;
    wire N__15868;
    wire N__15867;
    wire N__15864;
    wire N__15855;
    wire N__15852;
    wire N__15849;
    wire N__15846;
    wire N__15839;
    wire N__15836;
    wire N__15829;
    wire N__15818;
    wire N__15815;
    wire N__15814;
    wire N__15813;
    wire N__15812;
    wire N__15811;
    wire N__15810;
    wire N__15809;
    wire N__15808;
    wire N__15807;
    wire N__15804;
    wire N__15795;
    wire N__15792;
    wire N__15789;
    wire N__15788;
    wire N__15787;
    wire N__15782;
    wire N__15779;
    wire N__15778;
    wire N__15777;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15753;
    wire N__15750;
    wire N__15737;
    wire N__15736;
    wire N__15735;
    wire N__15734;
    wire N__15729;
    wire N__15726;
    wire N__15725;
    wire N__15724;
    wire N__15723;
    wire N__15722;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15712;
    wire N__15703;
    wire N__15700;
    wire N__15693;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15679;
    wire N__15676;
    wire N__15673;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15653;
    wire N__15652;
    wire N__15651;
    wire N__15650;
    wire N__15649;
    wire N__15648;
    wire N__15647;
    wire N__15646;
    wire N__15645;
    wire N__15644;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15636;
    wire N__15635;
    wire N__15632;
    wire N__15625;
    wire N__15622;
    wire N__15617;
    wire N__15612;
    wire N__15607;
    wire N__15602;
    wire N__15597;
    wire N__15584;
    wire N__15583;
    wire N__15582;
    wire N__15581;
    wire N__15576;
    wire N__15571;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15553;
    wire N__15550;
    wire N__15547;
    wire N__15542;
    wire N__15541;
    wire N__15540;
    wire N__15539;
    wire N__15538;
    wire N__15537;
    wire N__15532;
    wire N__15529;
    wire N__15526;
    wire N__15521;
    wire N__15512;
    wire N__15511;
    wire N__15510;
    wire N__15509;
    wire N__15508;
    wire N__15507;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15491;
    wire N__15482;
    wire N__15479;
    wire N__15476;
    wire N__15475;
    wire N__15472;
    wire N__15469;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15438;
    wire N__15435;
    wire N__15432;
    wire N__15429;
    wire N__15422;
    wire N__15419;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15407;
    wire N__15404;
    wire N__15401;
    wire N__15398;
    wire N__15395;
    wire N__15392;
    wire N__15389;
    wire N__15388;
    wire N__15385;
    wire N__15382;
    wire N__15377;
    wire N__15374;
    wire N__15373;
    wire N__15372;
    wire N__15369;
    wire N__15364;
    wire N__15359;
    wire N__15358;
    wire N__15357;
    wire N__15356;
    wire N__15355;
    wire N__15352;
    wire N__15351;
    wire N__15350;
    wire N__15347;
    wire N__15340;
    wire N__15337;
    wire N__15334;
    wire N__15331;
    wire N__15326;
    wire N__15323;
    wire N__15318;
    wire N__15315;
    wire N__15310;
    wire N__15307;
    wire N__15302;
    wire N__15301;
    wire N__15300;
    wire N__15299;
    wire N__15298;
    wire N__15295;
    wire N__15294;
    wire N__15293;
    wire N__15290;
    wire N__15289;
    wire N__15286;
    wire N__15283;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15259;
    wire N__15258;
    wire N__15255;
    wire N__15252;
    wire N__15241;
    wire N__15238;
    wire N__15235;
    wire N__15224;
    wire N__15223;
    wire N__15222;
    wire N__15221;
    wire N__15220;
    wire N__15217;
    wire N__15216;
    wire N__15213;
    wire N__15212;
    wire N__15211;
    wire N__15210;
    wire N__15209;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15190;
    wire N__15185;
    wire N__15180;
    wire N__15171;
    wire N__15164;
    wire N__15163;
    wire N__15162;
    wire N__15161;
    wire N__15158;
    wire N__15157;
    wire N__15152;
    wire N__15149;
    wire N__15148;
    wire N__15147;
    wire N__15144;
    wire N__15141;
    wire N__15138;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15128;
    wire N__15123;
    wire N__15120;
    wire N__15117;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15097;
    wire N__15094;
    wire N__15093;
    wire N__15092;
    wire N__15091;
    wire N__15090;
    wire N__15087;
    wire N__15086;
    wire N__15085;
    wire N__15084;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15070;
    wire N__15065;
    wire N__15058;
    wire N__15057;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15031;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15019;
    wire N__15016;
    wire N__15013;
    wire N__15012;
    wire N__15011;
    wire N__15010;
    wire N__15007;
    wire N__15004;
    wire N__15003;
    wire N__15002;
    wire N__14999;
    wire N__14994;
    wire N__14991;
    wire N__14988;
    wire N__14983;
    wire N__14978;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14960;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14939;
    wire N__14936;
    wire N__14933;
    wire N__14930;
    wire N__14927;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14902;
    wire N__14901;
    wire N__14898;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14854;
    wire N__14853;
    wire N__14852;
    wire N__14851;
    wire N__14850;
    wire N__14849;
    wire N__14848;
    wire N__14845;
    wire N__14844;
    wire N__14841;
    wire N__14840;
    wire N__14837;
    wire N__14836;
    wire N__14833;
    wire N__14832;
    wire N__14829;
    wire N__14828;
    wire N__14825;
    wire N__14824;
    wire N__14821;
    wire N__14820;
    wire N__14805;
    wire N__14804;
    wire N__14787;
    wire N__14784;
    wire N__14781;
    wire N__14778;
    wire N__14775;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14752;
    wire N__14751;
    wire N__14748;
    wire N__14745;
    wire N__14742;
    wire N__14741;
    wire N__14740;
    wire N__14737;
    wire N__14736;
    wire N__14733;
    wire N__14730;
    wire N__14727;
    wire N__14726;
    wire N__14723;
    wire N__14722;
    wire N__14719;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14707;
    wire N__14704;
    wire N__14701;
    wire N__14698;
    wire N__14693;
    wire N__14688;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14665;
    wire N__14662;
    wire N__14659;
    wire N__14658;
    wire N__14655;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14647;
    wire N__14646;
    wire N__14645;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14633;
    wire N__14630;
    wire N__14625;
    wire N__14622;
    wire N__14609;
    wire N__14606;
    wire N__14605;
    wire N__14604;
    wire N__14603;
    wire N__14602;
    wire N__14601;
    wire N__14598;
    wire N__14593;
    wire N__14590;
    wire N__14587;
    wire N__14586;
    wire N__14585;
    wire N__14582;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14570;
    wire N__14565;
    wire N__14560;
    wire N__14557;
    wire N__14546;
    wire N__14543;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14532;
    wire N__14531;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14523;
    wire N__14520;
    wire N__14517;
    wire N__14514;
    wire N__14511;
    wire N__14508;
    wire N__14505;
    wire N__14500;
    wire N__14497;
    wire N__14486;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14476;
    wire N__14473;
    wire N__14470;
    wire N__14467;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14455;
    wire N__14454;
    wire N__14451;
    wire N__14446;
    wire N__14445;
    wire N__14444;
    wire N__14443;
    wire N__14442;
    wire N__14437;
    wire N__14434;
    wire N__14427;
    wire N__14424;
    wire N__14417;
    wire N__14416;
    wire N__14411;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14398;
    wire N__14397;
    wire N__14396;
    wire N__14395;
    wire N__14394;
    wire N__14393;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14385;
    wire N__14382;
    wire N__14379;
    wire N__14374;
    wire N__14373;
    wire N__14370;
    wire N__14365;
    wire N__14362;
    wire N__14357;
    wire N__14354;
    wire N__14351;
    wire N__14348;
    wire N__14343;
    wire N__14338;
    wire N__14327;
    wire N__14324;
    wire N__14321;
    wire N__14318;
    wire N__14315;
    wire N__14312;
    wire N__14309;
    wire N__14306;
    wire N__14305;
    wire N__14304;
    wire N__14301;
    wire N__14296;
    wire N__14293;
    wire N__14290;
    wire N__14285;
    wire N__14282;
    wire N__14279;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14261;
    wire N__14258;
    wire N__14255;
    wire N__14252;
    wire N__14249;
    wire N__14246;
    wire N__14243;
    wire N__14240;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14197;
    wire N__14196;
    wire N__14195;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14182;
    wire N__14179;
    wire N__14178;
    wire N__14177;
    wire N__14174;
    wire N__14169;
    wire N__14166;
    wire N__14163;
    wire N__14160;
    wire N__14157;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14128;
    wire N__14127;
    wire N__14124;
    wire N__14123;
    wire N__14120;
    wire N__14119;
    wire N__14116;
    wire N__14113;
    wire N__14112;
    wire N__14111;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14088;
    wire N__14085;
    wire N__14082;
    wire N__14077;
    wire N__14072;
    wire N__14067;
    wire N__14062;
    wire N__14051;
    wire N__14048;
    wire N__14045;
    wire N__14042;
    wire N__14039;
    wire N__14036;
    wire N__14033;
    wire N__14030;
    wire N__14027;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14012;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14000;
    wire N__13997;
    wire N__13994;
    wire N__13993;
    wire N__13990;
    wire N__13987;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13964;
    wire N__13961;
    wire N__13958;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13937;
    wire N__13934;
    wire N__13931;
    wire N__13928;
    wire N__13927;
    wire N__13924;
    wire N__13921;
    wire N__13918;
    wire N__13913;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13901;
    wire N__13900;
    wire N__13897;
    wire N__13894;
    wire N__13889;
    wire N__13888;
    wire N__13885;
    wire N__13882;
    wire N__13879;
    wire N__13874;
    wire N__13873;
    wire N__13870;
    wire N__13867;
    wire N__13862;
    wire N__13859;
    wire N__13858;
    wire N__13855;
    wire N__13852;
    wire N__13847;
    wire N__13846;
    wire N__13843;
    wire N__13840;
    wire N__13837;
    wire N__13832;
    wire N__13831;
    wire N__13828;
    wire N__13825;
    wire N__13820;
    wire N__13817;
    wire N__13816;
    wire N__13813;
    wire N__13810;
    wire N__13805;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13793;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13781;
    wire N__13780;
    wire N__13777;
    wire N__13774;
    wire N__13771;
    wire N__13766;
    wire N__13765;
    wire N__13762;
    wire N__13759;
    wire N__13754;
    wire N__13753;
    wire N__13750;
    wire N__13747;
    wire N__13744;
    wire N__13739;
    wire N__13736;
    wire N__13733;
    wire N__13730;
    wire N__13727;
    wire N__13724;
    wire N__13721;
    wire N__13718;
    wire N__13715;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13702;
    wire N__13701;
    wire N__13700;
    wire N__13699;
    wire N__13698;
    wire N__13695;
    wire N__13690;
    wire N__13687;
    wire N__13684;
    wire N__13683;
    wire N__13680;
    wire N__13677;
    wire N__13674;
    wire N__13667;
    wire N__13658;
    wire N__13655;
    wire N__13654;
    wire N__13649;
    wire N__13646;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13631;
    wire N__13628;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13613;
    wire N__13610;
    wire N__13607;
    wire N__13606;
    wire N__13603;
    wire N__13600;
    wire N__13595;
    wire N__13594;
    wire N__13593;
    wire N__13590;
    wire N__13587;
    wire N__13586;
    wire N__13583;
    wire N__13576;
    wire N__13573;
    wire N__13570;
    wire N__13567;
    wire N__13564;
    wire N__13561;
    wire N__13556;
    wire N__13555;
    wire N__13550;
    wire N__13549;
    wire N__13548;
    wire N__13545;
    wire N__13540;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13528;
    wire N__13525;
    wire N__13522;
    wire N__13521;
    wire N__13518;
    wire N__13517;
    wire N__13514;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13456;
    wire N__13453;
    wire N__13450;
    wire N__13447;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13429;
    wire N__13426;
    wire N__13423;
    wire N__13422;
    wire N__13421;
    wire N__13418;
    wire N__13411;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13391;
    wire N__13388;
    wire N__13385;
    wire N__13382;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13367;
    wire N__13366;
    wire N__13363;
    wire N__13360;
    wire N__13355;
    wire N__13354;
    wire N__13351;
    wire N__13348;
    wire N__13345;
    wire N__13340;
    wire N__13339;
    wire N__13336;
    wire N__13333;
    wire N__13330;
    wire N__13325;
    wire N__13324;
    wire N__13321;
    wire N__13318;
    wire N__13313;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13274;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13246;
    wire N__13243;
    wire N__13240;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13222;
    wire N__13219;
    wire N__13218;
    wire N__13215;
    wire N__13212;
    wire N__13209;
    wire N__13202;
    wire N__13199;
    wire N__13198;
    wire N__13195;
    wire N__13192;
    wire N__13189;
    wire N__13184;
    wire N__13183;
    wire N__13180;
    wire N__13177;
    wire N__13174;
    wire N__13171;
    wire N__13168;
    wire N__13163;
    wire N__13160;
    wire N__13157;
    wire N__13156;
    wire N__13153;
    wire N__13150;
    wire N__13147;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13135;
    wire N__13132;
    wire N__13129;
    wire N__13126;
    wire N__13121;
    wire N__13118;
    wire N__13115;
    wire N__13114;
    wire N__13111;
    wire N__13108;
    wire N__13105;
    wire N__13100;
    wire N__13097;
    wire N__13096;
    wire N__13095;
    wire N__13092;
    wire N__13089;
    wire N__13088;
    wire N__13079;
    wire N__13076;
    wire N__13073;
    wire N__13070;
    wire N__13069;
    wire N__13068;
    wire N__13061;
    wire N__13058;
    wire N__13055;
    wire N__13052;
    wire N__13051;
    wire N__13046;
    wire N__13043;
    wire N__13042;
    wire N__13041;
    wire N__13038;
    wire N__13035;
    wire N__13032;
    wire N__13025;
    wire N__13022;
    wire N__13021;
    wire N__13018;
    wire N__13015;
    wire N__13012;
    wire N__13007;
    wire N__13006;
    wire N__13003;
    wire N__13000;
    wire N__12997;
    wire N__12992;
    wire N__12989;
    wire N__12986;
    wire N__12983;
    wire N__12980;
    wire N__12979;
    wire N__12976;
    wire N__12973;
    wire N__12968;
    wire N__12965;
    wire N__12962;
    wire N__12959;
    wire N__12956;
    wire N__12953;
    wire N__12950;
    wire N__12949;
    wire N__12946;
    wire N__12943;
    wire N__12940;
    wire N__12935;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12917;
    wire N__12916;
    wire N__12913;
    wire N__12910;
    wire N__12907;
    wire N__12904;
    wire N__12899;
    wire N__12896;
    wire N__12893;
    wire N__12890;
    wire N__12887;
    wire N__12884;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12874;
    wire N__12871;
    wire N__12868;
    wire N__12865;
    wire N__12862;
    wire N__12857;
    wire N__12854;
    wire N__12851;
    wire N__12848;
    wire N__12847;
    wire N__12844;
    wire N__12841;
    wire N__12838;
    wire N__12835;
    wire N__12832;
    wire N__12829;
    wire N__12826;
    wire N__12821;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12811;
    wire N__12808;
    wire N__12805;
    wire N__12802;
    wire N__12797;
    wire N__12794;
    wire N__12793;
    wire N__12790;
    wire N__12787;
    wire N__12784;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12764;
    wire N__12761;
    wire N__12758;
    wire N__12757;
    wire N__12754;
    wire N__12751;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12730;
    wire N__12727;
    wire N__12724;
    wire N__12721;
    wire N__12718;
    wire N__12715;
    wire N__12712;
    wire N__12707;
    wire N__12704;
    wire N__12701;
    wire N__12698;
    wire N__12697;
    wire N__12694;
    wire N__12691;
    wire N__12688;
    wire N__12683;
    wire N__12682;
    wire N__12679;
    wire N__12676;
    wire N__12671;
    wire N__12668;
    wire N__12665;
    wire N__12662;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12650;
    wire N__12647;
    wire N__12644;
    wire N__12641;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12626;
    wire N__12623;
    wire N__12622;
    wire N__12621;
    wire N__12620;
    wire N__12617;
    wire N__12614;
    wire N__12609;
    wire N__12606;
    wire N__12599;
    wire N__12596;
    wire N__12593;
    wire N__12592;
    wire N__12591;
    wire N__12590;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12575;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12557;
    wire N__12556;
    wire N__12553;
    wire N__12552;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12540;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12520;
    wire N__12519;
    wire N__12516;
    wire N__12515;
    wire N__12514;
    wire N__12511;
    wire N__12508;
    wire N__12505;
    wire N__12502;
    wire N__12499;
    wire N__12488;
    wire N__12485;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12472;
    wire N__12469;
    wire N__12468;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12456;
    wire N__12449;
    wire N__12446;
    wire N__12443;
    wire N__12442;
    wire N__12441;
    wire N__12440;
    wire N__12437;
    wire N__12434;
    wire N__12429;
    wire N__12426;
    wire N__12419;
    wire N__12416;
    wire N__12413;
    wire N__12412;
    wire N__12411;
    wire N__12410;
    wire N__12407;
    wire N__12404;
    wire N__12399;
    wire N__12396;
    wire N__12389;
    wire N__12386;
    wire N__12385;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12377;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12361;
    wire N__12356;
    wire N__12353;
    wire N__12352;
    wire N__12349;
    wire N__12348;
    wire N__12347;
    wire N__12344;
    wire N__12341;
    wire N__12336;
    wire N__12329;
    wire N__12326;
    wire N__12325;
    wire N__12322;
    wire N__12321;
    wire N__12320;
    wire N__12317;
    wire N__12314;
    wire N__12311;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12293;
    wire N__12290;
    wire N__12287;
    wire N__12286;
    wire N__12283;
    wire N__12282;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12270;
    wire N__12263;
    wire N__12260;
    wire N__12257;
    wire N__12256;
    wire N__12255;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12230;
    wire N__12227;
    wire N__12224;
    wire N__12223;
    wire N__12222;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12197;
    wire N__12194;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12179;
    wire N__12178;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12164;
    wire N__12163;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12149;
    wire N__12148;
    wire N__12145;
    wire N__12142;
    wire N__12139;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12122;
    wire N__12119;
    wire N__12118;
    wire N__12117;
    wire N__12116;
    wire N__12115;
    wire N__12114;
    wire N__12113;
    wire N__12112;
    wire N__12111;
    wire N__12110;
    wire N__12109;
    wire N__12108;
    wire N__12105;
    wire N__12098;
    wire N__12089;
    wire N__12080;
    wire N__12075;
    wire N__12068;
    wire N__12065;
    wire N__12064;
    wire N__12063;
    wire N__12062;
    wire N__12059;
    wire N__12052;
    wire N__12049;
    wire N__12046;
    wire N__12041;
    wire N__12040;
    wire N__12039;
    wire N__12038;
    wire N__12035;
    wire N__12030;
    wire N__12027;
    wire N__12024;
    wire N__12017;
    wire N__12016;
    wire N__12015;
    wire N__12012;
    wire N__12009;
    wire N__12006;
    wire N__12003;
    wire N__12000;
    wire N__11995;
    wire N__11990;
    wire N__11987;
    wire N__11986;
    wire N__11983;
    wire N__11982;
    wire N__11981;
    wire N__11978;
    wire N__11975;
    wire N__11970;
    wire N__11963;
    wire N__11960;
    wire N__11957;
    wire N__11956;
    wire N__11953;
    wire N__11952;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11940;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11909;
    wire N__11908;
    wire N__11905;
    wire N__11902;
    wire N__11897;
    wire N__11896;
    wire N__11893;
    wire N__11890;
    wire N__11885;
    wire N__11884;
    wire N__11881;
    wire N__11878;
    wire N__11875;
    wire N__11870;
    wire N__11869;
    wire N__11866;
    wire N__11863;
    wire N__11860;
    wire N__11855;
    wire N__11854;
    wire N__11851;
    wire N__11848;
    wire N__11843;
    wire N__11842;
    wire N__11839;
    wire N__11836;
    wire N__11833;
    wire N__11828;
    wire N__11827;
    wire N__11824;
    wire N__11821;
    wire N__11818;
    wire N__11813;
    wire N__11812;
    wire N__11809;
    wire N__11806;
    wire N__11801;
    wire N__11798;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11786;
    wire N__11783;
    wire N__11780;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11750;
    wire N__11747;
    wire N__11744;
    wire N__11743;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11714;
    wire N__11711;
    wire N__11708;
    wire N__11705;
    wire N__11702;
    wire N__11701;
    wire N__11698;
    wire N__11695;
    wire N__11690;
    wire N__11689;
    wire N__11684;
    wire N__11681;
    wire N__11678;
    wire N__11675;
    wire N__11672;
    wire N__11669;
    wire N__11666;
    wire N__11663;
    wire N__11660;
    wire N__11657;
    wire N__11654;
    wire N__11651;
    wire N__11648;
    wire N__11645;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11602;
    wire N__11601;
    wire N__11600;
    wire N__11597;
    wire N__11594;
    wire N__11591;
    wire N__11588;
    wire N__11585;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11560;
    wire N__11557;
    wire N__11552;
    wire N__11549;
    wire N__11546;
    wire N__11543;
    wire N__11540;
    wire N__11537;
    wire N__11534;
    wire N__11531;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11512;
    wire N__11509;
    wire N__11506;
    wire N__11501;
    wire N__11500;
    wire N__11499;
    wire N__11496;
    wire N__11495;
    wire N__11488;
    wire N__11485;
    wire N__11480;
    wire N__11477;
    wire N__11474;
    wire N__11471;
    wire N__11468;
    wire N__11465;
    wire N__11464;
    wire N__11461;
    wire N__11460;
    wire N__11457;
    wire N__11454;
    wire N__11449;
    wire N__11448;
    wire N__11447;
    wire N__11442;
    wire N__11439;
    wire N__11436;
    wire N__11429;
    wire N__11428;
    wire N__11425;
    wire N__11424;
    wire N__11421;
    wire N__11414;
    wire N__11411;
    wire N__11408;
    wire N__11405;
    wire N__11402;
    wire N__11399;
    wire N__11396;
    wire N__11393;
    wire N__11390;
    wire N__11387;
    wire N__11384;
    wire N__11381;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11356;
    wire N__11353;
    wire N__11350;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11332;
    wire N__11331;
    wire N__11330;
    wire N__11327;
    wire N__11326;
    wire N__11325;
    wire N__11320;
    wire N__11315;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11297;
    wire N__11294;
    wire N__11291;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11270;
    wire N__11267;
    wire N__11264;
    wire N__11261;
    wire N__11258;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11243;
    wire N__11240;
    wire N__11237;
    wire N__11234;
    wire N__11231;
    wire N__11228;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11180;
    wire N__11177;
    wire N__11176;
    wire N__11173;
    wire N__11172;
    wire N__11169;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11029;
    wire N__11026;
    wire N__11025;
    wire N__11022;
    wire N__11021;
    wire N__11018;
    wire N__11015;
    wire N__11012;
    wire N__11009;
    wire N__11006;
    wire N__11003;
    wire N__10998;
    wire N__10995;
    wire N__10990;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10907;
    wire N__10904;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10627;
    wire N__10626;
    wire N__10623;
    wire N__10622;
    wire N__10619;
    wire N__10614;
    wire N__10611;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10579;
    wire N__10576;
    wire N__10575;
    wire N__10572;
    wire N__10565;
    wire N__10562;
    wire N__10559;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10544;
    wire N__10543;
    wire N__10542;
    wire N__10539;
    wire N__10538;
    wire N__10535;
    wire N__10530;
    wire N__10527;
    wire N__10520;
    wire N__10517;
    wire N__10516;
    wire N__10513;
    wire N__10512;
    wire N__10509;
    wire N__10502;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10471;
    wire N__10468;
    wire N__10465;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10396;
    wire N__10393;
    wire N__10392;
    wire N__10389;
    wire N__10382;
    wire N__10379;
    wire N__10378;
    wire N__10377;
    wire N__10374;
    wire N__10373;
    wire N__10370;
    wire N__10365;
    wire N__10362;
    wire N__10355;
    wire N__10354;
    wire N__10353;
    wire N__10350;
    wire N__10349;
    wire N__10346;
    wire N__10341;
    wire N__10338;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10321;
    wire N__10318;
    wire N__10317;
    wire N__10314;
    wire N__10313;
    wire N__10310;
    wire N__10305;
    wire N__10302;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10238;
    wire N__10235;
    wire N__10234;
    wire N__10233;
    wire N__10230;
    wire N__10229;
    wire N__10226;
    wire N__10221;
    wire N__10218;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10186;
    wire N__10183;
    wire N__10182;
    wire N__10179;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10147;
    wire N__10144;
    wire N__10143;
    wire N__10140;
    wire N__10133;
    wire N__10130;
    wire N__10129;
    wire N__10126;
    wire N__10125;
    wire N__10122;
    wire N__10121;
    wire N__10118;
    wire N__10113;
    wire N__10110;
    wire N__10103;
    wire N__10102;
    wire N__10099;
    wire N__10098;
    wire N__10095;
    wire N__10094;
    wire N__10091;
    wire N__10086;
    wire N__10083;
    wire N__10076;
    wire N__10075;
    wire N__10074;
    wire N__10071;
    wire N__10070;
    wire N__10069;
    wire N__10066;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10046;
    wire N__10045;
    wire N__10042;
    wire N__10041;
    wire N__10038;
    wire N__10037;
    wire N__10034;
    wire N__10029;
    wire N__10026;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10012;
    wire N__10011;
    wire N__10008;
    wire N__10007;
    wire N__10004;
    wire N__9999;
    wire N__9996;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9973;
    wire N__9970;
    wire N__9969;
    wire N__9966;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9889;
    wire N__9886;
    wire N__9885;
    wire N__9882;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9863;
    wire N__9860;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9818;
    wire N__9815;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9796;
    wire N__9793;
    wire N__9790;
    wire N__9787;
    wire N__9782;
    wire N__9779;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9769;
    wire N__9768;
    wire N__9765;
    wire N__9762;
    wire N__9759;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9709;
    wire N__9706;
    wire N__9703;
    wire N__9698;
    wire N__9695;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9683;
    wire N__9680;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9670;
    wire N__9665;
    wire N__9662;
    wire N__9661;
    wire N__9658;
    wire N__9655;
    wire N__9650;
    wire N__9647;
    wire N__9646;
    wire N__9643;
    wire N__9640;
    wire N__9635;
    wire N__9632;
    wire N__9631;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9617;
    wire N__9614;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9604;
    wire N__9599;
    wire N__9596;
    wire N__9595;
    wire N__9592;
    wire N__9589;
    wire N__9584;
    wire N__9581;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9568;
    wire N__9565;
    wire N__9564;
    wire N__9561;
    wire N__9560;
    wire N__9557;
    wire N__9552;
    wire N__9549;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9523;
    wire N__9518;
    wire N__9515;
    wire N__9514;
    wire N__9511;
    wire N__9508;
    wire N__9503;
    wire N__9502;
    wire N__9499;
    wire N__9496;
    wire N__9491;
    wire N__9488;
    wire N__9487;
    wire N__9484;
    wire N__9481;
    wire N__9476;
    wire N__9473;
    wire N__9472;
    wire N__9469;
    wire N__9466;
    wire N__9461;
    wire N__9458;
    wire N__9457;
    wire N__9454;
    wire N__9451;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9418;
    wire N__9415;
    wire N__9414;
    wire N__9413;
    wire N__9410;
    wire N__9403;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9391;
    wire N__9388;
    wire N__9387;
    wire N__9384;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9283;
    wire N__9280;
    wire N__9279;
    wire N__9276;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9205;
    wire N__9202;
    wire N__9201;
    wire N__9198;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9166;
    wire N__9163;
    wire N__9162;
    wire N__9159;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9103;
    wire N__9100;
    wire N__9099;
    wire N__9096;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9019;
    wire N__9016;
    wire N__9015;
    wire N__9012;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8917;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8899;
    wire N__8898;
    wire N__8897;
    wire N__8896;
    wire N__8887;
    wire N__8884;
    wire N__8879;
    wire N__8878;
    wire N__8873;
    wire N__8870;
    wire N__8869;
    wire N__8866;
    wire N__8865;
    wire N__8862;
    wire N__8859;
    wire N__8856;
    wire N__8853;
    wire N__8846;
    wire N__8845;
    wire N__8844;
    wire N__8843;
    wire N__8842;
    wire N__8839;
    wire N__8830;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire VCCG0;
    wire \PCH_PWRGD.un4_count_11 ;
    wire \PCH_PWRGD.un4_count_9 ;
    wire \PCH_PWRGD.un4_count_10_cascade_ ;
    wire \PCH_PWRGD.N_1_i_cascade_ ;
    wire \PCH_PWRGD.un1_curr_state_0_sqmuxa_0_cascade_ ;
    wire \PCH_PWRGD.curr_state_RNI7N705Z0Z_0_cascade_ ;
    wire \PCH_PWRGD.un4_count_8 ;
    wire \PCH_PWRGD.N_3_i_cascade_ ;
    wire vr_ready_vccin;
    wire \PCH_PWRGD.curr_stateZ0Z_0 ;
    wire \PCH_PWRGD.N_1_i ;
    wire \PCH_PWRGD.N_3_i ;
    wire \PCH_PWRGD.curr_stateZ0Z_1 ;
    wire bfn_1_5_0_;
    wire \POWERLED.mult1_un89_sum_cry_2 ;
    wire \POWERLED.mult1_un89_sum_cry_3 ;
    wire \POWERLED.mult1_un89_sum_cry_4 ;
    wire \POWERLED.mult1_un89_sum_cry_5 ;
    wire \POWERLED.mult1_un89_sum_cry_6 ;
    wire \POWERLED.mult1_un89_sum_cry_7 ;
    wire \POWERLED.mult1_un89_sum_s_8_cascade_ ;
    wire bfn_1_6_0_;
    wire \POWERLED.mult1_un96_sum_cry_2 ;
    wire \POWERLED.mult1_un89_sum_cry_3_s ;
    wire \POWERLED.mult1_un96_sum_cry_3 ;
    wire \POWERLED.mult1_un89_sum_cry_4_s ;
    wire \POWERLED.mult1_un96_sum_cry_4 ;
    wire \POWERLED.mult1_un89_sum_cry_5_s ;
    wire \POWERLED.mult1_un96_sum_cry_5 ;
    wire \POWERLED.mult1_un89_sum_cry_6_s ;
    wire \POWERLED.mult1_un89_sum_i_0_8 ;
    wire \POWERLED.mult1_un96_sum_cry_6 ;
    wire \POWERLED.mult1_un96_sum_axb_8 ;
    wire \POWERLED.mult1_un96_sum_cry_7 ;
    wire \POWERLED.mult1_un96_sum_s_8_cascade_ ;
    wire bfn_1_7_0_;
    wire \POWERLED.mult1_un103_sum_cry_2 ;
    wire \POWERLED.mult1_un96_sum_cry_3_s ;
    wire \POWERLED.mult1_un103_sum_cry_3 ;
    wire \POWERLED.mult1_un96_sum_cry_4_s ;
    wire \POWERLED.mult1_un103_sum_cry_4 ;
    wire \POWERLED.mult1_un96_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_cry_5 ;
    wire \POWERLED.mult1_un96_sum_cry_6_s ;
    wire \POWERLED.mult1_un96_sum_i_0_8 ;
    wire \POWERLED.mult1_un103_sum_cry_6 ;
    wire \POWERLED.mult1_un103_sum_axb_8 ;
    wire \POWERLED.mult1_un103_sum_cry_7 ;
    wire \POWERLED.mult1_un103_sum_s_8_cascade_ ;
    wire bfn_1_8_0_;
    wire \POWERLED.mult1_un110_sum_cry_2 ;
    wire \POWERLED.mult1_un103_sum_cry_3_s ;
    wire \POWERLED.mult1_un110_sum_cry_3 ;
    wire \POWERLED.mult1_un103_sum_cry_4_s ;
    wire \POWERLED.mult1_un110_sum_cry_4 ;
    wire \POWERLED.mult1_un103_sum_cry_5_s ;
    wire \POWERLED.mult1_un110_sum_cry_5 ;
    wire \POWERLED.mult1_un103_sum_cry_6_s ;
    wire \POWERLED.mult1_un103_sum_i_0_8 ;
    wire \POWERLED.mult1_un110_sum_cry_6 ;
    wire \POWERLED.mult1_un110_sum_axb_8 ;
    wire \POWERLED.mult1_un110_sum_cry_7 ;
    wire \POWERLED.mult1_un110_sum_s_8_cascade_ ;
    wire bfn_1_9_0_;
    wire \POWERLED.mult1_un124_sum_cry_2 ;
    wire \POWERLED.mult1_un124_sum_cry_3 ;
    wire \POWERLED.mult1_un124_sum_cry_4 ;
    wire \POWERLED.mult1_un124_sum_cry_5 ;
    wire \POWERLED.mult1_un124_sum_cry_6 ;
    wire \POWERLED.mult1_un124_sum_cry_7 ;
    wire \POWERLED.mult1_un124_sum_s_8_cascade_ ;
    wire bfn_1_10_0_;
    wire \POWERLED.mult1_un131_sum_cry_2 ;
    wire \POWERLED.mult1_un124_sum_cry_3_s ;
    wire \POWERLED.mult1_un131_sum_cry_3 ;
    wire \POWERLED.mult1_un124_sum_cry_4_s ;
    wire \POWERLED.mult1_un131_sum_cry_4 ;
    wire \POWERLED.mult1_un124_sum_cry_5_s ;
    wire \POWERLED.mult1_un131_sum_cry_5 ;
    wire \POWERLED.mult1_un124_sum_cry_6_s ;
    wire \POWERLED.mult1_un124_sum_i_0_8 ;
    wire \POWERLED.mult1_un131_sum_cry_6 ;
    wire \POWERLED.mult1_un131_sum_axb_8 ;
    wire \POWERLED.mult1_un131_sum_cry_7 ;
    wire \POWERLED.mult1_un131_sum_s_8_cascade_ ;
    wire bfn_1_11_0_;
    wire \POWERLED.mult1_un138_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_cry_3_s ;
    wire \POWERLED.mult1_un138_sum_cry_3 ;
    wire \POWERLED.mult1_un131_sum_cry_4_s ;
    wire \POWERLED.mult1_un138_sum_cry_4 ;
    wire \POWERLED.mult1_un131_sum_cry_5_s ;
    wire \POWERLED.mult1_un138_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_cry_6_s ;
    wire \POWERLED.mult1_un131_sum_i_0_8 ;
    wire \POWERLED.mult1_un138_sum_cry_6 ;
    wire \POWERLED.mult1_un138_sum_axb_8 ;
    wire \POWERLED.mult1_un138_sum_cry_7 ;
    wire \POWERLED.mult1_un138_sum_s_8_cascade_ ;
    wire bfn_1_12_0_;
    wire \POWERLED.mult1_un159_sum_cry_1 ;
    wire \POWERLED.mult1_un159_sum_cry_2 ;
    wire \POWERLED.mult1_un159_sum_cry_3 ;
    wire \POWERLED.mult1_un159_sum_cry_4 ;
    wire \POWERLED.mult1_un159_sum_cry_5 ;
    wire \POWERLED.mult1_un159_sum_cry_6 ;
    wire \POWERLED.mult1_un159_sum_s_7_cascade_ ;
    wire bfn_1_13_0_;
    wire \POWERLED.mult1_un166_sum_cry_0 ;
    wire \POWERLED.mult1_un159_sum_cry_2_s ;
    wire \POWERLED.mult1_un166_sum_cry_1 ;
    wire \POWERLED.mult1_un159_sum_cry_3_s ;
    wire \POWERLED.mult1_un166_sum_cry_2 ;
    wire \POWERLED.mult1_un159_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_s_7 ;
    wire \POWERLED.mult1_un166_sum_cry_3 ;
    wire \POWERLED.mult1_un159_sum_cry_5_s ;
    wire G_407;
    wire \POWERLED.mult1_un166_sum_cry_4 ;
    wire \POWERLED.mult1_un166_sum_axb_6 ;
    wire \POWERLED.mult1_un166_sum_cry_5 ;
    wire \POWERLED.mult1_un96_sum_i ;
    wire \POWERLED.mult1_un96_sum_s_8 ;
    wire pwrbtn_led;
    wire \PCH_PWRGD.un1_curr_state10_0 ;
    wire \PCH_PWRGD.countZ0Z_0 ;
    wire bfn_2_2_0_;
    wire \PCH_PWRGD.countZ0Z_1 ;
    wire \PCH_PWRGD.un1_count_1_cry_0 ;
    wire \PCH_PWRGD.countZ0Z_2 ;
    wire \PCH_PWRGD.un1_count_1_cry_1 ;
    wire \PCH_PWRGD.countZ0Z_3 ;
    wire \PCH_PWRGD.un1_count_1_cry_2 ;
    wire \PCH_PWRGD.countZ0Z_4 ;
    wire \PCH_PWRGD.un1_count_1_cry_3 ;
    wire \PCH_PWRGD.countZ0Z_5 ;
    wire \PCH_PWRGD.un1_count_1_cry_4 ;
    wire \PCH_PWRGD.countZ0Z_6 ;
    wire \PCH_PWRGD.un1_count_1_cry_5 ;
    wire \PCH_PWRGD.countZ0Z_7 ;
    wire \PCH_PWRGD.un1_count_1_cry_6 ;
    wire \PCH_PWRGD.un1_count_1_cry_7 ;
    wire \PCH_PWRGD.countZ0Z_8 ;
    wire bfn_2_3_0_;
    wire \PCH_PWRGD.countZ0Z_9 ;
    wire \PCH_PWRGD.un1_count_1_cry_8 ;
    wire \PCH_PWRGD.countZ0Z_10 ;
    wire \PCH_PWRGD.un1_count_1_cry_9 ;
    wire \PCH_PWRGD.countZ0Z_11 ;
    wire \PCH_PWRGD.un1_count_1_cry_10 ;
    wire \PCH_PWRGD.countZ0Z_12 ;
    wire \PCH_PWRGD.un1_count_1_cry_11 ;
    wire \PCH_PWRGD.countZ0Z_13 ;
    wire \PCH_PWRGD.un1_count_1_cry_12 ;
    wire \PCH_PWRGD.countZ0Z_14 ;
    wire \PCH_PWRGD.un1_count_1_cry_13 ;
    wire \PCH_PWRGD.un1_count_1_cry_14 ;
    wire \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_2_4_0_;
    wire \PCH_PWRGD.countZ0Z_15 ;
    wire \PCH_PWRGD.N_65_3 ;
    wire \PCH_PWRGD.curr_state_RNI7N705Z0Z_0 ;
    wire bfn_2_5_0_;
    wire \POWERLED.mult1_un82_sum_cry_3_s ;
    wire \POWERLED.mult1_un82_sum_cry_2 ;
    wire \POWERLED.mult1_un82_sum_cry_4_s ;
    wire \POWERLED.mult1_un82_sum_cry_3 ;
    wire \POWERLED.mult1_un82_sum_cry_5_s ;
    wire \POWERLED.mult1_un82_sum_cry_4 ;
    wire \POWERLED.mult1_un82_sum_cry_6_s ;
    wire \POWERLED.mult1_un82_sum_cry_5 ;
    wire \POWERLED.mult1_un89_sum_axb_8 ;
    wire \POWERLED.mult1_un82_sum_cry_6 ;
    wire \POWERLED.mult1_un82_sum_cry_7 ;
    wire \POWERLED.mult1_un82_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un82_sum_i_0_8 ;
    wire bfn_2_6_0_;
    wire \POWERLED.mult1_un75_sum_cry_3_s ;
    wire \POWERLED.mult1_un75_sum_cry_2 ;
    wire \POWERLED.mult1_un75_sum_cry_4_s ;
    wire \POWERLED.mult1_un75_sum_cry_3 ;
    wire \POWERLED.mult1_un75_sum_cry_5_s ;
    wire \POWERLED.mult1_un75_sum_cry_4 ;
    wire \POWERLED.mult1_un75_sum_cry_6_s ;
    wire \POWERLED.mult1_un75_sum_cry_5 ;
    wire \POWERLED.mult1_un82_sum_axb_8 ;
    wire \POWERLED.mult1_un75_sum_cry_6 ;
    wire \POWERLED.mult1_un75_sum_cry_7 ;
    wire \POWERLED.mult1_un75_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un75_sum_i_0_8 ;
    wire bfn_2_7_0_;
    wire \POWERLED.mult1_un68_sum_cry_3_s ;
    wire \POWERLED.mult1_un68_sum_cry_2 ;
    wire \POWERLED.mult1_un68_sum_cry_4_s ;
    wire \POWERLED.mult1_un68_sum_cry_3 ;
    wire \POWERLED.mult1_un68_sum_cry_5_s ;
    wire \POWERLED.mult1_un68_sum_cry_4 ;
    wire \POWERLED.mult1_un68_sum_cry_6_s ;
    wire \POWERLED.mult1_un68_sum_cry_5 ;
    wire \POWERLED.mult1_un75_sum_axb_8 ;
    wire \POWERLED.mult1_un68_sum_cry_6 ;
    wire \POWERLED.mult1_un68_sum_cry_7 ;
    wire \POWERLED.mult1_un68_sum_i_0_8 ;
    wire \POWERLED.mult1_un89_sum_s_8 ;
    wire \POWERLED.mult1_un82_sum_s_8 ;
    wire \POWERLED.mult1_un68_sum_s_8 ;
    wire \POWERLED.mult1_un75_sum_s_8 ;
    wire \POWERLED.mult1_un103_sum_i ;
    wire \POWERLED.mult1_un103_sum_s_8 ;
    wire \POWERLED.mult1_un89_sum_i ;
    wire bfn_2_9_0_;
    wire \POWERLED.mult1_un117_sum_cry_3_s ;
    wire \POWERLED.mult1_un117_sum_cry_2 ;
    wire \POWERLED.mult1_un110_sum_cry_3_s ;
    wire \POWERLED.mult1_un117_sum_cry_4_s ;
    wire \POWERLED.mult1_un117_sum_cry_3 ;
    wire \POWERLED.mult1_un110_sum_cry_4_s ;
    wire \POWERLED.mult1_un117_sum_cry_5_s ;
    wire \POWERLED.mult1_un117_sum_cry_4 ;
    wire \POWERLED.mult1_un110_sum_s_8 ;
    wire \POWERLED.mult1_un110_sum_cry_5_s ;
    wire \POWERLED.mult1_un117_sum_cry_6_s ;
    wire \POWERLED.mult1_un117_sum_cry_5 ;
    wire \POWERLED.mult1_un110_sum_cry_6_s ;
    wire \POWERLED.mult1_un110_sum_i_0_8 ;
    wire \POWERLED.mult1_un124_sum_axb_8 ;
    wire \POWERLED.mult1_un117_sum_cry_6 ;
    wire \POWERLED.mult1_un117_sum_axb_8 ;
    wire \POWERLED.mult1_un117_sum_cry_7 ;
    wire \POWERLED.mult1_un117_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un117_sum_i_0_8 ;
    wire \POWERLED.mult1_un124_sum_s_8 ;
    wire \POWERLED.mult1_un131_sum_s_8 ;
    wire \POWERLED.mult1_un131_sum_i ;
    wire \POWERLED.mult1_un117_sum_s_8 ;
    wire bfn_2_11_0_;
    wire \POWERLED.mult1_un138_sum_i_0_8 ;
    wire \POWERLED.mult1_un145_sum_cry_2 ;
    wire \POWERLED.mult1_un138_sum_cry_3_s ;
    wire \POWERLED.mult1_un145_sum_axb_4_l_fx ;
    wire \POWERLED.mult1_un145_sum_cry_3 ;
    wire \POWERLED.mult1_un138_sum_cry_4_s ;
    wire \POWERLED.mult1_un145_sum_cry_4 ;
    wire \POWERLED.mult1_un138_sum_cry_5_s ;
    wire \POWERLED.mult1_un145_sum_cry_5 ;
    wire \POWERLED.mult1_un145_sum_cry_6 ;
    wire \POWERLED.mult1_un145_sum_axb_8 ;
    wire \POWERLED.mult1_un145_sum_cry_7 ;
    wire \POWERLED.mult1_un145_sum_s_8_cascade_ ;
    wire bfn_2_12_0_;
    wire \POWERLED.mult1_un145_sum_i ;
    wire \POWERLED.mult1_un152_sum_cry_3_s ;
    wire \POWERLED.mult1_un152_sum_cry_2 ;
    wire \POWERLED.mult1_un145_sum_cry_3_s ;
    wire \POWERLED.mult1_un152_sum_cry_4_s ;
    wire \POWERLED.mult1_un152_sum_cry_3 ;
    wire \POWERLED.mult1_un145_sum_cry_4_s ;
    wire \POWERLED.mult1_un152_sum_cry_5_s ;
    wire \POWERLED.mult1_un152_sum_cry_4 ;
    wire \POWERLED.mult1_un145_sum_s_8 ;
    wire \POWERLED.mult1_un145_sum_cry_5_s ;
    wire \POWERLED.mult1_un152_sum_cry_6_s ;
    wire \POWERLED.mult1_un152_sum_cry_5 ;
    wire \POWERLED.mult1_un145_sum_cry_6_s ;
    wire \POWERLED.mult1_un145_sum_i_0_8 ;
    wire \POWERLED.mult1_un159_sum_axb_7 ;
    wire \POWERLED.mult1_un152_sum_cry_6 ;
    wire \POWERLED.mult1_un152_sum_axb_8 ;
    wire \POWERLED.mult1_un152_sum_cry_7 ;
    wire \POWERLED.mult1_un152_sum_s_8 ;
    wire \POWERLED.mult1_un152_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un152_sum_i_0_8 ;
    wire \POWERLED.un1_count_2_0 ;
    wire \POWERLED.count_i_0_0 ;
    wire bfn_2_13_0_;
    wire \POWERLED.un1_count_2_1 ;
    wire \POWERLED.count_i_1 ;
    wire \POWERLED.un1_count_2_cry_0 ;
    wire \POWERLED.un1_count_2_2 ;
    wire \POWERLED.count_i_2 ;
    wire \POWERLED.un1_count_2_cry_1 ;
    wire \POWERLED.un1_count_2_3 ;
    wire \POWERLED.count_i_3 ;
    wire \POWERLED.un1_count_2_cry_2 ;
    wire \POWERLED.count_i_4 ;
    wire \POWERLED.un1_count_2_cry_3 ;
    wire \POWERLED.un1_count_2_5 ;
    wire \POWERLED.count_i_5 ;
    wire \POWERLED.un1_count_2_cry_4 ;
    wire \POWERLED.un1_count_2_6 ;
    wire \POWERLED.count_i_6 ;
    wire \POWERLED.un1_count_2_cry_5 ;
    wire \POWERLED.un1_count_2_7 ;
    wire \POWERLED.count_i_7 ;
    wire \POWERLED.un1_count_2_cry_6 ;
    wire \POWERLED.un1_count_2_cry_7 ;
    wire \POWERLED.un1_count_2_8 ;
    wire \POWERLED.count_i_8 ;
    wire bfn_2_14_0_;
    wire \POWERLED.un1_count_2_9 ;
    wire \POWERLED.count_i_9 ;
    wire \POWERLED.un1_count_2_cry_8 ;
    wire \POWERLED.un1_count_2_10 ;
    wire \POWERLED.count_i_10 ;
    wire \POWERLED.un1_count_2_cry_9 ;
    wire \POWERLED.un1_count_2_11 ;
    wire \POWERLED.count_i_11 ;
    wire \POWERLED.un1_count_2_cry_10 ;
    wire \POWERLED.un1_count_2_12 ;
    wire \POWERLED.count_i_12 ;
    wire \POWERLED.un1_count_2_cry_11 ;
    wire \POWERLED.un1_count_2_13 ;
    wire \POWERLED.count_i_13 ;
    wire \POWERLED.un1_count_2_cry_12 ;
    wire \POWERLED.un1_count_2_14 ;
    wire \POWERLED.count_i_14 ;
    wire \POWERLED.un1_count_2_cry_13 ;
    wire \POWERLED.un1_count_2_15 ;
    wire \POWERLED.count_i_15 ;
    wire \POWERLED.un1_count_2_cry_14 ;
    wire \POWERLED.un1_count_2_cry_15 ;
    wire bfn_2_15_0_;
    wire \POWERLED.un1_count_2_cry_15_THRU_CO ;
    wire \POWERLED.un1_count_2_cry_15_THRU_CO_cascade_ ;
    wire \POWERLED.pwm_out_RNOZ0 ;
    wire vpp_ok;
    wire vddq_en;
    wire gpio_fpga_soc_1;
    wire \HDA_STRAP.N_5_0_cascade_ ;
    wire pch_pwrok;
    wire \HDA_STRAP.m14_ns_1 ;
    wire bfn_4_5_0_;
    wire \POWERLED.mult1_un54_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6 ;
    wire \POWERLED.mult1_un54_sum_cry_7 ;
    wire bfn_4_6_0_;
    wire \POWERLED.mult1_un47_sum_cry_3_s ;
    wire \POWERLED.mult1_un47_sum_cry_2 ;
    wire \POWERLED.mult1_un47_sum_cry_4_s ;
    wire \POWERLED.mult1_un47_sum_cry_3 ;
    wire \POWERLED.mult1_un47_sum_cry_5_s ;
    wire \POWERLED.mult1_un47_sum_cry_4 ;
    wire \POWERLED.mult1_un47_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_7_THRU_CO ;
    wire \POWERLED.mult1_un47_sum_cry_6 ;
    wire \POWERLED.mult1_un68_sum_i ;
    wire bfn_4_7_0_;
    wire \POWERLED.mult1_un61_sum_cry_3_s ;
    wire \POWERLED.mult1_un61_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3_s ;
    wire \POWERLED.mult1_un61_sum_cry_4_s ;
    wire \POWERLED.mult1_un61_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4_s ;
    wire \POWERLED.mult1_un61_sum_cry_5_s ;
    wire \POWERLED.mult1_un61_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_cry_5_s ;
    wire \POWERLED.mult1_un61_sum_cry_6_s ;
    wire \POWERLED.mult1_un61_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6_s ;
    wire \POWERLED.mult1_un54_sum_i_8 ;
    wire \POWERLED.mult1_un68_sum_axb_8 ;
    wire \POWERLED.mult1_un61_sum_cry_6 ;
    wire \POWERLED.mult1_un47_sum_cry_6_s ;
    wire \POWERLED.mult1_un54_sum_s_8 ;
    wire \POWERLED.mult1_un54_sum_cry_6_THRU_CO ;
    wire \POWERLED.mult1_un61_sum_cry_7 ;
    wire \POWERLED.mult1_un61_sum_s_8 ;
    wire \POWERLED.mult1_un61_sum_i_0_8 ;
    wire \POWERLED.mult1_un110_sum_i ;
    wire \POWERLED.mult1_un138_sum_i ;
    wire \POWERLED.mult1_un124_sum_i ;
    wire \POWERLED.mult1_un117_sum_i ;
    wire \POWERLED.mult1_un138_sum_cry_6_s ;
    wire \POWERLED.mult1_un145_sum_axb_7_l_fx ;
    wire \POWERLED.mult1_un138_sum_s_8 ;
    wire \POWERLED.un1_count_2_4 ;
    wire v5s_enn;
    wire \POWERLED.mult1_un159_sum_i ;
    wire \POWERLED.mult1_un152_sum_i ;
    wire \POWERLED.un1_countlt6_0_cascade_ ;
    wire \POWERLED.g0_0_7_cascade_ ;
    wire \POWERLED.un1_count_0 ;
    wire \POWERLED.un1_countlto15_5_cascade_ ;
    wire \POWERLED.g0_0_4 ;
    wire \POWERLED.un1_countlt6 ;
    wire \POWERLED.g0_0_5 ;
    wire \POWERLED.un1_countlto15_4_cascade_ ;
    wire \POWERLED.un1_countlto15_7 ;
    wire \POWERLED.count_RNIOVT24Z0Z_11 ;
    wire \POWERLED.curr_stateZ0Z_0 ;
    wire \POWERLED.count_RNIOVT24Z0Z_11_cascade_ ;
    wire \HDA_STRAP.N_5_0 ;
    wire \HDA_STRAP.curr_stateZ0Z_2 ;
    wire hda_sdo_atp;
    wire \POWERLED.mult1_un82_sum_i ;
    wire \POWERLED.un1_dutycycle_1_i_28 ;
    wire \POWERLED.un1_dutycycle_1_19_0_cascade_ ;
    wire \POWERLED.mult1_un75_sum_i ;
    wire \POWERLED.N_53 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_4 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_5 ;
    wire \POWERLED.mult1_un47_sum_axb_4 ;
    wire \POWERLED.un1_dutycycle_1_i_29 ;
    wire \POWERLED.mult1_un61_sum_i ;
    wire \POWERLED.mult1_un54_sum_i ;
    wire bfn_5_9_0_;
    wire \POWERLED.un1_count_off_1_cry_0 ;
    wire \POWERLED.un1_count_off_1_cry_1 ;
    wire \POWERLED.un1_count_off_1_cry_2 ;
    wire \POWERLED.un1_count_off_1_cry_3 ;
    wire \POWERLED.un1_count_off_1_cry_4 ;
    wire \POWERLED.un1_count_off_1_cry_5 ;
    wire \POWERLED.un1_count_off_1_cry_6 ;
    wire \POWERLED.un1_count_off_1_cry_7 ;
    wire bfn_5_10_0_;
    wire \POWERLED.un1_count_off_1_cry_8 ;
    wire \POWERLED.un1_count_off_1_cry_9 ;
    wire \POWERLED.un1_count_off_1_cry_10 ;
    wire \POWERLED.un1_count_off_1_cry_11 ;
    wire \POWERLED.un1_count_off_1_cry_12 ;
    wire \POWERLED.un1_count_off_1_cry_13 ;
    wire \POWERLED.un1_count_off_1_cry_14 ;
    wire \POWERLED.count_offZ0Z_12 ;
    wire \POWERLED.count_offZ0Z_13 ;
    wire \POWERLED.count_offZ0Z_15 ;
    wire \POWERLED.count_offZ0Z_1 ;
    wire \POWERLED.count_offZ0Z_11 ;
    wire \POWERLED.count_offZ0Z_0 ;
    wire \POWERLED.count_offZ0Z_14 ;
    wire \POWERLED.count_offZ0Z_10 ;
    wire \POWERLED.count_offZ0Z_8 ;
    wire \POWERLED.count_offZ0Z_6 ;
    wire \POWERLED.count_offZ0Z_9 ;
    wire \POWERLED.count_offZ0Z_5 ;
    wire \POWERLED.func_state_ns_0_a2_11_0 ;
    wire \POWERLED.func_state_ns_0_a2_10_0 ;
    wire \POWERLED.func_state_ns_0_a2_9_0_cascade_ ;
    wire \POWERLED.count_off_0_sqmuxa ;
    wire \POWERLED.count_off_0_sqmuxa_cascade_ ;
    wire \POWERLED.N_85_1 ;
    wire \POWERLED.countZ0Z_0 ;
    wire \POWERLED.countZ0Z_1 ;
    wire bfn_5_14_0_;
    wire \POWERLED.countZ0Z_2 ;
    wire \POWERLED.un1_count_1_cry_1 ;
    wire \POWERLED.countZ0Z_3 ;
    wire \POWERLED.un1_count_1_cry_2 ;
    wire \POWERLED.countZ0Z_4 ;
    wire \POWERLED.un1_count_1_cry_3 ;
    wire \POWERLED.countZ0Z_5 ;
    wire \POWERLED.un1_count_1_cry_4 ;
    wire \POWERLED.countZ0Z_6 ;
    wire \POWERLED.un1_count_1_cry_5 ;
    wire \POWERLED.countZ0Z_7 ;
    wire \POWERLED.un1_count_1_cry_6 ;
    wire \POWERLED.countZ0Z_8 ;
    wire \POWERLED.un1_count_1_cry_7 ;
    wire \POWERLED.un1_count_1_cry_8 ;
    wire \POWERLED.countZ0Z_9 ;
    wire bfn_5_15_0_;
    wire \POWERLED.countZ0Z_10 ;
    wire \POWERLED.un1_count_1_cry_9 ;
    wire \POWERLED.countZ0Z_11 ;
    wire \POWERLED.un1_count_1_cry_10 ;
    wire \POWERLED.countZ0Z_12 ;
    wire \POWERLED.un1_count_1_cry_11 ;
    wire \POWERLED.countZ0Z_13 ;
    wire \POWERLED.un1_count_1_cry_12 ;
    wire \POWERLED.countZ0Z_14 ;
    wire \POWERLED.un1_count_1_cry_13 ;
    wire \POWERLED.un1_count_1_cry_14 ;
    wire \POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire \POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO ;
    wire bfn_5_16_0_;
    wire \POWERLED.countZ0Z_15 ;
    wire \POWERLED.N_65_5 ;
    wire \POWERLED.curr_state_RNI75RB5Z0Z_0 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_0 ;
    wire bfn_6_1_0_;
    wire \HDA_STRAP.un1_count_1_cry_0 ;
    wire \HDA_STRAP.un1_count_1_cry_1 ;
    wire \HDA_STRAP.un1_count_1_cry_2 ;
    wire \HDA_STRAP.un1_count_1_cry_3 ;
    wire \HDA_STRAP.un1_count_1_cry_4 ;
    wire \HDA_STRAP.un1_count_1_cry_5 ;
    wire \HDA_STRAP.un1_count_1_cry_6 ;
    wire \HDA_STRAP.un1_count_1_cry_7 ;
    wire bfn_6_2_0_;
    wire \HDA_STRAP.un1_count_1_cry_8 ;
    wire \HDA_STRAP.un1_count_1_cry_9 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_11 ;
    wire \HDA_STRAP.un1_count_1_cry_10 ;
    wire \HDA_STRAP.un1_count_1_cry_11 ;
    wire \HDA_STRAP.un1_count_1_cry_12 ;
    wire \HDA_STRAP.un1_count_1_cry_13 ;
    wire \HDA_STRAP.un1_count_1_cry_14 ;
    wire \HDA_STRAP.un1_count_1_cry_15 ;
    wire bfn_6_3_0_;
    wire \HDA_STRAP.un1_count_1_cry_16 ;
    wire \POWERLED.un1_dutycycle_1_axb_0 ;
    wire bfn_6_5_0_;
    wire \POWERLED.un1_dutycycle_1_axb_1 ;
    wire \POWERLED.mult1_un138_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_0 ;
    wire \POWERLED.dutycycle_RNI16B71Z0Z_5 ;
    wire \POWERLED.dutycycle_RNIFHLJZ0Z_0 ;
    wire \POWERLED.mult1_un131_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_1 ;
    wire \POWERLED.mult1_un124_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_2 ;
    wire \POWERLED.mult1_un117_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_3 ;
    wire \POWERLED.dutycycle_RNIEJ021Z0Z_4 ;
    wire \POWERLED.mult1_un110_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_4 ;
    wire \POWERLED.dutycycle_RNI6NI81Z0Z_5 ;
    wire \POWERLED.mult1_un103_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_5 ;
    wire \POWERLED.dutycycle_RNIJNBA1Z0Z_6 ;
    wire \POWERLED.mult1_un96_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_6 ;
    wire \POWERLED.un1_dutycycle_1_cry_7 ;
    wire \POWERLED.mult1_un89_sum ;
    wire bfn_6_6_0_;
    wire \POWERLED.mult1_un82_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_8 ;
    wire \POWERLED.mult1_un75_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_9 ;
    wire \POWERLED.mult1_un68_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_10 ;
    wire \POWERLED.mult1_un61_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_11 ;
    wire \POWERLED.mult1_un54_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_12 ;
    wire \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1 ;
    wire \POWERLED.un1_dutycycle_1_cry_13 ;
    wire \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1 ;
    wire \POWERLED.un1_dutycycle_1_cry_14 ;
    wire \POWERLED.un1_dutycycle_1_cry_15 ;
    wire \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71 ;
    wire bfn_6_7_0_;
    wire \POWERLED.CO2 ;
    wire \POWERLED.CO2_THRU_CO ;
    wire \POWERLED.dutycycle_fastZ0Z_5 ;
    wire \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5 ;
    wire \POWERLED.dutycycle_RNIE4FLZ0Z_9 ;
    wire \POWERLED.dutycycle_RNI53MGZ0Z_14 ;
    wire \POWERLED.dutycycle_RNI84C11Z0Z_14 ;
    wire \POWERLED.dutycycle_RNIB1FLZ0Z_8 ;
    wire \POWERLED.dutycycle_RNI75MGZ0Z_15 ;
    wire \POWERLED.un1_dutycycle_1_34_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_1_axb_8_cascade_ ;
    wire \POWERLED.dutycycle_fast_RNILMLMZ0Z_6 ;
    wire \POWERLED.dutycycle_RNIJL1R1Z0Z_6 ;
    wire \POWERLED.dutycycle_fastZ0Z_6 ;
    wire \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6 ;
    wire \POWERLED.dutycycle_RNI2V0PZ0Z_10 ;
    wire \POWERLED.dutycycle_RNI2V0PZ0Z_10_cascade_ ;
    wire \POWERLED.dutycycle_RNI712I1Z0Z_15 ;
    wire \POWERLED.dutycycle_RNIQ09G1Z0Z_10 ;
    wire \POWERLED.count_offZ0Z_3 ;
    wire \POWERLED.count_offZ0Z_7 ;
    wire \POWERLED.count_offZ0Z_4 ;
    wire \POWERLED.count_offZ0Z_2 ;
    wire \POWERLED.func_state_ns_0_a2_8_0 ;
    wire \POWERLED.un1_dutycycle_1_44_0_cascade_ ;
    wire \POWERLED.dutycycle_RNIF3561Z0Z_9 ;
    wire \POWERLED.dutycycle_RNIC8C11Z0Z_15 ;
    wire \POWERLED.dutycycle_RNI73C11Z0Z_15 ;
    wire \POWERLED.N_368_0_i_i_a6_0 ;
    wire \POWERLED.N_207_cascade_ ;
    wire \POWERLED.N_48 ;
    wire \POWERLED.N_149 ;
    wire \POWERLED.N_149_cascade_ ;
    wire \POWERLED.N_214 ;
    wire \POWERLED.N_213 ;
    wire \POWERLED.N_234 ;
    wire \POWERLED.N_218_cascade_ ;
    wire \POWERLED.N_248 ;
    wire \POWERLED.N_88_cascade_ ;
    wire \POWERLED.N_208_cascade_ ;
    wire \POWERLED.func_state_ns_i_0_1_1 ;
    wire \POWERLED.N_222 ;
    wire \POWERLED.N_222_cascade_ ;
    wire \POWERLED.N_228 ;
    wire \POWERLED.N_211_cascade_ ;
    wire \POWERLED.func_state_ns_i_0_0_1 ;
    wire \POWERLED.N_179 ;
    wire \POWERLED.N_178 ;
    wire \POWERLED.N_180 ;
    wire \POWERLED.N_250 ;
    wire \HDA_STRAP.curr_state_RNIH91AZ0Z_0 ;
    wire \HDA_STRAP.countZ0Z_2 ;
    wire \HDA_STRAP.countZ0Z_1 ;
    wire \HDA_STRAP.countZ0Z_3 ;
    wire \HDA_STRAP.countZ0Z_0 ;
    wire \HDA_STRAP.countZ0Z_14 ;
    wire \HDA_STRAP.countZ0Z_15 ;
    wire \HDA_STRAP.countZ0Z_12 ;
    wire \HDA_STRAP.un4_count_9_cascade_ ;
    wire \HDA_STRAP.countZ0Z_13 ;
    wire \HDA_STRAP.countZ0Z_7 ;
    wire \HDA_STRAP.countZ0Z_5 ;
    wire \HDA_STRAP.countZ0Z_9 ;
    wire \HDA_STRAP.countZ0Z_4 ;
    wire \HDA_STRAP.countZ0Z_11 ;
    wire \HDA_STRAP.un4_count_12 ;
    wire \HDA_STRAP.un4_count_11 ;
    wire \HDA_STRAP.un4_count_10_cascade_ ;
    wire \HDA_STRAP.un4_count_13 ;
    wire \HDA_STRAP.count_RNIB5IA5Z0Z_0_cascade_ ;
    wire \HDA_STRAP.curr_state_RNO_0Z0Z_2 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_10 ;
    wire \HDA_STRAP.countZ0Z_10 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_16 ;
    wire \HDA_STRAP.countZ0Z_16 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_17 ;
    wire \HDA_STRAP.countZ0Z_17 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_8 ;
    wire \HDA_STRAP.countZ0Z_8 ;
    wire \POWERLED.dutycycle_RNI31MG_0Z0Z_12 ;
    wire \POWERLED.dutycycle_RNI31MGZ0Z_12 ;
    wire \POWERLED.un1_dutycycle_1_39_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI34C41Z0Z_8 ;
    wire \POWERLED.N_117 ;
    wire \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5 ;
    wire \POWERLED.dutycycle_RNIK4I81Z0Z_6 ;
    wire \POWERLED.dutycycle_lm_0_1_2 ;
    wire \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6 ;
    wire \POWERLED.dutycycle_RNIQAI81Z0Z_4 ;
    wire \POWERLED.dutycycle_RNIOQLJZ0Z_4 ;
    wire bfn_7_7_0_;
    wire \POWERLED.dutycycleZ0Z_0 ;
    wire \POWERLED.dutycycle_s_0 ;
    wire \POWERLED.dutycycle_cry_c_0_THRU_CO ;
    wire \POWERLED.dutycycleZ0Z_1 ;
    wire \POWERLED.dutycycle_s_1 ;
    wire \POWERLED.dutycycle_cry_0 ;
    wire \POWERLED.dutycycleZ0Z_2 ;
    wire \POWERLED.dutycycle_s_2 ;
    wire \POWERLED.dutycycle_cry_1 ;
    wire \POWERLED.dutycycleZ0Z_3 ;
    wire \POWERLED.dutycycle_cry_2 ;
    wire \POWERLED.dutycycleZ0Z_4 ;
    wire \POWERLED.dutycycle_cry_3 ;
    wire \POWERLED.dutycycleZ0Z_5 ;
    wire \POWERLED.dutycycle_s_5 ;
    wire \POWERLED.dutycycle_cry_4 ;
    wire \POWERLED.dutycycleZ0Z_6 ;
    wire \POWERLED.dutycycle_s_6 ;
    wire \POWERLED.dutycycle_cry_5 ;
    wire \POWERLED.dutycycle_cry_6 ;
    wire \POWERLED.dutycycleZ0Z_7 ;
    wire bfn_7_8_0_;
    wire \POWERLED.dutycycle_cry_7 ;
    wire \POWERLED.dutycycle_cry_8 ;
    wire \POWERLED.dutycycle_cry_9 ;
    wire \POWERLED.dutycycle_cry_10 ;
    wire \POWERLED.dutycycle_cry_11 ;
    wire \POWERLED.dutycycle_cry_12 ;
    wire \POWERLED.dutycycle_cry_13 ;
    wire \POWERLED.dutycycle_cry_14 ;
    wire \POWERLED.N_177 ;
    wire bfn_7_9_0_;
    wire \POWERLED.N_246_cascade_ ;
    wire \POWERLED.N_203_4 ;
    wire \POWERLED.N_203_4_cascade_ ;
    wire \POWERLED.N_203_cascade_ ;
    wire \POWERLED.N_251_cascade_ ;
    wire \POWERLED.un2_slp_s3n_2_0_1_0 ;
    wire \POWERLED.count_clk_139_tz_0 ;
    wire \POWERLED.un2_slp_s3n_2_0_cascade_ ;
    wire \POWERLED.N_246 ;
    wire \POWERLED.N_205 ;
    wire \POWERLED.un2_slp_s3n_2_0_a6_3_0_cascade_ ;
    wire \POWERLED.un2_slp_s3n_2_0_1 ;
    wire \POWERLED.N_127 ;
    wire \POWERLED.count_clk_1_sqmuxa_5_0_1 ;
    wire \POWERLED.N_127_cascade_ ;
    wire \POWERLED.count_clk_1_sqmuxa_5_0_0 ;
    wire \POWERLED.N_88 ;
    wire \POWERLED.dutycycle_3_sqmuxa_1_i_0_1_1_cascade_ ;
    wire \POWERLED.N_200_2 ;
    wire \POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_1 ;
    wire \POWERLED.N_366_1_cascade_ ;
    wire \POWERLED.N_251 ;
    wire \POWERLED.dutycycle ;
    wire \POWERLED.N_243 ;
    wire slp_s4n;
    wire \POWERLED.func_stateZ0Z_1 ;
    wire \POWERLED.func_stateZ0Z_0 ;
    wire \POWERLED.count_off_RNIIKVR3Z0Z_10 ;
    wire \POWERLED.N_148 ;
    wire slp_s3n;
    wire vccst_en;
    wire vpp_en;
    wire N_55;
    wire \VPP_VDDQ.N_238 ;
    wire \VPP_VDDQ.N_238_cascade_ ;
    wire \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_ ;
    wire \VPP_VDDQ.G_127_0 ;
    wire \VPP_VDDQ.delayed_vddq_pwrgdZ0 ;
    wire \VPP_VDDQ.curr_stateZ0Z_1 ;
    wire \VPP_VDDQ.curr_stateZ0Z_0 ;
    wire \VPP_VDDQ.N_128 ;
    wire \VPP_VDDQ.N_154_cascade_ ;
    wire \HDA_STRAP.count_RNO_0Z0Z_6 ;
    wire \HDA_STRAP.curr_stateZ0Z_1 ;
    wire \HDA_STRAP.curr_stateZ0Z_0 ;
    wire \HDA_STRAP.count_RNIB5IA5Z0Z_0 ;
    wire \HDA_STRAP.countZ0Z_6 ;
    wire bfn_8_5_0_;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_0 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_1 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_2 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_3 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_4 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_5 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_6 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_7 ;
    wire bfn_8_6_0_;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_8 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_9 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_10 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_11 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_12 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_13 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_14 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_8_7_0_;
    wire \POWERLED.dutycycle_RNIO18NZ0Z_9 ;
    wire \POWERLED.dutycycleZ0Z_13 ;
    wire \POWERLED.dutycycleZ0Z_12 ;
    wire \POWERLED.dutycycleZ0Z_14 ;
    wire \POWERLED.dutycycleZ0Z_10 ;
    wire \POWERLED.dutycycleZ0Z_9 ;
    wire \POWERLED.dutycycleZ0Z_11 ;
    wire \POWERLED.dutycycleZ0Z_15 ;
    wire \POWERLED.dutycycleZ0Z_8 ;
    wire \POWERLED.un2_slp_s3n_2_0_o2_3_7 ;
    wire \POWERLED.un2_slp_s3n_2_0_o2_3_8_cascade_ ;
    wire \POWERLED.un2_slp_s3n_2_0_o2_3_6 ;
    wire \POWERLED.N_112 ;
    wire \POWERLED.N_366_1 ;
    wire \POWERLED.un1_dutycycle_4_sqmuxa_0 ;
    wire \POWERLED.N_177_5 ;
    wire \POWERLED.count_clk_0_sqmuxa_5_0_o2_0_0_cascade_ ;
    wire \POWERLED.N_141 ;
    wire \POWERLED.N_136_cascade_ ;
    wire \POWERLED.N_146 ;
    wire \POWERLED.count_clk_0_sqmuxa_5_0_a6_1 ;
    wire \POWERLED.count_clk_0_sqmuxa_5_0_o2_4 ;
    wire gpio_fpga_soc_4;
    wire \POWERLED.count_off_1_sqmuxa_i_a6_0_1_cascade_ ;
    wire \POWERLED.N_136 ;
    wire \POWERLED.count_off_1_sqmuxa_i_a6_0_3 ;
    wire bfn_8_11_0_;
    wire \RSMRST_PWRGD.un1_count_1_cry_0 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_1 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_2 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_3 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_4 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_5 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_6 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_7 ;
    wire bfn_8_12_0_;
    wire \RSMRST_PWRGD.un1_count_1_cry_8 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_9 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_10 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_11 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_12 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_13 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_8_13_0_;
    wire \VPP_VDDQ.N_108_i ;
    wire bfn_8_14_0_;
    wire \VPP_VDDQ.un1_count_1_cry_0 ;
    wire \VPP_VDDQ.un1_count_1_cry_1 ;
    wire \VPP_VDDQ.un1_count_1_cry_2 ;
    wire \VPP_VDDQ.un1_count_1_cry_3 ;
    wire \VPP_VDDQ.un1_count_1_cry_4 ;
    wire \VPP_VDDQ.un1_count_1_cry_5 ;
    wire \VPP_VDDQ.un1_count_1_cry_6 ;
    wire \VPP_VDDQ.un1_count_1_cry_7 ;
    wire bfn_8_15_0_;
    wire \VPP_VDDQ.un1_count_1_cry_8 ;
    wire \VPP_VDDQ.un1_count_1_cry_9 ;
    wire \VPP_VDDQ.un1_count_1_cry_10 ;
    wire \VPP_VDDQ.un1_count_1_cry_11 ;
    wire \VPP_VDDQ.un1_count_1_cry_12 ;
    wire \VPP_VDDQ.un1_count_1_cry_13 ;
    wire \VPP_VDDQ.un1_count_1_cry_14 ;
    wire \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_8_16_0_;
    wire \VPP_VDDQ.N_65_1 ;
    wire \VPP_VDDQ.curr_state_RNIGR9S7Z0Z_0 ;
    wire \COUNTER.counterZ0Z_1 ;
    wire bfn_9_1_0_;
    wire \COUNTER.counter_1_cry_1 ;
    wire \COUNTER.counter_1_cry_2 ;
    wire \COUNTER.counter_1_cry_3 ;
    wire \COUNTER.counterZ0Z_5 ;
    wire \COUNTER.counter_1_cry_4_THRU_CO ;
    wire \COUNTER.counter_1_cry_4 ;
    wire \COUNTER.counterZ0Z_6 ;
    wire \COUNTER.counter_1_cry_5_THRU_CO ;
    wire \COUNTER.counter_1_cry_5 ;
    wire \COUNTER.counterZ0Z_7 ;
    wire \COUNTER.counter_1_cry_6 ;
    wire \COUNTER.counter_1_cry_7 ;
    wire \COUNTER.counter_1_cry_8 ;
    wire bfn_9_2_0_;
    wire \COUNTER.counter_1_cry_9 ;
    wire \COUNTER.counter_1_cry_10 ;
    wire \COUNTER.counter_1_cry_11 ;
    wire \COUNTER.counter_1_cry_12 ;
    wire \COUNTER.counter_1_cry_13 ;
    wire \COUNTER.counter_1_cry_14 ;
    wire \COUNTER.counter_1_cry_15 ;
    wire \COUNTER.counter_1_cry_16 ;
    wire bfn_9_3_0_;
    wire \COUNTER.counter_1_cry_17 ;
    wire \COUNTER.counter_1_cry_18 ;
    wire \COUNTER.counter_1_cry_19 ;
    wire \COUNTER.counter_1_cry_20 ;
    wire \COUNTER.counter_1_cry_21 ;
    wire \COUNTER.counter_1_cry_22 ;
    wire \COUNTER.counter_1_cry_23 ;
    wire \COUNTER.counter_1_cry_24 ;
    wire bfn_9_4_0_;
    wire \COUNTER.counter_1_cry_25 ;
    wire \COUNTER.counter_1_cry_26 ;
    wire \COUNTER.counter_1_cry_27 ;
    wire \COUNTER.counter_1_cry_28 ;
    wire \COUNTER.counter_1_cry_29 ;
    wire \COUNTER.counter_1_cry_30 ;
    wire \COUNTER.counterZ0Z_22 ;
    wire \COUNTER.counterZ0Z_21 ;
    wire \COUNTER.counterZ0Z_23 ;
    wire \COUNTER.counterZ0Z_20 ;
    wire \ALL_SYS_PWRGD.countZ0Z_5 ;
    wire \ALL_SYS_PWRGD.countZ0Z_3 ;
    wire \ALL_SYS_PWRGD.countZ0Z_11 ;
    wire \ALL_SYS_PWRGD.countZ0Z_2 ;
    wire \COUNTER.counterZ0Z_26 ;
    wire \COUNTER.counterZ0Z_25 ;
    wire \COUNTER.counterZ0Z_27 ;
    wire \COUNTER.counterZ0Z_24 ;
    wire \COUNTER.counterZ0Z_30 ;
    wire \COUNTER.counterZ0Z_28 ;
    wire \COUNTER.counterZ0Z_29 ;
    wire \COUNTER.counterZ0Z_31 ;
    wire \COUNTER.counter_1_cry_3_THRU_CO ;
    wire \COUNTER.counterZ0Z_4 ;
    wire \COUNTER.counterZ0Z_0 ;
    wire \COUNTER.counter_1_cry_1_THRU_CO ;
    wire \COUNTER.counterZ0Z_2 ;
    wire \COUNTER.counter_1_cry_2_THRU_CO ;
    wire \COUNTER.counterZ0Z_3 ;
    wire \ALL_SYS_PWRGD.countZ0Z_7 ;
    wire \ALL_SYS_PWRGD.countZ0Z_8 ;
    wire \ALL_SYS_PWRGD.countZ0Z_6 ;
    wire \ALL_SYS_PWRGD.countZ0Z_4 ;
    wire \ALL_SYS_PWRGD.countZ0Z_14 ;
    wire \ALL_SYS_PWRGD.countZ0Z_15 ;
    wire \ALL_SYS_PWRGD.countZ0Z_13 ;
    wire \ALL_SYS_PWRGD.countZ0Z_12 ;
    wire \ALL_SYS_PWRGD.un4_count_10 ;
    wire \ALL_SYS_PWRGD.un4_count_11_cascade_ ;
    wire \ALL_SYS_PWRGD.un4_count_8 ;
    wire \ALL_SYS_PWRGD.countZ0Z_1 ;
    wire \ALL_SYS_PWRGD.countZ0Z_9 ;
    wire \ALL_SYS_PWRGD.countZ0Z_10 ;
    wire \ALL_SYS_PWRGD.countZ0Z_0 ;
    wire \ALL_SYS_PWRGD.un4_count_9 ;
    wire \ALL_SYS_PWRGD.curr_state_RNIKNST6Z0Z_0 ;
    wire \ALL_SYS_PWRGD.curr_state_RNIKNST6Z0Z_0_cascade_ ;
    wire \ALL_SYS_PWRGD.N_65_4 ;
    wire slp_susn;
    wire v5a_ok;
    wire v33a_ok;
    wire v1p8a_ok;
    wire \COUNTER.tmp_i ;
    wire tmp_RNIRH3P;
    wire \POWERLED.count_clk_1_sqmuxa_5_i ;
    wire \POWERLED.count_clkZ0Z_0 ;
    wire bfn_9_9_0_;
    wire \POWERLED.count_clkZ0Z_1 ;
    wire \POWERLED.un1_count_clk_1_cry_0 ;
    wire \POWERLED.count_clkZ0Z_2 ;
    wire \POWERLED.un1_count_clk_1_cry_1 ;
    wire \POWERLED.count_clkZ0Z_3 ;
    wire \POWERLED.un1_count_clk_1_cry_2 ;
    wire \POWERLED.count_clkZ0Z_4 ;
    wire \POWERLED.un1_count_clk_1_cry_3 ;
    wire \POWERLED.count_clkZ0Z_5 ;
    wire \POWERLED.un1_count_clk_1_cry_4 ;
    wire \POWERLED.count_clkZ0Z_6 ;
    wire \POWERLED.un1_count_clk_1_cry_5 ;
    wire \POWERLED.count_clkZ0Z_7 ;
    wire \POWERLED.un1_count_clk_1_cry_6 ;
    wire \POWERLED.un1_count_clk_1_cry_7 ;
    wire \POWERLED.count_clkZ0Z_8 ;
    wire bfn_9_10_0_;
    wire \POWERLED.count_clkZ0Z_9 ;
    wire \POWERLED.un1_count_clk_1_cry_8 ;
    wire \POWERLED.count_clkZ0Z_10 ;
    wire \POWERLED.un1_count_clk_1_cry_9 ;
    wire \POWERLED.count_clkZ0Z_11 ;
    wire \POWERLED.un1_count_clk_1_cry_10 ;
    wire \POWERLED.count_clkZ0Z_12 ;
    wire \POWERLED.un1_count_clk_1_cry_11 ;
    wire \POWERLED.count_clkZ0Z_13 ;
    wire \POWERLED.un1_count_clk_1_cry_12 ;
    wire \POWERLED.count_clkZ0Z_14 ;
    wire \POWERLED.un1_count_clk_1_cry_13 ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \POWERLED.un1_count_clk_1_cry_14 ;
    wire \POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_9_11_0_;
    wire \POWERLED.count_clkZ0Z_15 ;
    wire \POWERLED.N_65_0 ;
    wire \POWERLED.count_clk_RNIOH1J11Z0Z_7 ;
    wire \RSMRST_PWRGD.countZ0Z_11 ;
    wire \RSMRST_PWRGD.countZ0Z_10 ;
    wire \RSMRST_PWRGD.countZ0Z_13 ;
    wire \RSMRST_PWRGD.countZ0Z_6 ;
    wire \RSMRST_PWRGD.countZ0Z_0 ;
    wire \RSMRST_PWRGD.countZ0Z_8 ;
    wire \RSMRST_PWRGD.countZ0Z_9 ;
    wire \RSMRST_PWRGD.countZ0Z_12 ;
    wire \RSMRST_PWRGD.m4_i_i_a2_0_11 ;
    wire \RSMRST_PWRGD.m4_i_i_a2_0_9_cascade_ ;
    wire \RSMRST_PWRGD.countZ0Z_15 ;
    wire \RSMRST_PWRGD.countZ0Z_14 ;
    wire \RSMRST_PWRGD.countZ0Z_7 ;
    wire \RSMRST_PWRGD.m4_i_i_a2_0_7_cascade_ ;
    wire \RSMRST_PWRGD.countZ0Z_3 ;
    wire \RSMRST_PWRGD.m4_i_i_a2_0_12 ;
    wire \RSMRST_PWRGD.countZ0Z_4 ;
    wire \RSMRST_PWRGD.countZ0Z_2 ;
    wire \RSMRST_PWRGD.countZ0Z_5 ;
    wire \RSMRST_PWRGD.countZ0Z_1 ;
    wire \RSMRST_PWRGD.m4_i_i_a2_0_10 ;
    wire \RSMRST_PWRGD.N_240_cascade_ ;
    wire \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0 ;
    wire \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0_cascade_ ;
    wire \RSMRST_PWRGD.N_65_2 ;
    wire \RSMRST_PWRGD.N_37 ;
    wire \VPP_VDDQ.countZ0Z_5 ;
    wire \VPP_VDDQ.countZ0Z_4 ;
    wire \VPP_VDDQ.countZ0Z_7 ;
    wire \VPP_VDDQ.countZ0Z_3 ;
    wire \VPP_VDDQ.countZ0Z_14 ;
    wire \VPP_VDDQ.countZ0Z_15 ;
    wire \VPP_VDDQ.countZ0Z_13 ;
    wire \VPP_VDDQ.countZ0Z_12 ;
    wire \VPP_VDDQ.countZ0Z_6 ;
    wire \VPP_VDDQ.countZ0Z_2 ;
    wire \VPP_VDDQ.countZ0Z_10 ;
    wire \VPP_VDDQ.countZ0Z_1 ;
    wire \VPP_VDDQ.countZ0Z_9 ;
    wire \VPP_VDDQ.countZ0Z_8 ;
    wire \VPP_VDDQ.countZ0Z_11 ;
    wire \VPP_VDDQ.countZ0Z_0 ;
    wire \VPP_VDDQ.un6_count_11 ;
    wire \VPP_VDDQ.un6_count_10 ;
    wire \VPP_VDDQ.un6_count_9_cascade_ ;
    wire \VPP_VDDQ.un6_count_8 ;
    wire \VPP_VDDQ.count_esr_RNIRFM64Z0Z_15 ;
    wire \COUNTER.counterZ0Z_14 ;
    wire \COUNTER.counterZ0Z_13 ;
    wire \COUNTER.counterZ0Z_15 ;
    wire \COUNTER.counterZ0Z_12 ;
    wire \COUNTER.counterZ0Z_18 ;
    wire \COUNTER.counterZ0Z_17 ;
    wire \COUNTER.counterZ0Z_19 ;
    wire \COUNTER.counterZ0Z_16 ;
    wire \COUNTER.counterZ0Z_10 ;
    wire \COUNTER.counterZ0Z_9 ;
    wire \COUNTER.counterZ0Z_11 ;
    wire \COUNTER.counterZ0Z_8 ;
    wire \COUNTER.un4_counter_0_and ;
    wire bfn_11_5_0_;
    wire \COUNTER.un4_counter_1_and ;
    wire \COUNTER.un4_counter_0 ;
    wire \COUNTER.un4_counter_2_and ;
    wire \COUNTER.un4_counter_1 ;
    wire \COUNTER.un4_counter_3_and ;
    wire \COUNTER.un4_counter_2 ;
    wire \COUNTER.un4_counter_4_and ;
    wire \COUNTER.un4_counter_3 ;
    wire \COUNTER.un4_counter_5_and ;
    wire \COUNTER.un4_counter_4 ;
    wire \COUNTER.un4_counter_6_and ;
    wire \COUNTER.un4_counter_5 ;
    wire \COUNTER.un4_counter_7_and ;
    wire \COUNTER.un4_counter_6 ;
    wire \COUNTER.un4_counter_7 ;
    wire bfn_11_6_0_;
    wire \COUNTER.un4_counter_7_THRU_CO ;
    wire \ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa_cascade_ ;
    wire \ALL_SYS_PWRGD.un1_curr_state10_0 ;
    wire \ALL_SYS_PWRGD.N_1_i ;
    wire \ALL_SYS_PWRGD.N_36 ;
    wire \ALL_SYS_PWRGD.curr_stateZ0Z_0 ;
    wire \ALL_SYS_PWRGD.curr_stateZ0Z_1 ;
    wire vccst_pwrgd;
    wire \RSMRST_PWRGD.curr_stateZ0Z_1 ;
    wire \RSMRST_PWRGD.N_241 ;
    wire \RSMRST_PWRGD.N_240 ;
    wire \RSMRST_PWRGD.curr_stateZ0Z_0 ;
    wire rsmrstn;
    wire fpga_osc;
    wire N_65_g;
    wire vddq_ok;
    wire v5s_ok;
    wire rsmrst_pwrgd_signal;
    wire vccst_cpu_ok;
    wire \ALL_SYS_PWRGD.m4_0_0_a2_1_cascade_ ;
    wire v33s_ok;
    wire \ALL_SYS_PWRGD.N_245 ;
    wire _gnd_net_;

    defparam ipInertedIOPad_VR_READY_VCCINAUX_iopad.PULLUP=1'b0;
    IO_PAD ipInertedIOPad_VR_READY_VCCINAUX_iopad (
            .OE(N__21309),
            .DIN(N__21308),
            .DOUT(N__21307),
            .PACKAGEPIN(VR_READY_VCCINAUX));
    defparam ipInertedIOPad_VR_READY_VCCINAUX_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCINAUX_preio (
            .PADOEN(N__21309),
            .PADOUT(N__21308),
            .PADIN(N__21307),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_ENn_iopad (
            .OE(N__21300),
            .DIN(N__21299),
            .DOUT(N__21298),
            .PACKAGEPIN(V33A_ENn));
    defparam ipInertedIOPad_V33A_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33A_ENn_preio (
            .PADOEN(N__21300),
            .PADOUT(N__21299),
            .PADIN(N__21298),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V1P8A_EN_iopad (
            .OE(N__21291),
            .DIN(N__21290),
            .DOUT(N__21289),
            .PACKAGEPIN(V1P8A_EN));
    defparam ipInertedIOPad_V1P8A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V1P8A_EN_preio (
            .PADOEN(N__21291),
            .PADOUT(N__21290),
            .PADIN(N__21289),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17852),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDDQ_EN_iopad (
            .OE(N__21282),
            .DIN(N__21281),
            .DOUT(N__21280),
            .PACKAGEPIN(VDDQ_EN));
    defparam ipInertedIOPad_VDDQ_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDDQ_EN_preio (
            .PADOEN(N__21282),
            .PADOUT(N__21281),
            .PADIN(N__21280),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__11063),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad (
            .OE(N__21273),
            .DIN(N__21272),
            .DOUT(N__21271),
            .PACKAGEPIN(VCCST_OVERRIDE_3V3));
    defparam ipInertedIOPad_VCCST_OVERRIDE_3V3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_OVERRIDE_3V3_preio (
            .PADOEN(N__21273),
            .PADOUT(N__21272),
            .PADIN(N__21271),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_OK_iopad (
            .OE(N__21264),
            .DIN(N__21263),
            .DOUT(N__21262),
            .PACKAGEPIN(V5S_OK));
    defparam ipInertedIOPad_V5S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5S_OK_preio (
            .PADOEN(N__21264),
            .PADOUT(N__21263),
            .PADIN(N__21262),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S3n_iopad (
            .OE(N__21255),
            .DIN(N__21254),
            .DOUT(N__21253),
            .PACKAGEPIN(SLP_S3n));
    defparam ipInertedIOPad_SLP_S3n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S3n_preio (
            .PADOEN(N__21255),
            .PADOUT(N__21254),
            .PADIN(N__21253),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s3n),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S0n_iopad (
            .OE(N__21246),
            .DIN(N__21245),
            .DOUT(N__21244),
            .PACKAGEPIN(SLP_S0n));
    defparam ipInertedIOPad_SLP_S0n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S0n_preio (
            .PADOEN(N__21246),
            .PADOUT(N__21245),
            .PADIN(N__21244),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_ENn_iopad (
            .OE(N__21237),
            .DIN(N__21236),
            .DOUT(N__21235),
            .PACKAGEPIN(V5S_ENn));
    defparam ipInertedIOPad_V5S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5S_ENn_preio (
            .PADOEN(N__21237),
            .PADOUT(N__21236),
            .PADIN(N__21235),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__11573),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V1P8A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V1P8A_OK_iopad (
            .OE(N__21228),
            .DIN(N__21227),
            .DOUT(N__21226),
            .PACKAGEPIN(V1P8A_OK));
    defparam ipInertedIOPad_V1P8A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V1P8A_OK_preio (
            .PADOEN(N__21228),
            .PADOUT(N__21227),
            .PADIN(N__21226),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v1p8a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTNn_iopad (
            .OE(N__21219),
            .DIN(N__21218),
            .DOUT(N__21217),
            .PACKAGEPIN(PWRBTNn));
    defparam ipInertedIOPad_PWRBTNn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PWRBTNn_preio (
            .PADOEN(N__21219),
            .PADOUT(N__21218),
            .PADIN(N__21217),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTN_LED_iopad (
            .OE(N__21210),
            .DIN(N__21209),
            .DOUT(N__21208),
            .PACKAGEPIN(PWRBTN_LED));
    defparam ipInertedIOPad_PWRBTN_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PWRBTN_LED_preio (
            .PADOEN(N__21210),
            .PADOUT(N__21209),
            .PADIN(N__21208),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__9542),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_2_iopad (
            .OE(N__21201),
            .DIN(N__21200),
            .DOUT(N__21199),
            .PACKAGEPIN(GPIO_FPGA_SoC_2));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_2_preio (
            .PADOEN(N__21201),
            .PADOUT(N__21200),
            .PADIN(N__21199),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad (
            .OE(N__21192),
            .DIN(N__21191),
            .DOUT(N__21190),
            .PACKAGEPIN(VCCIN_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__21192),
            .PADOUT(N__21191),
            .PADIN(N__21190),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_SLP_SUSn_iopad.PULLUP=1'b0;
    IO_PAD ipInertedIOPad_SLP_SUSn_iopad (
            .OE(N__21183),
            .DIN(N__21182),
            .DOUT(N__21181),
            .PACKAGEPIN(SLP_SUSn));
    defparam ipInertedIOPad_SLP_SUSn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_SUSn_preio (
            .PADOEN(N__21183),
            .PADOUT(N__21182),
            .PADIN(N__21181),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_susn),
            .DIN1());
    IO_PAD ipInertedIOPad_CPU_C10_GATE_N_iopad (
            .OE(N__21174),
            .DIN(N__21173),
            .DOUT(N__21172),
            .PACKAGEPIN(CPU_C10_GATE_N));
    defparam ipInertedIOPad_CPU_C10_GATE_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_CPU_C10_GATE_N_preio (
            .PADOEN(N__21174),
            .PADOUT(N__21173),
            .PADIN(N__21172),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_EN_iopad (
            .OE(N__21165),
            .DIN(N__21164),
            .DOUT(N__21163),
            .PACKAGEPIN(VCCST_EN));
    defparam ipInertedIOPad_VCCST_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_EN_preio (
            .PADOEN(N__21165),
            .PADOUT(N__21164),
            .PADIN(N__21163),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__15023),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V33DSW_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V33DSW_OK_iopad (
            .OE(N__21156),
            .DIN(N__21155),
            .DOUT(N__21154),
            .PACKAGEPIN(V33DSW_OK));
    defparam ipInertedIOPad_V33DSW_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33DSW_OK_preio (
            .PADOEN(N__21156),
            .PADOUT(N__21155),
            .PADIN(N__21154),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_TPM_GPIO_iopad (
            .OE(N__21147),
            .DIN(N__21146),
            .DOUT(N__21145),
            .PACKAGEPIN(TPM_GPIO));
    defparam ipInertedIOPad_TPM_GPIO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_TPM_GPIO_preio (
            .PADOEN(N__21147),
            .PADOUT(N__21146),
            .PADIN(N__21145),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSWARN_N_iopad (
            .OE(N__21138),
            .DIN(N__21137),
            .DOUT(N__21136),
            .PACKAGEPIN(SUSWARN_N));
    defparam ipInertedIOPad_SUSWARN_N_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SUSWARN_N_preio (
            .PADOEN(N__21138),
            .PADOUT(N__21137),
            .PADIN(N__21136),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16592),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PLTRSTn_iopad (
            .OE(N__21129),
            .DIN(N__21128),
            .DOUT(N__21127),
            .PACKAGEPIN(PLTRSTn));
    defparam ipInertedIOPad_PLTRSTn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PLTRSTn_preio (
            .PADOEN(N__21129),
            .PADOUT(N__21128),
            .PADIN(N__21127),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_4_iopad (
            .OE(N__21120),
            .DIN(N__21119),
            .DOUT(N__21118),
            .PACKAGEPIN(GPIO_FPGA_SoC_4));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_4_preio (
            .PADOEN(N__21120),
            .PADOUT(N__21119),
            .PADIN(N__21118),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_4),
            .DIN1());
    defparam ipInertedIOPad_VR_READY_VCCIN_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VR_READY_VCCIN_iopad (
            .OE(N__21111),
            .DIN(N__21110),
            .DOUT(N__21109),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam ipInertedIOPad_VR_READY_VCCIN_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCIN_preio (
            .PADOEN(N__21111),
            .PADOUT(N__21110),
            .PADIN(N__21109),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccin),
            .DIN1());
    defparam ipInertedIOPad_V5A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V5A_OK_iopad (
            .OE(N__21102),
            .DIN(N__21101),
            .DOUT(N__21100),
            .PACKAGEPIN(V5A_OK));
    defparam ipInertedIOPad_V5A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5A_OK_preio (
            .PADOEN(N__21102),
            .PADOUT(N__21101),
            .PADIN(N__21100),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_RSMRSTn_iopad (
            .OE(N__21093),
            .DIN(N__21092),
            .DOUT(N__21091),
            .PACKAGEPIN(RSMRSTn));
    defparam ipInertedIOPad_RSMRSTn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RSMRSTn_preio (
            .PADOEN(N__21093),
            .PADOUT(N__21092),
            .PADIN(N__21091),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20717),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_OSC_iopad (
            .OE(N__21084),
            .DIN(N__21083),
            .DOUT(N__21082),
            .PACKAGEPIN(FPGA_OSC));
    defparam ipInertedIOPad_FPGA_OSC_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_OSC_preio (
            .PADOEN(N__21084),
            .PADOUT(N__21083),
            .PADIN(N__21082),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(fpga_osc),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_PWRGD_iopad (
            .OE(N__21075),
            .DIN(N__21074),
            .DOUT(N__21073),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam ipInertedIOPad_VCCST_PWRGD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_PWRGD_preio (
            .PADOEN(N__21075),
            .PADOUT(N__21074),
            .PADIN(N__21073),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19285),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SYS_PWROK_iopad (
            .OE(N__21066),
            .DIN(N__21065),
            .DOUT(N__21064),
            .PACKAGEPIN(SYS_PWROK));
    defparam ipInertedIOPad_SYS_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SYS_PWROK_preio (
            .PADOEN(N__21066),
            .PADOUT(N__21065),
            .PADIN(N__21064),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__11033),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO2_iopad (
            .OE(N__21057),
            .DIN(N__21056),
            .DOUT(N__21055),
            .PACKAGEPIN(SPI_FP_IO2));
    defparam ipInertedIOPad_SPI_FP_IO2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO2_preio (
            .PADOEN(N__21057),
            .PADOUT(N__21056),
            .PADIN(N__21055),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE1_FPGA_iopad (
            .OE(N__21048),
            .DIN(N__21047),
            .DOUT(N__21046),
            .PACKAGEPIN(SATAXPCIE1_FPGA));
    defparam ipInertedIOPad_SATAXPCIE1_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE1_FPGA_preio (
            .PADOEN(N__21048),
            .PADOUT(N__21047),
            .PADIN(N__21046),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_1_iopad (
            .OE(N__21039),
            .DIN(N__21038),
            .DOUT(N__21037),
            .PACKAGEPIN(GPIO_FPGA_EXP_1));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_1_preio (
            .PADOEN(N__21039),
            .PADOUT(N__21038),
            .PADIN(N__21037),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad (
            .OE(N__21030),
            .DIN(N__21029),
            .DOUT(N__21028),
            .PACKAGEPIN(VCCINAUX_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__21030),
            .PADOUT(N__21029),
            .PADIN(N__21028),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PE_iopad (
            .OE(N__21021),
            .DIN(N__21020),
            .DOUT(N__21019),
            .PACKAGEPIN(VCCINAUX_VR_PE));
    defparam ipInertedIOPad_VCCINAUX_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PE_preio (
            .PADOEN(N__21021),
            .PADOUT(N__21020),
            .PADIN(N__21019),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_HDA_SDO_ATP_iopad (
            .OE(N__21012),
            .DIN(N__21011),
            .DOUT(N__21010),
            .PACKAGEPIN(HDA_SDO_ATP));
    defparam ipInertedIOPad_HDA_SDO_ATP_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_HDA_SDO_ATP_preio (
            .PADOEN(N__21012),
            .PADOUT(N__21011),
            .PADIN(N__21010),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__11681),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_2_iopad (
            .OE(N__21003),
            .DIN(N__21002),
            .DOUT(N__21001),
            .PACKAGEPIN(GPIO_FPGA_EXP_2));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_2_preio (
            .PADOEN(N__21003),
            .PADOUT(N__21002),
            .PADIN(N__21001),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VPP_EN_iopad (
            .OE(N__20994),
            .DIN(N__20993),
            .DOUT(N__20992),
            .PACKAGEPIN(VPP_EN));
    defparam ipInertedIOPad_VPP_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VPP_EN_preio (
            .PADOEN(N__20994),
            .PADOUT(N__20993),
            .PADIN(N__20992),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__14969),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VDDQ_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VDDQ_OK_iopad (
            .OE(N__20985),
            .DIN(N__20984),
            .DOUT(N__20983),
            .PACKAGEPIN(VDDQ_OK));
    defparam ipInertedIOPad_VDDQ_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDDQ_OK_preio (
            .PADOEN(N__20985),
            .PADOUT(N__20984),
            .PADIN(N__20983),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vddq_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSACK_N_iopad (
            .OE(N__20976),
            .DIN(N__20975),
            .DOUT(N__20974),
            .PACKAGEPIN(SUSACK_N));
    defparam ipInertedIOPad_SUSACK_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSACK_N_preio (
            .PADOEN(N__20976),
            .PADOUT(N__20975),
            .PADIN(N__20974),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S4n_iopad (
            .OE(N__20967),
            .DIN(N__20966),
            .DOUT(N__20965),
            .PACKAGEPIN(SLP_S4n));
    defparam ipInertedIOPad_SLP_S4n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S4n_preio (
            .PADOEN(N__20967),
            .PADOUT(N__20966),
            .PADIN(N__20965),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s4n),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_CPU_OK_iopad (
            .OE(N__20958),
            .DIN(N__20957),
            .DOUT(N__20956),
            .PACKAGEPIN(VCCST_CPU_OK));
    defparam ipInertedIOPad_VCCST_CPU_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_CPU_OK_preio (
            .PADOEN(N__20958),
            .PADOUT(N__20957),
            .PADIN(N__20956),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vccst_cpu_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_EN_iopad (
            .OE(N__20949),
            .DIN(N__20948),
            .DOUT(N__20947),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam ipInertedIOPad_VCCINAUX_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_EN_preio (
            .PADOEN(N__20949),
            .PADOUT(N__20948),
            .PADIN(N__20947),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17783),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_OK_iopad (
            .OE(N__20940),
            .DIN(N__20939),
            .DOUT(N__20938),
            .PACKAGEPIN(V33S_OK));
    defparam ipInertedIOPad_V33S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33S_OK_preio (
            .PADOEN(N__20940),
            .PADOUT(N__20939),
            .PADIN(N__20938),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_ENn_iopad (
            .OE(N__20931),
            .DIN(N__20930),
            .DOUT(N__20929),
            .PACKAGEPIN(V33S_ENn));
    defparam ipInertedIOPad_V33S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33S_ENn_preio (
            .PADOEN(N__20931),
            .PADOUT(N__20930),
            .PADIN(N__20929),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__11569),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_1_iopad (
            .OE(N__20922),
            .DIN(N__20921),
            .DOUT(N__20920),
            .PACKAGEPIN(GPIO_FPGA_SoC_1));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_1_preio (
            .PADOEN(N__20922),
            .PADOUT(N__20921),
            .PADIN(N__20920),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_1),
            .DIN1());
    defparam ipInertedIOPad_DSW_PWROK_iopad.PULLUP=1'b0;
    IO_PAD ipInertedIOPad_DSW_PWROK_iopad (
            .OE(N__20913),
            .DIN(N__20912),
            .DOUT(N__20911),
            .PACKAGEPIN(DSW_PWROK));
    defparam ipInertedIOPad_DSW_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DSW_PWROK_preio (
            .PADOEN(N__20913),
            .PADOUT(N__20912),
            .PADIN(N__20911),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__18374),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5A_EN_iopad (
            .OE(N__20904),
            .DIN(N__20903),
            .DOUT(N__20902),
            .PACKAGEPIN(V5A_EN));
    defparam ipInertedIOPad_V5A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5A_EN_preio (
            .PADOEN(N__20904),
            .PADOUT(N__20903),
            .PADIN(N__20902),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17848),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_3_iopad (
            .OE(N__20895),
            .DIN(N__20894),
            .DOUT(N__20893),
            .PACKAGEPIN(GPIO_FPGA_SoC_3));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_3_preio (
            .PADOEN(N__20895),
            .PADOUT(N__20894),
            .PADIN(N__20893),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad (
            .OE(N__20886),
            .DIN(N__20885),
            .DOUT(N__20884),
            .PACKAGEPIN(VR_PROCHOT_FPGA_OUT_N));
    defparam ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio (
            .PADOEN(N__20886),
            .PADOUT(N__20885),
            .PADIN(N__20884),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VPP_OK_iopad.PULLUP=1'b0;
    IO_PAD ipInertedIOPad_VPP_OK_iopad (
            .OE(N__20877),
            .DIN(N__20876),
            .DOUT(N__20875),
            .PACKAGEPIN(VPP_OK));
    defparam ipInertedIOPad_VPP_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VPP_OK_preio (
            .PADOEN(N__20877),
            .PADOUT(N__20876),
            .PADIN(N__20875),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vpp_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PE_iopad (
            .OE(N__20868),
            .DIN(N__20867),
            .DOUT(N__20866),
            .PACKAGEPIN(VCCIN_VR_PE));
    defparam ipInertedIOPad_VCCIN_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PE_preio (
            .PADOEN(N__20868),
            .PADOUT(N__20867),
            .PADIN(N__20866),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_EN_iopad (
            .OE(N__20859),
            .DIN(N__20858),
            .DOUT(N__20857),
            .PACKAGEPIN(VCCIN_EN));
    defparam ipInertedIOPad_VCCIN_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_EN_preio (
            .PADOEN(N__20859),
            .PADOUT(N__20858),
            .PADIN(N__20857),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19284),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SOC_SPKR_iopad (
            .OE(N__20850),
            .DIN(N__20849),
            .DOUT(N__20848),
            .PACKAGEPIN(SOC_SPKR));
    defparam ipInertedIOPad_SOC_SPKR_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SOC_SPKR_preio (
            .PADOEN(N__20850),
            .PADOUT(N__20849),
            .PADIN(N__20848),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S5n_iopad (
            .OE(N__20841),
            .DIN(N__20840),
            .DOUT(N__20839),
            .PACKAGEPIN(SLP_S5n));
    defparam ipInertedIOPad_SLP_S5n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S5n_preio (
            .PADOEN(N__20841),
            .PADOUT(N__20840),
            .PADIN(N__20839),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V12_MAIN_MON_iopad (
            .OE(N__20832),
            .DIN(N__20831),
            .DOUT(N__20830),
            .PACKAGEPIN(V12_MAIN_MON));
    defparam ipInertedIOPad_V12_MAIN_MON_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V12_MAIN_MON_preio (
            .PADOEN(N__20832),
            .PADOUT(N__20831),
            .PADIN(N__20830),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO3_iopad (
            .OE(N__20823),
            .DIN(N__20822),
            .DOUT(N__20821),
            .PACKAGEPIN(SPI_FP_IO3));
    defparam ipInertedIOPad_SPI_FP_IO3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO3_preio (
            .PADOEN(N__20823),
            .PADOUT(N__20822),
            .PADIN(N__20821),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE0_FPGA_iopad (
            .OE(N__20814),
            .DIN(N__20813),
            .DOUT(N__20812),
            .PACKAGEPIN(SATAXPCIE0_FPGA));
    defparam ipInertedIOPad_SATAXPCIE0_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE0_FPGA_preio (
            .PADOEN(N__20814),
            .PADOUT(N__20813),
            .PADIN(N__20812),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_OK_iopad (
            .OE(N__20805),
            .DIN(N__20804),
            .DOUT(N__20803),
            .PACKAGEPIN(V33A_OK));
    defparam ipInertedIOPad_V33A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33A_OK_preio (
            .PADOEN(N__20805),
            .PADOUT(N__20804),
            .PADIN(N__20803),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PCH_PWROK_iopad (
            .OE(N__20796),
            .DIN(N__20795),
            .DOUT(N__20794),
            .PACKAGEPIN(PCH_PWROK));
    defparam ipInertedIOPad_PCH_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PCH_PWROK_preio (
            .PADOEN(N__20796),
            .PADOUT(N__20795),
            .PADIN(N__20794),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__11025),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_SLP_WLAN_N_iopad (
            .OE(N__20787),
            .DIN(N__20786),
            .DOUT(N__20785),
            .PACKAGEPIN(FPGA_SLP_WLAN_N));
    defparam ipInertedIOPad_FPGA_SLP_WLAN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_SLP_WLAN_N_preio (
            .PADOEN(N__20787),
            .PADOUT(N__20786),
            .PADIN(N__20785),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    InMux I__4744 (
            .O(N__20768),
            .I(N__20765));
    LocalMux I__4743 (
            .O(N__20765),
            .I(N__20761));
    InMux I__4742 (
            .O(N__20764),
            .I(N__20758));
    Span4Mux_s2_h I__4741 (
            .O(N__20761),
            .I(N__20755));
    LocalMux I__4740 (
            .O(N__20758),
            .I(N__20752));
    Odrv4 I__4739 (
            .O(N__20755),
            .I(\RSMRST_PWRGD.N_240 ));
    Odrv12 I__4738 (
            .O(N__20752),
            .I(\RSMRST_PWRGD.N_240 ));
    InMux I__4737 (
            .O(N__20747),
            .I(N__20740));
    InMux I__4736 (
            .O(N__20746),
            .I(N__20737));
    InMux I__4735 (
            .O(N__20745),
            .I(N__20734));
    InMux I__4734 (
            .O(N__20744),
            .I(N__20729));
    InMux I__4733 (
            .O(N__20743),
            .I(N__20729));
    LocalMux I__4732 (
            .O(N__20740),
            .I(N__20724));
    LocalMux I__4731 (
            .O(N__20737),
            .I(N__20724));
    LocalMux I__4730 (
            .O(N__20734),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__4729 (
            .O(N__20729),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    Odrv4 I__4728 (
            .O(N__20724),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    IoInMux I__4727 (
            .O(N__20717),
            .I(N__20712));
    InMux I__4726 (
            .O(N__20716),
            .I(N__20709));
    InMux I__4725 (
            .O(N__20715),
            .I(N__20705));
    LocalMux I__4724 (
            .O(N__20712),
            .I(N__20699));
    LocalMux I__4723 (
            .O(N__20709),
            .I(N__20696));
    InMux I__4722 (
            .O(N__20708),
            .I(N__20693));
    LocalMux I__4721 (
            .O(N__20705),
            .I(N__20690));
    InMux I__4720 (
            .O(N__20704),
            .I(N__20687));
    InMux I__4719 (
            .O(N__20703),
            .I(N__20684));
    InMux I__4718 (
            .O(N__20702),
            .I(N__20681));
    IoSpan4Mux I__4717 (
            .O(N__20699),
            .I(N__20678));
    Span4Mux_h I__4716 (
            .O(N__20696),
            .I(N__20675));
    LocalMux I__4715 (
            .O(N__20693),
            .I(N__20672));
    Span4Mux_v I__4714 (
            .O(N__20690),
            .I(N__20663));
    LocalMux I__4713 (
            .O(N__20687),
            .I(N__20663));
    LocalMux I__4712 (
            .O(N__20684),
            .I(N__20663));
    LocalMux I__4711 (
            .O(N__20681),
            .I(N__20663));
    IoSpan4Mux I__4710 (
            .O(N__20678),
            .I(N__20660));
    Span4Mux_v I__4709 (
            .O(N__20675),
            .I(N__20657));
    Span12Mux_s10_h I__4708 (
            .O(N__20672),
            .I(N__20654));
    Span4Mux_v I__4707 (
            .O(N__20663),
            .I(N__20651));
    Odrv4 I__4706 (
            .O(N__20660),
            .I(rsmrstn));
    Odrv4 I__4705 (
            .O(N__20657),
            .I(rsmrstn));
    Odrv12 I__4704 (
            .O(N__20654),
            .I(rsmrstn));
    Odrv4 I__4703 (
            .O(N__20651),
            .I(rsmrstn));
    ClkMux I__4702 (
            .O(N__20642),
            .I(N__20638));
    ClkMux I__4701 (
            .O(N__20641),
            .I(N__20632));
    LocalMux I__4700 (
            .O(N__20638),
            .I(N__20625));
    ClkMux I__4699 (
            .O(N__20637),
            .I(N__20622));
    ClkMux I__4698 (
            .O(N__20636),
            .I(N__20619));
    ClkMux I__4697 (
            .O(N__20635),
            .I(N__20616));
    LocalMux I__4696 (
            .O(N__20632),
            .I(N__20612));
    ClkMux I__4695 (
            .O(N__20631),
            .I(N__20609));
    ClkMux I__4694 (
            .O(N__20630),
            .I(N__20606));
    ClkMux I__4693 (
            .O(N__20629),
            .I(N__20601));
    ClkMux I__4692 (
            .O(N__20628),
            .I(N__20597));
    Span4Mux_s3_v I__4691 (
            .O(N__20625),
            .I(N__20586));
    LocalMux I__4690 (
            .O(N__20622),
            .I(N__20586));
    LocalMux I__4689 (
            .O(N__20619),
            .I(N__20586));
    LocalMux I__4688 (
            .O(N__20616),
            .I(N__20582));
    ClkMux I__4687 (
            .O(N__20615),
            .I(N__20579));
    Span4Mux_s3_v I__4686 (
            .O(N__20612),
            .I(N__20574));
    LocalMux I__4685 (
            .O(N__20609),
            .I(N__20574));
    LocalMux I__4684 (
            .O(N__20606),
            .I(N__20571));
    ClkMux I__4683 (
            .O(N__20605),
            .I(N__20568));
    ClkMux I__4682 (
            .O(N__20604),
            .I(N__20565));
    LocalMux I__4681 (
            .O(N__20601),
            .I(N__20561));
    ClkMux I__4680 (
            .O(N__20600),
            .I(N__20554));
    LocalMux I__4679 (
            .O(N__20597),
            .I(N__20551));
    ClkMux I__4678 (
            .O(N__20596),
            .I(N__20548));
    ClkMux I__4677 (
            .O(N__20595),
            .I(N__20544));
    ClkMux I__4676 (
            .O(N__20594),
            .I(N__20539));
    ClkMux I__4675 (
            .O(N__20593),
            .I(N__20535));
    Span4Mux_v I__4674 (
            .O(N__20586),
            .I(N__20529));
    ClkMux I__4673 (
            .O(N__20585),
            .I(N__20526));
    Span4Mux_s3_v I__4672 (
            .O(N__20582),
            .I(N__20521));
    LocalMux I__4671 (
            .O(N__20579),
            .I(N__20521));
    Span4Mux_v I__4670 (
            .O(N__20574),
            .I(N__20518));
    Span4Mux_s3_v I__4669 (
            .O(N__20571),
            .I(N__20511));
    LocalMux I__4668 (
            .O(N__20568),
            .I(N__20511));
    LocalMux I__4667 (
            .O(N__20565),
            .I(N__20511));
    ClkMux I__4666 (
            .O(N__20564),
            .I(N__20508));
    Span4Mux_v I__4665 (
            .O(N__20561),
            .I(N__20505));
    ClkMux I__4664 (
            .O(N__20560),
            .I(N__20502));
    ClkMux I__4663 (
            .O(N__20559),
            .I(N__20499));
    ClkMux I__4662 (
            .O(N__20558),
            .I(N__20496));
    ClkMux I__4661 (
            .O(N__20557),
            .I(N__20492));
    LocalMux I__4660 (
            .O(N__20554),
            .I(N__20488));
    Span4Mux_s2_h I__4659 (
            .O(N__20551),
            .I(N__20483));
    LocalMux I__4658 (
            .O(N__20548),
            .I(N__20483));
    ClkMux I__4657 (
            .O(N__20547),
            .I(N__20480));
    LocalMux I__4656 (
            .O(N__20544),
            .I(N__20477));
    ClkMux I__4655 (
            .O(N__20543),
            .I(N__20474));
    ClkMux I__4654 (
            .O(N__20542),
            .I(N__20468));
    LocalMux I__4653 (
            .O(N__20539),
            .I(N__20462));
    ClkMux I__4652 (
            .O(N__20538),
            .I(N__20459));
    LocalMux I__4651 (
            .O(N__20535),
            .I(N__20455));
    ClkMux I__4650 (
            .O(N__20534),
            .I(N__20452));
    ClkMux I__4649 (
            .O(N__20533),
            .I(N__20447));
    ClkMux I__4648 (
            .O(N__20532),
            .I(N__20444));
    Span4Mux_h I__4647 (
            .O(N__20529),
            .I(N__20438));
    LocalMux I__4646 (
            .O(N__20526),
            .I(N__20438));
    Span4Mux_v I__4645 (
            .O(N__20521),
            .I(N__20429));
    Span4Mux_h I__4644 (
            .O(N__20518),
            .I(N__20429));
    Span4Mux_v I__4643 (
            .O(N__20511),
            .I(N__20429));
    LocalMux I__4642 (
            .O(N__20508),
            .I(N__20429));
    Span4Mux_v I__4641 (
            .O(N__20505),
            .I(N__20423));
    LocalMux I__4640 (
            .O(N__20502),
            .I(N__20423));
    LocalMux I__4639 (
            .O(N__20499),
            .I(N__20418));
    LocalMux I__4638 (
            .O(N__20496),
            .I(N__20418));
    ClkMux I__4637 (
            .O(N__20495),
            .I(N__20415));
    LocalMux I__4636 (
            .O(N__20492),
            .I(N__20412));
    ClkMux I__4635 (
            .O(N__20491),
            .I(N__20409));
    Span4Mux_h I__4634 (
            .O(N__20488),
            .I(N__20404));
    Span4Mux_h I__4633 (
            .O(N__20483),
            .I(N__20399));
    LocalMux I__4632 (
            .O(N__20480),
            .I(N__20399));
    Span4Mux_v I__4631 (
            .O(N__20477),
            .I(N__20394));
    LocalMux I__4630 (
            .O(N__20474),
            .I(N__20394));
    ClkMux I__4629 (
            .O(N__20473),
            .I(N__20391));
    ClkMux I__4628 (
            .O(N__20472),
            .I(N__20388));
    ClkMux I__4627 (
            .O(N__20471),
            .I(N__20385));
    LocalMux I__4626 (
            .O(N__20468),
            .I(N__20381));
    ClkMux I__4625 (
            .O(N__20467),
            .I(N__20378));
    ClkMux I__4624 (
            .O(N__20466),
            .I(N__20374));
    ClkMux I__4623 (
            .O(N__20465),
            .I(N__20371));
    Span4Mux_v I__4622 (
            .O(N__20462),
            .I(N__20365));
    LocalMux I__4621 (
            .O(N__20459),
            .I(N__20365));
    ClkMux I__4620 (
            .O(N__20458),
            .I(N__20362));
    Span4Mux_s3_v I__4619 (
            .O(N__20455),
            .I(N__20357));
    LocalMux I__4618 (
            .O(N__20452),
            .I(N__20357));
    ClkMux I__4617 (
            .O(N__20451),
            .I(N__20354));
    ClkMux I__4616 (
            .O(N__20450),
            .I(N__20351));
    LocalMux I__4615 (
            .O(N__20447),
            .I(N__20348));
    LocalMux I__4614 (
            .O(N__20444),
            .I(N__20345));
    ClkMux I__4613 (
            .O(N__20443),
            .I(N__20342));
    Span4Mux_v I__4612 (
            .O(N__20438),
            .I(N__20336));
    Span4Mux_v I__4611 (
            .O(N__20429),
            .I(N__20336));
    ClkMux I__4610 (
            .O(N__20428),
            .I(N__20333));
    Span4Mux_v I__4609 (
            .O(N__20423),
            .I(N__20330));
    Span4Mux_v I__4608 (
            .O(N__20418),
            .I(N__20325));
    LocalMux I__4607 (
            .O(N__20415),
            .I(N__20325));
    Span4Mux_h I__4606 (
            .O(N__20412),
            .I(N__20320));
    LocalMux I__4605 (
            .O(N__20409),
            .I(N__20320));
    ClkMux I__4604 (
            .O(N__20408),
            .I(N__20317));
    ClkMux I__4603 (
            .O(N__20407),
            .I(N__20314));
    Span4Mux_v I__4602 (
            .O(N__20404),
            .I(N__20305));
    Span4Mux_v I__4601 (
            .O(N__20399),
            .I(N__20305));
    Span4Mux_h I__4600 (
            .O(N__20394),
            .I(N__20305));
    LocalMux I__4599 (
            .O(N__20391),
            .I(N__20305));
    LocalMux I__4598 (
            .O(N__20388),
            .I(N__20302));
    LocalMux I__4597 (
            .O(N__20385),
            .I(N__20299));
    ClkMux I__4596 (
            .O(N__20384),
            .I(N__20296));
    Span4Mux_v I__4595 (
            .O(N__20381),
            .I(N__20291));
    LocalMux I__4594 (
            .O(N__20378),
            .I(N__20291));
    ClkMux I__4593 (
            .O(N__20377),
            .I(N__20288));
    LocalMux I__4592 (
            .O(N__20374),
            .I(N__20285));
    LocalMux I__4591 (
            .O(N__20371),
            .I(N__20282));
    ClkMux I__4590 (
            .O(N__20370),
            .I(N__20279));
    Span4Mux_v I__4589 (
            .O(N__20365),
            .I(N__20274));
    LocalMux I__4588 (
            .O(N__20362),
            .I(N__20274));
    Span4Mux_v I__4587 (
            .O(N__20357),
            .I(N__20265));
    LocalMux I__4586 (
            .O(N__20354),
            .I(N__20265));
    LocalMux I__4585 (
            .O(N__20351),
            .I(N__20265));
    Span4Mux_h I__4584 (
            .O(N__20348),
            .I(N__20265));
    Span4Mux_v I__4583 (
            .O(N__20345),
            .I(N__20260));
    LocalMux I__4582 (
            .O(N__20342),
            .I(N__20260));
    ClkMux I__4581 (
            .O(N__20341),
            .I(N__20257));
    Span4Mux_v I__4580 (
            .O(N__20336),
            .I(N__20254));
    LocalMux I__4579 (
            .O(N__20333),
            .I(N__20251));
    IoSpan4Mux I__4578 (
            .O(N__20330),
            .I(N__20248));
    Span4Mux_v I__4577 (
            .O(N__20325),
            .I(N__20241));
    Span4Mux_v I__4576 (
            .O(N__20320),
            .I(N__20241));
    LocalMux I__4575 (
            .O(N__20317),
            .I(N__20241));
    LocalMux I__4574 (
            .O(N__20314),
            .I(N__20238));
    Span4Mux_v I__4573 (
            .O(N__20305),
            .I(N__20233));
    Span4Mux_h I__4572 (
            .O(N__20302),
            .I(N__20233));
    Span4Mux_h I__4571 (
            .O(N__20299),
            .I(N__20228));
    LocalMux I__4570 (
            .O(N__20296),
            .I(N__20228));
    Span4Mux_h I__4569 (
            .O(N__20291),
            .I(N__20223));
    LocalMux I__4568 (
            .O(N__20288),
            .I(N__20223));
    Span4Mux_s2_h I__4567 (
            .O(N__20285),
            .I(N__20216));
    Span4Mux_h I__4566 (
            .O(N__20282),
            .I(N__20216));
    LocalMux I__4565 (
            .O(N__20279),
            .I(N__20216));
    Span4Mux_h I__4564 (
            .O(N__20274),
            .I(N__20207));
    Span4Mux_v I__4563 (
            .O(N__20265),
            .I(N__20207));
    Span4Mux_h I__4562 (
            .O(N__20260),
            .I(N__20207));
    LocalMux I__4561 (
            .O(N__20257),
            .I(N__20207));
    IoSpan4Mux I__4560 (
            .O(N__20254),
            .I(N__20202));
    Span4Mux_h I__4559 (
            .O(N__20251),
            .I(N__20199));
    IoSpan4Mux I__4558 (
            .O(N__20248),
            .I(N__20192));
    IoSpan4Mux I__4557 (
            .O(N__20241),
            .I(N__20192));
    IoSpan4Mux I__4556 (
            .O(N__20238),
            .I(N__20192));
    Span4Mux_v I__4555 (
            .O(N__20233),
            .I(N__20183));
    Span4Mux_v I__4554 (
            .O(N__20228),
            .I(N__20183));
    Span4Mux_h I__4553 (
            .O(N__20223),
            .I(N__20183));
    Span4Mux_h I__4552 (
            .O(N__20216),
            .I(N__20183));
    Sp12to4 I__4551 (
            .O(N__20207),
            .I(N__20180));
    ClkMux I__4550 (
            .O(N__20206),
            .I(N__20177));
    ClkMux I__4549 (
            .O(N__20205),
            .I(N__20174));
    Odrv4 I__4548 (
            .O(N__20202),
            .I(fpga_osc));
    Odrv4 I__4547 (
            .O(N__20199),
            .I(fpga_osc));
    Odrv4 I__4546 (
            .O(N__20192),
            .I(fpga_osc));
    Odrv4 I__4545 (
            .O(N__20183),
            .I(fpga_osc));
    Odrv12 I__4544 (
            .O(N__20180),
            .I(fpga_osc));
    LocalMux I__4543 (
            .O(N__20177),
            .I(fpga_osc));
    LocalMux I__4542 (
            .O(N__20174),
            .I(fpga_osc));
    InMux I__4541 (
            .O(N__20159),
            .I(N__20047));
    InMux I__4540 (
            .O(N__20158),
            .I(N__20047));
    InMux I__4539 (
            .O(N__20157),
            .I(N__20047));
    InMux I__4538 (
            .O(N__20156),
            .I(N__20047));
    InMux I__4537 (
            .O(N__20155),
            .I(N__20040));
    InMux I__4536 (
            .O(N__20154),
            .I(N__20040));
    InMux I__4535 (
            .O(N__20153),
            .I(N__20040));
    InMux I__4534 (
            .O(N__20152),
            .I(N__20033));
    InMux I__4533 (
            .O(N__20151),
            .I(N__20033));
    InMux I__4532 (
            .O(N__20150),
            .I(N__20033));
    InMux I__4531 (
            .O(N__20149),
            .I(N__20024));
    InMux I__4530 (
            .O(N__20148),
            .I(N__20024));
    InMux I__4529 (
            .O(N__20147),
            .I(N__20024));
    InMux I__4528 (
            .O(N__20146),
            .I(N__20024));
    InMux I__4527 (
            .O(N__20145),
            .I(N__20015));
    InMux I__4526 (
            .O(N__20144),
            .I(N__20015));
    InMux I__4525 (
            .O(N__20143),
            .I(N__20015));
    InMux I__4524 (
            .O(N__20142),
            .I(N__20015));
    InMux I__4523 (
            .O(N__20141),
            .I(N__20008));
    InMux I__4522 (
            .O(N__20140),
            .I(N__20008));
    InMux I__4521 (
            .O(N__20139),
            .I(N__20008));
    InMux I__4520 (
            .O(N__20138),
            .I(N__20001));
    InMux I__4519 (
            .O(N__20137),
            .I(N__20001));
    InMux I__4518 (
            .O(N__20136),
            .I(N__20001));
    InMux I__4517 (
            .O(N__20135),
            .I(N__19992));
    InMux I__4516 (
            .O(N__20134),
            .I(N__19992));
    InMux I__4515 (
            .O(N__20133),
            .I(N__19992));
    InMux I__4514 (
            .O(N__20132),
            .I(N__19992));
    InMux I__4513 (
            .O(N__20131),
            .I(N__19983));
    InMux I__4512 (
            .O(N__20130),
            .I(N__19983));
    InMux I__4511 (
            .O(N__20129),
            .I(N__19983));
    InMux I__4510 (
            .O(N__20128),
            .I(N__19983));
    InMux I__4509 (
            .O(N__20127),
            .I(N__19974));
    InMux I__4508 (
            .O(N__20126),
            .I(N__19974));
    InMux I__4507 (
            .O(N__20125),
            .I(N__19974));
    InMux I__4506 (
            .O(N__20124),
            .I(N__19974));
    InMux I__4505 (
            .O(N__20123),
            .I(N__19969));
    InMux I__4504 (
            .O(N__20122),
            .I(N__19969));
    InMux I__4503 (
            .O(N__20121),
            .I(N__19960));
    InMux I__4502 (
            .O(N__20120),
            .I(N__19960));
    InMux I__4501 (
            .O(N__20119),
            .I(N__19960));
    InMux I__4500 (
            .O(N__20118),
            .I(N__19960));
    InMux I__4499 (
            .O(N__20117),
            .I(N__19951));
    InMux I__4498 (
            .O(N__20116),
            .I(N__19951));
    InMux I__4497 (
            .O(N__20115),
            .I(N__19951));
    InMux I__4496 (
            .O(N__20114),
            .I(N__19951));
    InMux I__4495 (
            .O(N__20113),
            .I(N__19942));
    InMux I__4494 (
            .O(N__20112),
            .I(N__19942));
    InMux I__4493 (
            .O(N__20111),
            .I(N__19942));
    InMux I__4492 (
            .O(N__20110),
            .I(N__19942));
    InMux I__4491 (
            .O(N__20109),
            .I(N__19935));
    InMux I__4490 (
            .O(N__20108),
            .I(N__19935));
    InMux I__4489 (
            .O(N__20107),
            .I(N__19935));
    InMux I__4488 (
            .O(N__20106),
            .I(N__19926));
    InMux I__4487 (
            .O(N__20105),
            .I(N__19926));
    InMux I__4486 (
            .O(N__20104),
            .I(N__19926));
    InMux I__4485 (
            .O(N__20103),
            .I(N__19926));
    InMux I__4484 (
            .O(N__20102),
            .I(N__19919));
    InMux I__4483 (
            .O(N__20101),
            .I(N__19919));
    InMux I__4482 (
            .O(N__20100),
            .I(N__19919));
    InMux I__4481 (
            .O(N__20099),
            .I(N__19910));
    InMux I__4480 (
            .O(N__20098),
            .I(N__19910));
    InMux I__4479 (
            .O(N__20097),
            .I(N__19910));
    InMux I__4478 (
            .O(N__20096),
            .I(N__19910));
    InMux I__4477 (
            .O(N__20095),
            .I(N__19901));
    InMux I__4476 (
            .O(N__20094),
            .I(N__19901));
    InMux I__4475 (
            .O(N__20093),
            .I(N__19901));
    InMux I__4474 (
            .O(N__20092),
            .I(N__19901));
    InMux I__4473 (
            .O(N__20091),
            .I(N__19894));
    InMux I__4472 (
            .O(N__20090),
            .I(N__19894));
    InMux I__4471 (
            .O(N__20089),
            .I(N__19894));
    InMux I__4470 (
            .O(N__20088),
            .I(N__19885));
    InMux I__4469 (
            .O(N__20087),
            .I(N__19885));
    InMux I__4468 (
            .O(N__20086),
            .I(N__19885));
    InMux I__4467 (
            .O(N__20085),
            .I(N__19885));
    InMux I__4466 (
            .O(N__20084),
            .I(N__19880));
    InMux I__4465 (
            .O(N__20083),
            .I(N__19880));
    InMux I__4464 (
            .O(N__20082),
            .I(N__19871));
    InMux I__4463 (
            .O(N__20081),
            .I(N__19871));
    InMux I__4462 (
            .O(N__20080),
            .I(N__19871));
    InMux I__4461 (
            .O(N__20079),
            .I(N__19871));
    InMux I__4460 (
            .O(N__20078),
            .I(N__19868));
    InMux I__4459 (
            .O(N__20077),
            .I(N__19859));
    InMux I__4458 (
            .O(N__20076),
            .I(N__19859));
    InMux I__4457 (
            .O(N__20075),
            .I(N__19859));
    InMux I__4456 (
            .O(N__20074),
            .I(N__19859));
    InMux I__4455 (
            .O(N__20073),
            .I(N__19852));
    InMux I__4454 (
            .O(N__20072),
            .I(N__19852));
    InMux I__4453 (
            .O(N__20071),
            .I(N__19852));
    InMux I__4452 (
            .O(N__20070),
            .I(N__19843));
    InMux I__4451 (
            .O(N__20069),
            .I(N__19843));
    InMux I__4450 (
            .O(N__20068),
            .I(N__19843));
    InMux I__4449 (
            .O(N__20067),
            .I(N__19843));
    InMux I__4448 (
            .O(N__20066),
            .I(N__19840));
    InMux I__4447 (
            .O(N__20065),
            .I(N__19835));
    InMux I__4446 (
            .O(N__20064),
            .I(N__19835));
    InMux I__4445 (
            .O(N__20063),
            .I(N__19832));
    InMux I__4444 (
            .O(N__20062),
            .I(N__19829));
    InMux I__4443 (
            .O(N__20061),
            .I(N__19826));
    InMux I__4442 (
            .O(N__20060),
            .I(N__19821));
    InMux I__4441 (
            .O(N__20059),
            .I(N__19821));
    InMux I__4440 (
            .O(N__20058),
            .I(N__19816));
    InMux I__4439 (
            .O(N__20057),
            .I(N__19816));
    InMux I__4438 (
            .O(N__20056),
            .I(N__19813));
    LocalMux I__4437 (
            .O(N__20047),
            .I(N__19803));
    LocalMux I__4436 (
            .O(N__20040),
            .I(N__19799));
    LocalMux I__4435 (
            .O(N__20033),
            .I(N__19794));
    LocalMux I__4434 (
            .O(N__20024),
            .I(N__19791));
    LocalMux I__4433 (
            .O(N__20015),
            .I(N__19788));
    LocalMux I__4432 (
            .O(N__20008),
            .I(N__19781));
    LocalMux I__4431 (
            .O(N__20001),
            .I(N__19778));
    LocalMux I__4430 (
            .O(N__19992),
            .I(N__19775));
    LocalMux I__4429 (
            .O(N__19983),
            .I(N__19770));
    LocalMux I__4428 (
            .O(N__19974),
            .I(N__19767));
    LocalMux I__4427 (
            .O(N__19969),
            .I(N__19764));
    LocalMux I__4426 (
            .O(N__19960),
            .I(N__19759));
    LocalMux I__4425 (
            .O(N__19951),
            .I(N__19756));
    LocalMux I__4424 (
            .O(N__19942),
            .I(N__19753));
    LocalMux I__4423 (
            .O(N__19935),
            .I(N__19750));
    LocalMux I__4422 (
            .O(N__19926),
            .I(N__19746));
    LocalMux I__4421 (
            .O(N__19919),
            .I(N__19743));
    LocalMux I__4420 (
            .O(N__19910),
            .I(N__19737));
    LocalMux I__4419 (
            .O(N__19901),
            .I(N__19734));
    LocalMux I__4418 (
            .O(N__19894),
            .I(N__19731));
    LocalMux I__4417 (
            .O(N__19885),
            .I(N__19728));
    LocalMux I__4416 (
            .O(N__19880),
            .I(N__19725));
    LocalMux I__4415 (
            .O(N__19871),
            .I(N__19722));
    LocalMux I__4414 (
            .O(N__19868),
            .I(N__19719));
    LocalMux I__4413 (
            .O(N__19859),
            .I(N__19716));
    LocalMux I__4412 (
            .O(N__19852),
            .I(N__19713));
    LocalMux I__4411 (
            .O(N__19843),
            .I(N__19709));
    LocalMux I__4410 (
            .O(N__19840),
            .I(N__19706));
    LocalMux I__4409 (
            .O(N__19835),
            .I(N__19703));
    LocalMux I__4408 (
            .O(N__19832),
            .I(N__19700));
    LocalMux I__4407 (
            .O(N__19829),
            .I(N__19697));
    LocalMux I__4406 (
            .O(N__19826),
            .I(N__19694));
    LocalMux I__4405 (
            .O(N__19821),
            .I(N__19691));
    LocalMux I__4404 (
            .O(N__19816),
            .I(N__19688));
    LocalMux I__4403 (
            .O(N__19813),
            .I(N__19685));
    CEMux I__4402 (
            .O(N__19812),
            .I(N__19568));
    CEMux I__4401 (
            .O(N__19811),
            .I(N__19568));
    CEMux I__4400 (
            .O(N__19810),
            .I(N__19568));
    CEMux I__4399 (
            .O(N__19809),
            .I(N__19568));
    CEMux I__4398 (
            .O(N__19808),
            .I(N__19568));
    CEMux I__4397 (
            .O(N__19807),
            .I(N__19568));
    CEMux I__4396 (
            .O(N__19806),
            .I(N__19568));
    Glb2LocalMux I__4395 (
            .O(N__19803),
            .I(N__19568));
    CEMux I__4394 (
            .O(N__19802),
            .I(N__19568));
    Glb2LocalMux I__4393 (
            .O(N__19799),
            .I(N__19568));
    CEMux I__4392 (
            .O(N__19798),
            .I(N__19568));
    CEMux I__4391 (
            .O(N__19797),
            .I(N__19568));
    Glb2LocalMux I__4390 (
            .O(N__19794),
            .I(N__19568));
    Glb2LocalMux I__4389 (
            .O(N__19791),
            .I(N__19568));
    Glb2LocalMux I__4388 (
            .O(N__19788),
            .I(N__19568));
    CEMux I__4387 (
            .O(N__19787),
            .I(N__19568));
    CEMux I__4386 (
            .O(N__19786),
            .I(N__19568));
    CEMux I__4385 (
            .O(N__19785),
            .I(N__19568));
    CEMux I__4384 (
            .O(N__19784),
            .I(N__19568));
    Glb2LocalMux I__4383 (
            .O(N__19781),
            .I(N__19568));
    Glb2LocalMux I__4382 (
            .O(N__19778),
            .I(N__19568));
    Glb2LocalMux I__4381 (
            .O(N__19775),
            .I(N__19568));
    CEMux I__4380 (
            .O(N__19774),
            .I(N__19568));
    CEMux I__4379 (
            .O(N__19773),
            .I(N__19568));
    Glb2LocalMux I__4378 (
            .O(N__19770),
            .I(N__19568));
    Glb2LocalMux I__4377 (
            .O(N__19767),
            .I(N__19568));
    Glb2LocalMux I__4376 (
            .O(N__19764),
            .I(N__19568));
    CEMux I__4375 (
            .O(N__19763),
            .I(N__19568));
    CEMux I__4374 (
            .O(N__19762),
            .I(N__19568));
    Glb2LocalMux I__4373 (
            .O(N__19759),
            .I(N__19568));
    Glb2LocalMux I__4372 (
            .O(N__19756),
            .I(N__19568));
    Glb2LocalMux I__4371 (
            .O(N__19753),
            .I(N__19568));
    Glb2LocalMux I__4370 (
            .O(N__19750),
            .I(N__19568));
    CEMux I__4369 (
            .O(N__19749),
            .I(N__19568));
    Glb2LocalMux I__4368 (
            .O(N__19746),
            .I(N__19568));
    Glb2LocalMux I__4367 (
            .O(N__19743),
            .I(N__19568));
    CEMux I__4366 (
            .O(N__19742),
            .I(N__19568));
    CEMux I__4365 (
            .O(N__19741),
            .I(N__19568));
    CEMux I__4364 (
            .O(N__19740),
            .I(N__19568));
    Glb2LocalMux I__4363 (
            .O(N__19737),
            .I(N__19568));
    Glb2LocalMux I__4362 (
            .O(N__19734),
            .I(N__19568));
    Glb2LocalMux I__4361 (
            .O(N__19731),
            .I(N__19568));
    Glb2LocalMux I__4360 (
            .O(N__19728),
            .I(N__19568));
    Glb2LocalMux I__4359 (
            .O(N__19725),
            .I(N__19568));
    Glb2LocalMux I__4358 (
            .O(N__19722),
            .I(N__19568));
    Glb2LocalMux I__4357 (
            .O(N__19719),
            .I(N__19568));
    Glb2LocalMux I__4356 (
            .O(N__19716),
            .I(N__19568));
    Glb2LocalMux I__4355 (
            .O(N__19713),
            .I(N__19568));
    CEMux I__4354 (
            .O(N__19712),
            .I(N__19568));
    Glb2LocalMux I__4353 (
            .O(N__19709),
            .I(N__19568));
    Glb2LocalMux I__4352 (
            .O(N__19706),
            .I(N__19568));
    Glb2LocalMux I__4351 (
            .O(N__19703),
            .I(N__19568));
    Glb2LocalMux I__4350 (
            .O(N__19700),
            .I(N__19568));
    Glb2LocalMux I__4349 (
            .O(N__19697),
            .I(N__19568));
    Glb2LocalMux I__4348 (
            .O(N__19694),
            .I(N__19568));
    Glb2LocalMux I__4347 (
            .O(N__19691),
            .I(N__19568));
    Glb2LocalMux I__4346 (
            .O(N__19688),
            .I(N__19568));
    Glb2LocalMux I__4345 (
            .O(N__19685),
            .I(N__19568));
    GlobalMux I__4344 (
            .O(N__19568),
            .I(N__19565));
    gio2CtrlBuf I__4343 (
            .O(N__19565),
            .I(N_65_g));
    InMux I__4342 (
            .O(N__19562),
            .I(N__19559));
    LocalMux I__4341 (
            .O(N__19559),
            .I(N__19556));
    Span4Mux_v I__4340 (
            .O(N__19556),
            .I(N__19552));
    InMux I__4339 (
            .O(N__19555),
            .I(N__19549));
    Span4Mux_v I__4338 (
            .O(N__19552),
            .I(N__19546));
    LocalMux I__4337 (
            .O(N__19549),
            .I(N__19543));
    Odrv4 I__4336 (
            .O(N__19546),
            .I(vddq_ok));
    Odrv12 I__4335 (
            .O(N__19543),
            .I(vddq_ok));
    InMux I__4334 (
            .O(N__19538),
            .I(N__19535));
    LocalMux I__4333 (
            .O(N__19535),
            .I(v5s_ok));
    InMux I__4332 (
            .O(N__19532),
            .I(N__19529));
    LocalMux I__4331 (
            .O(N__19529),
            .I(N__19526));
    Span4Mux_s3_h I__4330 (
            .O(N__19526),
            .I(N__19520));
    InMux I__4329 (
            .O(N__19525),
            .I(N__19515));
    InMux I__4328 (
            .O(N__19524),
            .I(N__19515));
    InMux I__4327 (
            .O(N__19523),
            .I(N__19512));
    Sp12to4 I__4326 (
            .O(N__19520),
            .I(N__19507));
    LocalMux I__4325 (
            .O(N__19515),
            .I(N__19507));
    LocalMux I__4324 (
            .O(N__19512),
            .I(N__19504));
    Odrv12 I__4323 (
            .O(N__19507),
            .I(rsmrst_pwrgd_signal));
    Odrv4 I__4322 (
            .O(N__19504),
            .I(rsmrst_pwrgd_signal));
    InMux I__4321 (
            .O(N__19499),
            .I(N__19496));
    LocalMux I__4320 (
            .O(N__19496),
            .I(N__19493));
    Span4Mux_v I__4319 (
            .O(N__19493),
            .I(N__19490));
    Odrv4 I__4318 (
            .O(N__19490),
            .I(vccst_cpu_ok));
    CascadeMux I__4317 (
            .O(N__19487),
            .I(\ALL_SYS_PWRGD.m4_0_0_a2_1_cascade_ ));
    InMux I__4316 (
            .O(N__19484),
            .I(N__19481));
    LocalMux I__4315 (
            .O(N__19481),
            .I(N__19478));
    Span12Mux_v I__4314 (
            .O(N__19478),
            .I(N__19475));
    Odrv12 I__4313 (
            .O(N__19475),
            .I(v33s_ok));
    CascadeMux I__4312 (
            .O(N__19472),
            .I(N__19467));
    InMux I__4311 (
            .O(N__19471),
            .I(N__19460));
    InMux I__4310 (
            .O(N__19470),
            .I(N__19460));
    InMux I__4309 (
            .O(N__19467),
            .I(N__19453));
    InMux I__4308 (
            .O(N__19466),
            .I(N__19453));
    InMux I__4307 (
            .O(N__19465),
            .I(N__19453));
    LocalMux I__4306 (
            .O(N__19460),
            .I(\ALL_SYS_PWRGD.N_245 ));
    LocalMux I__4305 (
            .O(N__19453),
            .I(\ALL_SYS_PWRGD.N_245 ));
    InMux I__4304 (
            .O(N__19448),
            .I(bfn_11_6_0_));
    InMux I__4303 (
            .O(N__19445),
            .I(N__19436));
    InMux I__4302 (
            .O(N__19444),
            .I(N__19436));
    InMux I__4301 (
            .O(N__19443),
            .I(N__19436));
    LocalMux I__4300 (
            .O(N__19436),
            .I(N__19427));
    InMux I__4299 (
            .O(N__19435),
            .I(N__19418));
    InMux I__4298 (
            .O(N__19434),
            .I(N__19418));
    InMux I__4297 (
            .O(N__19433),
            .I(N__19418));
    InMux I__4296 (
            .O(N__19432),
            .I(N__19418));
    InMux I__4295 (
            .O(N__19431),
            .I(N__19413));
    InMux I__4294 (
            .O(N__19430),
            .I(N__19413));
    Span4Mux_s1_v I__4293 (
            .O(N__19427),
            .I(N__19410));
    LocalMux I__4292 (
            .O(N__19418),
            .I(N__19407));
    LocalMux I__4291 (
            .O(N__19413),
            .I(N__19404));
    Span4Mux_h I__4290 (
            .O(N__19410),
            .I(N__19401));
    Span4Mux_v I__4289 (
            .O(N__19407),
            .I(N__19398));
    Span4Mux_h I__4288 (
            .O(N__19404),
            .I(N__19395));
    Odrv4 I__4287 (
            .O(N__19401),
            .I(\COUNTER.un4_counter_7_THRU_CO ));
    Odrv4 I__4286 (
            .O(N__19398),
            .I(\COUNTER.un4_counter_7_THRU_CO ));
    Odrv4 I__4285 (
            .O(N__19395),
            .I(\COUNTER.un4_counter_7_THRU_CO ));
    CascadeMux I__4284 (
            .O(N__19388),
            .I(\ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa_cascade_ ));
    InMux I__4283 (
            .O(N__19385),
            .I(N__19381));
    CascadeMux I__4282 (
            .O(N__19384),
            .I(N__19378));
    LocalMux I__4281 (
            .O(N__19381),
            .I(N__19375));
    InMux I__4280 (
            .O(N__19378),
            .I(N__19372));
    Span4Mux_v I__4279 (
            .O(N__19375),
            .I(N__19367));
    LocalMux I__4278 (
            .O(N__19372),
            .I(N__19367));
    Span4Mux_h I__4277 (
            .O(N__19367),
            .I(N__19364));
    Odrv4 I__4276 (
            .O(N__19364),
            .I(\ALL_SYS_PWRGD.un1_curr_state10_0 ));
    CascadeMux I__4275 (
            .O(N__19361),
            .I(N__19357));
    InMux I__4274 (
            .O(N__19360),
            .I(N__19353));
    InMux I__4273 (
            .O(N__19357),
            .I(N__19348));
    InMux I__4272 (
            .O(N__19356),
            .I(N__19348));
    LocalMux I__4271 (
            .O(N__19353),
            .I(N__19343));
    LocalMux I__4270 (
            .O(N__19348),
            .I(N__19343));
    Span4Mux_v I__4269 (
            .O(N__19343),
            .I(N__19340));
    Odrv4 I__4268 (
            .O(N__19340),
            .I(\ALL_SYS_PWRGD.N_1_i ));
    InMux I__4267 (
            .O(N__19337),
            .I(N__19334));
    LocalMux I__4266 (
            .O(N__19334),
            .I(N__19331));
    Odrv4 I__4265 (
            .O(N__19331),
            .I(\ALL_SYS_PWRGD.N_36 ));
    InMux I__4264 (
            .O(N__19328),
            .I(N__19310));
    InMux I__4263 (
            .O(N__19327),
            .I(N__19310));
    InMux I__4262 (
            .O(N__19326),
            .I(N__19310));
    InMux I__4261 (
            .O(N__19325),
            .I(N__19310));
    InMux I__4260 (
            .O(N__19324),
            .I(N__19310));
    InMux I__4259 (
            .O(N__19323),
            .I(N__19310));
    LocalMux I__4258 (
            .O(N__19310),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_0 ));
    InMux I__4257 (
            .O(N__19307),
            .I(N__19289));
    InMux I__4256 (
            .O(N__19306),
            .I(N__19289));
    InMux I__4255 (
            .O(N__19305),
            .I(N__19289));
    InMux I__4254 (
            .O(N__19304),
            .I(N__19289));
    InMux I__4253 (
            .O(N__19303),
            .I(N__19289));
    InMux I__4252 (
            .O(N__19302),
            .I(N__19289));
    LocalMux I__4251 (
            .O(N__19289),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__4250 (
            .O(N__19286),
            .I(N__19280));
    IoInMux I__4249 (
            .O(N__19285),
            .I(N__19277));
    IoInMux I__4248 (
            .O(N__19284),
            .I(N__19274));
    InMux I__4247 (
            .O(N__19283),
            .I(N__19269));
    InMux I__4246 (
            .O(N__19280),
            .I(N__19269));
    LocalMux I__4245 (
            .O(N__19277),
            .I(N__19266));
    LocalMux I__4244 (
            .O(N__19274),
            .I(N__19263));
    LocalMux I__4243 (
            .O(N__19269),
            .I(N__19260));
    Span4Mux_s2_v I__4242 (
            .O(N__19266),
            .I(N__19257));
    Span4Mux_s1_v I__4241 (
            .O(N__19263),
            .I(N__19254));
    Span4Mux_s2_h I__4240 (
            .O(N__19260),
            .I(N__19251));
    Span4Mux_v I__4239 (
            .O(N__19257),
            .I(N__19248));
    Span4Mux_v I__4238 (
            .O(N__19254),
            .I(N__19245));
    Span4Mux_h I__4237 (
            .O(N__19251),
            .I(N__19242));
    Span4Mux_h I__4236 (
            .O(N__19248),
            .I(N__19237));
    Span4Mux_v I__4235 (
            .O(N__19245),
            .I(N__19237));
    Span4Mux_h I__4234 (
            .O(N__19242),
            .I(N__19234));
    Odrv4 I__4233 (
            .O(N__19237),
            .I(vccst_pwrgd));
    Odrv4 I__4232 (
            .O(N__19234),
            .I(vccst_pwrgd));
    InMux I__4231 (
            .O(N__19229),
            .I(N__19223));
    CascadeMux I__4230 (
            .O(N__19228),
            .I(N__19220));
    InMux I__4229 (
            .O(N__19227),
            .I(N__19215));
    InMux I__4228 (
            .O(N__19226),
            .I(N__19215));
    LocalMux I__4227 (
            .O(N__19223),
            .I(N__19212));
    InMux I__4226 (
            .O(N__19220),
            .I(N__19209));
    LocalMux I__4225 (
            .O(N__19215),
            .I(N__19206));
    Span4Mux_h I__4224 (
            .O(N__19212),
            .I(N__19203));
    LocalMux I__4223 (
            .O(N__19209),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    Odrv4 I__4222 (
            .O(N__19206),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    Odrv4 I__4221 (
            .O(N__19203),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    InMux I__4220 (
            .O(N__19196),
            .I(N__19190));
    InMux I__4219 (
            .O(N__19195),
            .I(N__19190));
    LocalMux I__4218 (
            .O(N__19190),
            .I(N__19187));
    Span4Mux_v I__4217 (
            .O(N__19187),
            .I(N__19183));
    InMux I__4216 (
            .O(N__19186),
            .I(N__19180));
    Odrv4 I__4215 (
            .O(N__19183),
            .I(\RSMRST_PWRGD.N_241 ));
    LocalMux I__4214 (
            .O(N__19180),
            .I(\RSMRST_PWRGD.N_241 ));
    InMux I__4213 (
            .O(N__19175),
            .I(N__19172));
    LocalMux I__4212 (
            .O(N__19172),
            .I(N__19169));
    Odrv4 I__4211 (
            .O(N__19169),
            .I(\COUNTER.un4_counter_0_and ));
    InMux I__4210 (
            .O(N__19166),
            .I(N__19163));
    LocalMux I__4209 (
            .O(N__19163),
            .I(N__19160));
    Span4Mux_v I__4208 (
            .O(N__19160),
            .I(N__19157));
    Odrv4 I__4207 (
            .O(N__19157),
            .I(\COUNTER.un4_counter_1_and ));
    InMux I__4206 (
            .O(N__19154),
            .I(N__19151));
    LocalMux I__4205 (
            .O(N__19151),
            .I(N__19148));
    Odrv4 I__4204 (
            .O(N__19148),
            .I(\COUNTER.un4_counter_2_and ));
    InMux I__4203 (
            .O(N__19145),
            .I(N__19142));
    LocalMux I__4202 (
            .O(N__19142),
            .I(N__19139));
    Odrv12 I__4201 (
            .O(N__19139),
            .I(\COUNTER.un4_counter_3_and ));
    InMux I__4200 (
            .O(N__19136),
            .I(N__19133));
    LocalMux I__4199 (
            .O(N__19133),
            .I(N__19130));
    Odrv4 I__4198 (
            .O(N__19130),
            .I(\COUNTER.un4_counter_4_and ));
    InMux I__4197 (
            .O(N__19127),
            .I(N__19124));
    LocalMux I__4196 (
            .O(N__19124),
            .I(N__19121));
    Span4Mux_s2_h I__4195 (
            .O(N__19121),
            .I(N__19118));
    Odrv4 I__4194 (
            .O(N__19118),
            .I(\COUNTER.un4_counter_5_and ));
    InMux I__4193 (
            .O(N__19115),
            .I(N__19112));
    LocalMux I__4192 (
            .O(N__19112),
            .I(N__19109));
    Odrv4 I__4191 (
            .O(N__19109),
            .I(\COUNTER.un4_counter_6_and ));
    InMux I__4190 (
            .O(N__19106),
            .I(N__19103));
    LocalMux I__4189 (
            .O(N__19103),
            .I(N__19100));
    Odrv4 I__4188 (
            .O(N__19100),
            .I(\COUNTER.un4_counter_7_and ));
    InMux I__4187 (
            .O(N__19097),
            .I(N__19093));
    InMux I__4186 (
            .O(N__19096),
            .I(N__19090));
    LocalMux I__4185 (
            .O(N__19093),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    LocalMux I__4184 (
            .O(N__19090),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    CascadeMux I__4183 (
            .O(N__19085),
            .I(N__19081));
    InMux I__4182 (
            .O(N__19084),
            .I(N__19078));
    InMux I__4181 (
            .O(N__19081),
            .I(N__19075));
    LocalMux I__4180 (
            .O(N__19078),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    LocalMux I__4179 (
            .O(N__19075),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    InMux I__4178 (
            .O(N__19070),
            .I(N__19066));
    InMux I__4177 (
            .O(N__19069),
            .I(N__19063));
    LocalMux I__4176 (
            .O(N__19066),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    LocalMux I__4175 (
            .O(N__19063),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    InMux I__4174 (
            .O(N__19058),
            .I(N__19054));
    InMux I__4173 (
            .O(N__19057),
            .I(N__19051));
    LocalMux I__4172 (
            .O(N__19054),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    LocalMux I__4171 (
            .O(N__19051),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    InMux I__4170 (
            .O(N__19046),
            .I(N__19042));
    InMux I__4169 (
            .O(N__19045),
            .I(N__19039));
    LocalMux I__4168 (
            .O(N__19042),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    LocalMux I__4167 (
            .O(N__19039),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    CascadeMux I__4166 (
            .O(N__19034),
            .I(N__19030));
    InMux I__4165 (
            .O(N__19033),
            .I(N__19027));
    InMux I__4164 (
            .O(N__19030),
            .I(N__19024));
    LocalMux I__4163 (
            .O(N__19027),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    LocalMux I__4162 (
            .O(N__19024),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    InMux I__4161 (
            .O(N__19019),
            .I(N__19015));
    InMux I__4160 (
            .O(N__19018),
            .I(N__19012));
    LocalMux I__4159 (
            .O(N__19015),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    LocalMux I__4158 (
            .O(N__19012),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    InMux I__4157 (
            .O(N__19007),
            .I(N__19003));
    InMux I__4156 (
            .O(N__19006),
            .I(N__19000));
    LocalMux I__4155 (
            .O(N__19003),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    LocalMux I__4154 (
            .O(N__19000),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    InMux I__4153 (
            .O(N__18995),
            .I(N__18991));
    InMux I__4152 (
            .O(N__18994),
            .I(N__18988));
    LocalMux I__4151 (
            .O(N__18991),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    LocalMux I__4150 (
            .O(N__18988),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    CascadeMux I__4149 (
            .O(N__18983),
            .I(N__18979));
    InMux I__4148 (
            .O(N__18982),
            .I(N__18976));
    InMux I__4147 (
            .O(N__18979),
            .I(N__18973));
    LocalMux I__4146 (
            .O(N__18976),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    LocalMux I__4145 (
            .O(N__18973),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    InMux I__4144 (
            .O(N__18968),
            .I(N__18964));
    InMux I__4143 (
            .O(N__18967),
            .I(N__18961));
    LocalMux I__4142 (
            .O(N__18964),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    LocalMux I__4141 (
            .O(N__18961),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    InMux I__4140 (
            .O(N__18956),
            .I(N__18952));
    InMux I__4139 (
            .O(N__18955),
            .I(N__18949));
    LocalMux I__4138 (
            .O(N__18952),
            .I(N__18946));
    LocalMux I__4137 (
            .O(N__18949),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    Odrv4 I__4136 (
            .O(N__18946),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    InMux I__4135 (
            .O(N__18941),
            .I(N__18937));
    InMux I__4134 (
            .O(N__18940),
            .I(N__18934));
    LocalMux I__4133 (
            .O(N__18937),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    LocalMux I__4132 (
            .O(N__18934),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    CascadeMux I__4131 (
            .O(N__18929),
            .I(N__18925));
    InMux I__4130 (
            .O(N__18928),
            .I(N__18922));
    InMux I__4129 (
            .O(N__18925),
            .I(N__18919));
    LocalMux I__4128 (
            .O(N__18922),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    LocalMux I__4127 (
            .O(N__18919),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    InMux I__4126 (
            .O(N__18914),
            .I(N__18910));
    InMux I__4125 (
            .O(N__18913),
            .I(N__18907));
    LocalMux I__4124 (
            .O(N__18910),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    LocalMux I__4123 (
            .O(N__18907),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    InMux I__4122 (
            .O(N__18902),
            .I(N__18899));
    LocalMux I__4121 (
            .O(N__18899),
            .I(\VPP_VDDQ.un6_count_11 ));
    InMux I__4120 (
            .O(N__18896),
            .I(N__18893));
    LocalMux I__4119 (
            .O(N__18893),
            .I(\VPP_VDDQ.un6_count_10 ));
    CascadeMux I__4118 (
            .O(N__18890),
            .I(\VPP_VDDQ.un6_count_9_cascade_ ));
    InMux I__4117 (
            .O(N__18887),
            .I(N__18884));
    LocalMux I__4116 (
            .O(N__18884),
            .I(\VPP_VDDQ.un6_count_8 ));
    CascadeMux I__4115 (
            .O(N__18881),
            .I(N__18878));
    InMux I__4114 (
            .O(N__18878),
            .I(N__18874));
    InMux I__4113 (
            .O(N__18877),
            .I(N__18871));
    LocalMux I__4112 (
            .O(N__18874),
            .I(N__18868));
    LocalMux I__4111 (
            .O(N__18871),
            .I(N__18865));
    Odrv4 I__4110 (
            .O(N__18868),
            .I(\VPP_VDDQ.count_esr_RNIRFM64Z0Z_15 ));
    Odrv4 I__4109 (
            .O(N__18865),
            .I(\VPP_VDDQ.count_esr_RNIRFM64Z0Z_15 ));
    InMux I__4108 (
            .O(N__18860),
            .I(N__18856));
    InMux I__4107 (
            .O(N__18859),
            .I(N__18853));
    LocalMux I__4106 (
            .O(N__18856),
            .I(N__18850));
    LocalMux I__4105 (
            .O(N__18853),
            .I(\COUNTER.counterZ0Z_14 ));
    Odrv4 I__4104 (
            .O(N__18850),
            .I(\COUNTER.counterZ0Z_14 ));
    InMux I__4103 (
            .O(N__18845),
            .I(N__18841));
    InMux I__4102 (
            .O(N__18844),
            .I(N__18838));
    LocalMux I__4101 (
            .O(N__18841),
            .I(N__18835));
    LocalMux I__4100 (
            .O(N__18838),
            .I(\COUNTER.counterZ0Z_13 ));
    Odrv4 I__4099 (
            .O(N__18835),
            .I(\COUNTER.counterZ0Z_13 ));
    CascadeMux I__4098 (
            .O(N__18830),
            .I(N__18827));
    InMux I__4097 (
            .O(N__18827),
            .I(N__18823));
    InMux I__4096 (
            .O(N__18826),
            .I(N__18820));
    LocalMux I__4095 (
            .O(N__18823),
            .I(N__18817));
    LocalMux I__4094 (
            .O(N__18820),
            .I(\COUNTER.counterZ0Z_15 ));
    Odrv12 I__4093 (
            .O(N__18817),
            .I(\COUNTER.counterZ0Z_15 ));
    InMux I__4092 (
            .O(N__18812),
            .I(N__18808));
    InMux I__4091 (
            .O(N__18811),
            .I(N__18805));
    LocalMux I__4090 (
            .O(N__18808),
            .I(N__18802));
    LocalMux I__4089 (
            .O(N__18805),
            .I(\COUNTER.counterZ0Z_12 ));
    Odrv4 I__4088 (
            .O(N__18802),
            .I(\COUNTER.counterZ0Z_12 ));
    InMux I__4087 (
            .O(N__18797),
            .I(N__18793));
    InMux I__4086 (
            .O(N__18796),
            .I(N__18790));
    LocalMux I__4085 (
            .O(N__18793),
            .I(N__18787));
    LocalMux I__4084 (
            .O(N__18790),
            .I(\COUNTER.counterZ0Z_18 ));
    Odrv4 I__4083 (
            .O(N__18787),
            .I(\COUNTER.counterZ0Z_18 ));
    InMux I__4082 (
            .O(N__18782),
            .I(N__18778));
    InMux I__4081 (
            .O(N__18781),
            .I(N__18775));
    LocalMux I__4080 (
            .O(N__18778),
            .I(N__18772));
    LocalMux I__4079 (
            .O(N__18775),
            .I(\COUNTER.counterZ0Z_17 ));
    Odrv4 I__4078 (
            .O(N__18772),
            .I(\COUNTER.counterZ0Z_17 ));
    CascadeMux I__4077 (
            .O(N__18767),
            .I(N__18763));
    InMux I__4076 (
            .O(N__18766),
            .I(N__18760));
    InMux I__4075 (
            .O(N__18763),
            .I(N__18757));
    LocalMux I__4074 (
            .O(N__18760),
            .I(N__18752));
    LocalMux I__4073 (
            .O(N__18757),
            .I(N__18752));
    Odrv4 I__4072 (
            .O(N__18752),
            .I(\COUNTER.counterZ0Z_19 ));
    InMux I__4071 (
            .O(N__18749),
            .I(N__18746));
    LocalMux I__4070 (
            .O(N__18746),
            .I(N__18742));
    InMux I__4069 (
            .O(N__18745),
            .I(N__18739));
    Span4Mux_s2_h I__4068 (
            .O(N__18742),
            .I(N__18736));
    LocalMux I__4067 (
            .O(N__18739),
            .I(\COUNTER.counterZ0Z_16 ));
    Odrv4 I__4066 (
            .O(N__18736),
            .I(\COUNTER.counterZ0Z_16 ));
    InMux I__4065 (
            .O(N__18731),
            .I(N__18728));
    LocalMux I__4064 (
            .O(N__18728),
            .I(N__18724));
    InMux I__4063 (
            .O(N__18727),
            .I(N__18721));
    Span4Mux_s2_h I__4062 (
            .O(N__18724),
            .I(N__18718));
    LocalMux I__4061 (
            .O(N__18721),
            .I(\COUNTER.counterZ0Z_10 ));
    Odrv4 I__4060 (
            .O(N__18718),
            .I(\COUNTER.counterZ0Z_10 ));
    InMux I__4059 (
            .O(N__18713),
            .I(N__18710));
    LocalMux I__4058 (
            .O(N__18710),
            .I(N__18706));
    InMux I__4057 (
            .O(N__18709),
            .I(N__18703));
    Span4Mux_s2_h I__4056 (
            .O(N__18706),
            .I(N__18700));
    LocalMux I__4055 (
            .O(N__18703),
            .I(\COUNTER.counterZ0Z_9 ));
    Odrv4 I__4054 (
            .O(N__18700),
            .I(\COUNTER.counterZ0Z_9 ));
    CascadeMux I__4053 (
            .O(N__18695),
            .I(N__18692));
    InMux I__4052 (
            .O(N__18692),
            .I(N__18689));
    LocalMux I__4051 (
            .O(N__18689),
            .I(N__18685));
    InMux I__4050 (
            .O(N__18688),
            .I(N__18682));
    Span4Mux_s2_h I__4049 (
            .O(N__18685),
            .I(N__18679));
    LocalMux I__4048 (
            .O(N__18682),
            .I(\COUNTER.counterZ0Z_11 ));
    Odrv4 I__4047 (
            .O(N__18679),
            .I(\COUNTER.counterZ0Z_11 ));
    InMux I__4046 (
            .O(N__18674),
            .I(N__18671));
    LocalMux I__4045 (
            .O(N__18671),
            .I(N__18667));
    InMux I__4044 (
            .O(N__18670),
            .I(N__18664));
    Span4Mux_s2_h I__4043 (
            .O(N__18667),
            .I(N__18661));
    LocalMux I__4042 (
            .O(N__18664),
            .I(\COUNTER.counterZ0Z_8 ));
    Odrv4 I__4041 (
            .O(N__18661),
            .I(\COUNTER.counterZ0Z_8 ));
    InMux I__4040 (
            .O(N__18656),
            .I(N__18653));
    LocalMux I__4039 (
            .O(N__18653),
            .I(\RSMRST_PWRGD.m4_i_i_a2_0_11 ));
    CascadeMux I__4038 (
            .O(N__18650),
            .I(\RSMRST_PWRGD.m4_i_i_a2_0_9_cascade_ ));
    InMux I__4037 (
            .O(N__18647),
            .I(N__18643));
    InMux I__4036 (
            .O(N__18646),
            .I(N__18640));
    LocalMux I__4035 (
            .O(N__18643),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    LocalMux I__4034 (
            .O(N__18640),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    InMux I__4033 (
            .O(N__18635),
            .I(N__18631));
    InMux I__4032 (
            .O(N__18634),
            .I(N__18628));
    LocalMux I__4031 (
            .O(N__18631),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    LocalMux I__4030 (
            .O(N__18628),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    InMux I__4029 (
            .O(N__18623),
            .I(N__18619));
    InMux I__4028 (
            .O(N__18622),
            .I(N__18616));
    LocalMux I__4027 (
            .O(N__18619),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    LocalMux I__4026 (
            .O(N__18616),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    CascadeMux I__4025 (
            .O(N__18611),
            .I(\RSMRST_PWRGD.m4_i_i_a2_0_7_cascade_ ));
    InMux I__4024 (
            .O(N__18608),
            .I(N__18604));
    InMux I__4023 (
            .O(N__18607),
            .I(N__18601));
    LocalMux I__4022 (
            .O(N__18604),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    LocalMux I__4021 (
            .O(N__18601),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    InMux I__4020 (
            .O(N__18596),
            .I(N__18593));
    LocalMux I__4019 (
            .O(N__18593),
            .I(\RSMRST_PWRGD.m4_i_i_a2_0_12 ));
    InMux I__4018 (
            .O(N__18590),
            .I(N__18586));
    InMux I__4017 (
            .O(N__18589),
            .I(N__18583));
    LocalMux I__4016 (
            .O(N__18586),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    LocalMux I__4015 (
            .O(N__18583),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    InMux I__4014 (
            .O(N__18578),
            .I(N__18574));
    InMux I__4013 (
            .O(N__18577),
            .I(N__18571));
    LocalMux I__4012 (
            .O(N__18574),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    LocalMux I__4011 (
            .O(N__18571),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    CascadeMux I__4010 (
            .O(N__18566),
            .I(N__18562));
    InMux I__4009 (
            .O(N__18565),
            .I(N__18559));
    InMux I__4008 (
            .O(N__18562),
            .I(N__18556));
    LocalMux I__4007 (
            .O(N__18559),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    LocalMux I__4006 (
            .O(N__18556),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    InMux I__4005 (
            .O(N__18551),
            .I(N__18547));
    InMux I__4004 (
            .O(N__18550),
            .I(N__18544));
    LocalMux I__4003 (
            .O(N__18547),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    LocalMux I__4002 (
            .O(N__18544),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    InMux I__4001 (
            .O(N__18539),
            .I(N__18536));
    LocalMux I__4000 (
            .O(N__18536),
            .I(\RSMRST_PWRGD.m4_i_i_a2_0_10 ));
    CascadeMux I__3999 (
            .O(N__18533),
            .I(\RSMRST_PWRGD.N_240_cascade_ ));
    SRMux I__3998 (
            .O(N__18530),
            .I(N__18526));
    SRMux I__3997 (
            .O(N__18529),
            .I(N__18523));
    LocalMux I__3996 (
            .O(N__18526),
            .I(N__18519));
    LocalMux I__3995 (
            .O(N__18523),
            .I(N__18516));
    SRMux I__3994 (
            .O(N__18522),
            .I(N__18513));
    Span4Mux_v I__3993 (
            .O(N__18519),
            .I(N__18506));
    Span4Mux_v I__3992 (
            .O(N__18516),
            .I(N__18506));
    LocalMux I__3991 (
            .O(N__18513),
            .I(N__18506));
    Sp12to4 I__3990 (
            .O(N__18506),
            .I(N__18503));
    Odrv12 I__3989 (
            .O(N__18503),
            .I(\RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0 ));
    CascadeMux I__3988 (
            .O(N__18500),
            .I(\RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0_cascade_ ));
    CEMux I__3987 (
            .O(N__18497),
            .I(N__18494));
    LocalMux I__3986 (
            .O(N__18494),
            .I(\RSMRST_PWRGD.N_65_2 ));
    CascadeMux I__3985 (
            .O(N__18491),
            .I(N__18487));
    InMux I__3984 (
            .O(N__18490),
            .I(N__18484));
    InMux I__3983 (
            .O(N__18487),
            .I(N__18481));
    LocalMux I__3982 (
            .O(N__18484),
            .I(N__18476));
    LocalMux I__3981 (
            .O(N__18481),
            .I(N__18476));
    Span4Mux_h I__3980 (
            .O(N__18476),
            .I(N__18473));
    Odrv4 I__3979 (
            .O(N__18473),
            .I(\RSMRST_PWRGD.N_37 ));
    InMux I__3978 (
            .O(N__18470),
            .I(N__18466));
    InMux I__3977 (
            .O(N__18469),
            .I(N__18463));
    LocalMux I__3976 (
            .O(N__18466),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    LocalMux I__3975 (
            .O(N__18463),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    InMux I__3974 (
            .O(N__18458),
            .I(N__18454));
    InMux I__3973 (
            .O(N__18457),
            .I(N__18451));
    LocalMux I__3972 (
            .O(N__18454),
            .I(\POWERLED.count_clkZ0Z_11 ));
    LocalMux I__3971 (
            .O(N__18451),
            .I(\POWERLED.count_clkZ0Z_11 ));
    InMux I__3970 (
            .O(N__18446),
            .I(\POWERLED.un1_count_clk_1_cry_10 ));
    InMux I__3969 (
            .O(N__18443),
            .I(N__18439));
    InMux I__3968 (
            .O(N__18442),
            .I(N__18436));
    LocalMux I__3967 (
            .O(N__18439),
            .I(\POWERLED.count_clkZ0Z_12 ));
    LocalMux I__3966 (
            .O(N__18436),
            .I(\POWERLED.count_clkZ0Z_12 ));
    InMux I__3965 (
            .O(N__18431),
            .I(\POWERLED.un1_count_clk_1_cry_11 ));
    CascadeMux I__3964 (
            .O(N__18428),
            .I(N__18424));
    InMux I__3963 (
            .O(N__18427),
            .I(N__18421));
    InMux I__3962 (
            .O(N__18424),
            .I(N__18418));
    LocalMux I__3961 (
            .O(N__18421),
            .I(\POWERLED.count_clkZ0Z_13 ));
    LocalMux I__3960 (
            .O(N__18418),
            .I(\POWERLED.count_clkZ0Z_13 ));
    InMux I__3959 (
            .O(N__18413),
            .I(\POWERLED.un1_count_clk_1_cry_12 ));
    InMux I__3958 (
            .O(N__18410),
            .I(N__18406));
    InMux I__3957 (
            .O(N__18409),
            .I(N__18403));
    LocalMux I__3956 (
            .O(N__18406),
            .I(\POWERLED.count_clkZ0Z_14 ));
    LocalMux I__3955 (
            .O(N__18403),
            .I(\POWERLED.count_clkZ0Z_14 ));
    InMux I__3954 (
            .O(N__18398),
            .I(\POWERLED.un1_count_clk_1_cry_13 ));
    InMux I__3953 (
            .O(N__18395),
            .I(N__18392));
    LocalMux I__3952 (
            .O(N__18392),
            .I(N__18389));
    Span4Mux_v I__3951 (
            .O(N__18389),
            .I(N__18384));
    InMux I__3950 (
            .O(N__18388),
            .I(N__18381));
    InMux I__3949 (
            .O(N__18387),
            .I(N__18378));
    IoSpan4Mux I__3948 (
            .O(N__18384),
            .I(N__18371));
    LocalMux I__3947 (
            .O(N__18381),
            .I(N__18366));
    LocalMux I__3946 (
            .O(N__18378),
            .I(N__18366));
    InMux I__3945 (
            .O(N__18377),
            .I(N__18363));
    InMux I__3944 (
            .O(N__18376),
            .I(N__18360));
    InMux I__3943 (
            .O(N__18375),
            .I(N__18357));
    IoInMux I__3942 (
            .O(N__18374),
            .I(N__18353));
    Span4Mux_s3_h I__3941 (
            .O(N__18371),
            .I(N__18344));
    Span4Mux_v I__3940 (
            .O(N__18366),
            .I(N__18344));
    LocalMux I__3939 (
            .O(N__18363),
            .I(N__18344));
    LocalMux I__3938 (
            .O(N__18360),
            .I(N__18344));
    LocalMux I__3937 (
            .O(N__18357),
            .I(N__18341));
    InMux I__3936 (
            .O(N__18356),
            .I(N__18338));
    LocalMux I__3935 (
            .O(N__18353),
            .I(N__18333));
    Span4Mux_h I__3934 (
            .O(N__18344),
            .I(N__18328));
    Span4Mux_v I__3933 (
            .O(N__18341),
            .I(N__18328));
    LocalMux I__3932 (
            .O(N__18338),
            .I(N__18325));
    InMux I__3931 (
            .O(N__18337),
            .I(N__18322));
    InMux I__3930 (
            .O(N__18336),
            .I(N__18319));
    Span4Mux_s3_h I__3929 (
            .O(N__18333),
            .I(N__18315));
    Span4Mux_v I__3928 (
            .O(N__18328),
            .I(N__18308));
    Span4Mux_h I__3927 (
            .O(N__18325),
            .I(N__18308));
    LocalMux I__3926 (
            .O(N__18322),
            .I(N__18308));
    LocalMux I__3925 (
            .O(N__18319),
            .I(N__18305));
    CascadeMux I__3924 (
            .O(N__18318),
            .I(N__18302));
    Span4Mux_v I__3923 (
            .O(N__18315),
            .I(N__18294));
    Span4Mux_v I__3922 (
            .O(N__18308),
            .I(N__18294));
    Span4Mux_s2_v I__3921 (
            .O(N__18305),
            .I(N__18294));
    InMux I__3920 (
            .O(N__18302),
            .I(N__18289));
    InMux I__3919 (
            .O(N__18301),
            .I(N__18289));
    Odrv4 I__3918 (
            .O(N__18294),
            .I(CONSTANT_ONE_NET));
    LocalMux I__3917 (
            .O(N__18289),
            .I(CONSTANT_ONE_NET));
    InMux I__3916 (
            .O(N__18284),
            .I(bfn_9_11_0_));
    CascadeMux I__3915 (
            .O(N__18281),
            .I(N__18277));
    InMux I__3914 (
            .O(N__18280),
            .I(N__18274));
    InMux I__3913 (
            .O(N__18277),
            .I(N__18271));
    LocalMux I__3912 (
            .O(N__18274),
            .I(\POWERLED.count_clkZ0Z_15 ));
    LocalMux I__3911 (
            .O(N__18271),
            .I(\POWERLED.count_clkZ0Z_15 ));
    CEMux I__3910 (
            .O(N__18266),
            .I(N__18263));
    LocalMux I__3909 (
            .O(N__18263),
            .I(N__18260));
    Span4Mux_v I__3908 (
            .O(N__18260),
            .I(N__18257));
    Span4Mux_s2_h I__3907 (
            .O(N__18257),
            .I(N__18254));
    Odrv4 I__3906 (
            .O(N__18254),
            .I(\POWERLED.N_65_0 ));
    SRMux I__3905 (
            .O(N__18251),
            .I(N__18247));
    SRMux I__3904 (
            .O(N__18250),
            .I(N__18244));
    LocalMux I__3903 (
            .O(N__18247),
            .I(N__18240));
    LocalMux I__3902 (
            .O(N__18244),
            .I(N__18237));
    SRMux I__3901 (
            .O(N__18243),
            .I(N__18234));
    Span4Mux_v I__3900 (
            .O(N__18240),
            .I(N__18226));
    Span4Mux_v I__3899 (
            .O(N__18237),
            .I(N__18226));
    LocalMux I__3898 (
            .O(N__18234),
            .I(N__18226));
    InMux I__3897 (
            .O(N__18233),
            .I(N__18223));
    Odrv4 I__3896 (
            .O(N__18226),
            .I(\POWERLED.count_clk_RNIOH1J11Z0Z_7 ));
    LocalMux I__3895 (
            .O(N__18223),
            .I(\POWERLED.count_clk_RNIOH1J11Z0Z_7 ));
    InMux I__3894 (
            .O(N__18218),
            .I(N__18214));
    InMux I__3893 (
            .O(N__18217),
            .I(N__18211));
    LocalMux I__3892 (
            .O(N__18214),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    LocalMux I__3891 (
            .O(N__18211),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    InMux I__3890 (
            .O(N__18206),
            .I(N__18202));
    InMux I__3889 (
            .O(N__18205),
            .I(N__18199));
    LocalMux I__3888 (
            .O(N__18202),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    LocalMux I__3887 (
            .O(N__18199),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    CascadeMux I__3886 (
            .O(N__18194),
            .I(N__18190));
    InMux I__3885 (
            .O(N__18193),
            .I(N__18187));
    InMux I__3884 (
            .O(N__18190),
            .I(N__18184));
    LocalMux I__3883 (
            .O(N__18187),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    LocalMux I__3882 (
            .O(N__18184),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    InMux I__3881 (
            .O(N__18179),
            .I(N__18175));
    InMux I__3880 (
            .O(N__18178),
            .I(N__18172));
    LocalMux I__3879 (
            .O(N__18175),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    LocalMux I__3878 (
            .O(N__18172),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    InMux I__3877 (
            .O(N__18167),
            .I(N__18163));
    InMux I__3876 (
            .O(N__18166),
            .I(N__18160));
    LocalMux I__3875 (
            .O(N__18163),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    LocalMux I__3874 (
            .O(N__18160),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    InMux I__3873 (
            .O(N__18155),
            .I(N__18151));
    InMux I__3872 (
            .O(N__18154),
            .I(N__18148));
    LocalMux I__3871 (
            .O(N__18151),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    LocalMux I__3870 (
            .O(N__18148),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    CascadeMux I__3869 (
            .O(N__18143),
            .I(N__18139));
    InMux I__3868 (
            .O(N__18142),
            .I(N__18136));
    InMux I__3867 (
            .O(N__18139),
            .I(N__18133));
    LocalMux I__3866 (
            .O(N__18136),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    LocalMux I__3865 (
            .O(N__18133),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    InMux I__3864 (
            .O(N__18128),
            .I(N__18124));
    InMux I__3863 (
            .O(N__18127),
            .I(N__18121));
    LocalMux I__3862 (
            .O(N__18124),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    LocalMux I__3861 (
            .O(N__18121),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    InMux I__3860 (
            .O(N__18116),
            .I(N__18111));
    InMux I__3859 (
            .O(N__18115),
            .I(N__18106));
    InMux I__3858 (
            .O(N__18114),
            .I(N__18106));
    LocalMux I__3857 (
            .O(N__18111),
            .I(\POWERLED.count_clkZ0Z_3 ));
    LocalMux I__3856 (
            .O(N__18106),
            .I(\POWERLED.count_clkZ0Z_3 ));
    InMux I__3855 (
            .O(N__18101),
            .I(\POWERLED.un1_count_clk_1_cry_2 ));
    InMux I__3854 (
            .O(N__18098),
            .I(N__18093));
    InMux I__3853 (
            .O(N__18097),
            .I(N__18088));
    InMux I__3852 (
            .O(N__18096),
            .I(N__18088));
    LocalMux I__3851 (
            .O(N__18093),
            .I(\POWERLED.count_clkZ0Z_4 ));
    LocalMux I__3850 (
            .O(N__18088),
            .I(\POWERLED.count_clkZ0Z_4 ));
    InMux I__3849 (
            .O(N__18083),
            .I(\POWERLED.un1_count_clk_1_cry_3 ));
    InMux I__3848 (
            .O(N__18080),
            .I(N__18074));
    InMux I__3847 (
            .O(N__18079),
            .I(N__18069));
    InMux I__3846 (
            .O(N__18078),
            .I(N__18069));
    InMux I__3845 (
            .O(N__18077),
            .I(N__18066));
    LocalMux I__3844 (
            .O(N__18074),
            .I(\POWERLED.count_clkZ0Z_5 ));
    LocalMux I__3843 (
            .O(N__18069),
            .I(\POWERLED.count_clkZ0Z_5 ));
    LocalMux I__3842 (
            .O(N__18066),
            .I(\POWERLED.count_clkZ0Z_5 ));
    InMux I__3841 (
            .O(N__18059),
            .I(\POWERLED.un1_count_clk_1_cry_4 ));
    InMux I__3840 (
            .O(N__18056),
            .I(N__18052));
    InMux I__3839 (
            .O(N__18055),
            .I(N__18048));
    LocalMux I__3838 (
            .O(N__18052),
            .I(N__18045));
    InMux I__3837 (
            .O(N__18051),
            .I(N__18041));
    LocalMux I__3836 (
            .O(N__18048),
            .I(N__18038));
    Span4Mux_h I__3835 (
            .O(N__18045),
            .I(N__18035));
    InMux I__3834 (
            .O(N__18044),
            .I(N__18032));
    LocalMux I__3833 (
            .O(N__18041),
            .I(\POWERLED.count_clkZ0Z_6 ));
    Odrv4 I__3832 (
            .O(N__18038),
            .I(\POWERLED.count_clkZ0Z_6 ));
    Odrv4 I__3831 (
            .O(N__18035),
            .I(\POWERLED.count_clkZ0Z_6 ));
    LocalMux I__3830 (
            .O(N__18032),
            .I(\POWERLED.count_clkZ0Z_6 ));
    InMux I__3829 (
            .O(N__18023),
            .I(\POWERLED.un1_count_clk_1_cry_5 ));
    InMux I__3828 (
            .O(N__18020),
            .I(N__18013));
    InMux I__3827 (
            .O(N__18019),
            .I(N__18008));
    InMux I__3826 (
            .O(N__18018),
            .I(N__18008));
    InMux I__3825 (
            .O(N__18017),
            .I(N__18001));
    InMux I__3824 (
            .O(N__18016),
            .I(N__18001));
    LocalMux I__3823 (
            .O(N__18013),
            .I(N__17997));
    LocalMux I__3822 (
            .O(N__18008),
            .I(N__17994));
    InMux I__3821 (
            .O(N__18007),
            .I(N__17991));
    CascadeMux I__3820 (
            .O(N__18006),
            .I(N__17987));
    LocalMux I__3819 (
            .O(N__18001),
            .I(N__17984));
    InMux I__3818 (
            .O(N__18000),
            .I(N__17981));
    Span4Mux_h I__3817 (
            .O(N__17997),
            .I(N__17978));
    Span12Mux_s7_v I__3816 (
            .O(N__17994),
            .I(N__17973));
    LocalMux I__3815 (
            .O(N__17991),
            .I(N__17973));
    InMux I__3814 (
            .O(N__17990),
            .I(N__17968));
    InMux I__3813 (
            .O(N__17987),
            .I(N__17968));
    Span4Mux_h I__3812 (
            .O(N__17984),
            .I(N__17965));
    LocalMux I__3811 (
            .O(N__17981),
            .I(\POWERLED.count_clkZ0Z_7 ));
    Odrv4 I__3810 (
            .O(N__17978),
            .I(\POWERLED.count_clkZ0Z_7 ));
    Odrv12 I__3809 (
            .O(N__17973),
            .I(\POWERLED.count_clkZ0Z_7 ));
    LocalMux I__3808 (
            .O(N__17968),
            .I(\POWERLED.count_clkZ0Z_7 ));
    Odrv4 I__3807 (
            .O(N__17965),
            .I(\POWERLED.count_clkZ0Z_7 ));
    InMux I__3806 (
            .O(N__17954),
            .I(\POWERLED.un1_count_clk_1_cry_6 ));
    InMux I__3805 (
            .O(N__17951),
            .I(N__17946));
    InMux I__3804 (
            .O(N__17950),
            .I(N__17941));
    InMux I__3803 (
            .O(N__17949),
            .I(N__17941));
    LocalMux I__3802 (
            .O(N__17946),
            .I(\POWERLED.count_clkZ0Z_8 ));
    LocalMux I__3801 (
            .O(N__17941),
            .I(\POWERLED.count_clkZ0Z_8 ));
    InMux I__3800 (
            .O(N__17936),
            .I(bfn_9_10_0_));
    InMux I__3799 (
            .O(N__17933),
            .I(N__17927));
    InMux I__3798 (
            .O(N__17932),
            .I(N__17920));
    InMux I__3797 (
            .O(N__17931),
            .I(N__17920));
    InMux I__3796 (
            .O(N__17930),
            .I(N__17920));
    LocalMux I__3795 (
            .O(N__17927),
            .I(\POWERLED.count_clkZ0Z_9 ));
    LocalMux I__3794 (
            .O(N__17920),
            .I(\POWERLED.count_clkZ0Z_9 ));
    InMux I__3793 (
            .O(N__17915),
            .I(\POWERLED.un1_count_clk_1_cry_8 ));
    InMux I__3792 (
            .O(N__17912),
            .I(N__17908));
    InMux I__3791 (
            .O(N__17911),
            .I(N__17905));
    LocalMux I__3790 (
            .O(N__17908),
            .I(\POWERLED.count_clkZ0Z_10 ));
    LocalMux I__3789 (
            .O(N__17905),
            .I(\POWERLED.count_clkZ0Z_10 ));
    InMux I__3788 (
            .O(N__17900),
            .I(\POWERLED.un1_count_clk_1_cry_9 ));
    InMux I__3787 (
            .O(N__17897),
            .I(N__17894));
    LocalMux I__3786 (
            .O(N__17894),
            .I(\ALL_SYS_PWRGD.un4_count_9 ));
    SRMux I__3785 (
            .O(N__17891),
            .I(N__17887));
    SRMux I__3784 (
            .O(N__17890),
            .I(N__17884));
    LocalMux I__3783 (
            .O(N__17887),
            .I(N__17880));
    LocalMux I__3782 (
            .O(N__17884),
            .I(N__17877));
    SRMux I__3781 (
            .O(N__17883),
            .I(N__17874));
    Span4Mux_v I__3780 (
            .O(N__17880),
            .I(N__17867));
    Span4Mux_v I__3779 (
            .O(N__17877),
            .I(N__17867));
    LocalMux I__3778 (
            .O(N__17874),
            .I(N__17867));
    Sp12to4 I__3777 (
            .O(N__17867),
            .I(N__17864));
    Odrv12 I__3776 (
            .O(N__17864),
            .I(\ALL_SYS_PWRGD.curr_state_RNIKNST6Z0Z_0 ));
    CascadeMux I__3775 (
            .O(N__17861),
            .I(\ALL_SYS_PWRGD.curr_state_RNIKNST6Z0Z_0_cascade_ ));
    CEMux I__3774 (
            .O(N__17858),
            .I(N__17855));
    LocalMux I__3773 (
            .O(N__17855),
            .I(\ALL_SYS_PWRGD.N_65_4 ));
    IoInMux I__3772 (
            .O(N__17852),
            .I(N__17849));
    LocalMux I__3771 (
            .O(N__17849),
            .I(N__17845));
    IoInMux I__3770 (
            .O(N__17848),
            .I(N__17842));
    IoSpan4Mux I__3769 (
            .O(N__17845),
            .I(N__17838));
    LocalMux I__3768 (
            .O(N__17842),
            .I(N__17835));
    InMux I__3767 (
            .O(N__17841),
            .I(N__17832));
    IoSpan4Mux I__3766 (
            .O(N__17838),
            .I(N__17829));
    Span12Mux_s8_h I__3765 (
            .O(N__17835),
            .I(N__17824));
    LocalMux I__3764 (
            .O(N__17832),
            .I(N__17824));
    Odrv4 I__3763 (
            .O(N__17829),
            .I(slp_susn));
    Odrv12 I__3762 (
            .O(N__17824),
            .I(slp_susn));
    InMux I__3761 (
            .O(N__17819),
            .I(N__17816));
    LocalMux I__3760 (
            .O(N__17816),
            .I(N__17813));
    Span4Mux_v I__3759 (
            .O(N__17813),
            .I(N__17810));
    Sp12to4 I__3758 (
            .O(N__17810),
            .I(N__17807));
    Odrv12 I__3757 (
            .O(N__17807),
            .I(v5a_ok));
    CascadeMux I__3756 (
            .O(N__17804),
            .I(N__17801));
    InMux I__3755 (
            .O(N__17801),
            .I(N__17798));
    LocalMux I__3754 (
            .O(N__17798),
            .I(N__17795));
    Span4Mux_h I__3753 (
            .O(N__17795),
            .I(N__17792));
    Span4Mux_v I__3752 (
            .O(N__17792),
            .I(N__17789));
    Span4Mux_v I__3751 (
            .O(N__17789),
            .I(N__17786));
    Odrv4 I__3750 (
            .O(N__17786),
            .I(v33a_ok));
    IoInMux I__3749 (
            .O(N__17783),
            .I(N__17780));
    LocalMux I__3748 (
            .O(N__17780),
            .I(N__17777));
    IoSpan4Mux I__3747 (
            .O(N__17777),
            .I(N__17773));
    InMux I__3746 (
            .O(N__17776),
            .I(N__17770));
    IoSpan4Mux I__3745 (
            .O(N__17773),
            .I(N__17767));
    LocalMux I__3744 (
            .O(N__17770),
            .I(N__17764));
    Span4Mux_s3_h I__3743 (
            .O(N__17767),
            .I(N__17761));
    Sp12to4 I__3742 (
            .O(N__17764),
            .I(N__17758));
    Sp12to4 I__3741 (
            .O(N__17761),
            .I(N__17753));
    Span12Mux_s11_v I__3740 (
            .O(N__17758),
            .I(N__17753));
    Odrv12 I__3739 (
            .O(N__17753),
            .I(v1p8a_ok));
    CascadeMux I__3738 (
            .O(N__17750),
            .I(N__17747));
    InMux I__3737 (
            .O(N__17747),
            .I(N__17741));
    InMux I__3736 (
            .O(N__17746),
            .I(N__17741));
    LocalMux I__3735 (
            .O(N__17741),
            .I(\COUNTER.tmp_i ));
    InMux I__3734 (
            .O(N__17738),
            .I(N__17734));
    IoInMux I__3733 (
            .O(N__17737),
            .I(N__17731));
    LocalMux I__3732 (
            .O(N__17734),
            .I(N__17728));
    LocalMux I__3731 (
            .O(N__17731),
            .I(N__17725));
    Span4Mux_v I__3730 (
            .O(N__17728),
            .I(N__17722));
    Span4Mux_s0_h I__3729 (
            .O(N__17725),
            .I(N__17719));
    Span4Mux_h I__3728 (
            .O(N__17722),
            .I(N__17716));
    Span4Mux_h I__3727 (
            .O(N__17719),
            .I(N__17713));
    Span4Mux_v I__3726 (
            .O(N__17716),
            .I(N__17710));
    Span4Mux_h I__3725 (
            .O(N__17713),
            .I(N__17707));
    Odrv4 I__3724 (
            .O(N__17710),
            .I(tmp_RNIRH3P));
    Odrv4 I__3723 (
            .O(N__17707),
            .I(tmp_RNIRH3P));
    CascadeMux I__3722 (
            .O(N__17702),
            .I(N__17698));
    InMux I__3721 (
            .O(N__17701),
            .I(N__17695));
    InMux I__3720 (
            .O(N__17698),
            .I(N__17692));
    LocalMux I__3719 (
            .O(N__17695),
            .I(N__17687));
    LocalMux I__3718 (
            .O(N__17692),
            .I(N__17687));
    Span4Mux_h I__3717 (
            .O(N__17687),
            .I(N__17684));
    Odrv4 I__3716 (
            .O(N__17684),
            .I(\POWERLED.count_clk_1_sqmuxa_5_i ));
    InMux I__3715 (
            .O(N__17681),
            .I(N__17677));
    InMux I__3714 (
            .O(N__17680),
            .I(N__17674));
    LocalMux I__3713 (
            .O(N__17677),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__3712 (
            .O(N__17674),
            .I(\POWERLED.count_clkZ0Z_0 ));
    InMux I__3711 (
            .O(N__17669),
            .I(N__17663));
    InMux I__3710 (
            .O(N__17668),
            .I(N__17656));
    InMux I__3709 (
            .O(N__17667),
            .I(N__17656));
    InMux I__3708 (
            .O(N__17666),
            .I(N__17656));
    LocalMux I__3707 (
            .O(N__17663),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__3706 (
            .O(N__17656),
            .I(\POWERLED.count_clkZ0Z_1 ));
    InMux I__3705 (
            .O(N__17651),
            .I(\POWERLED.un1_count_clk_1_cry_0 ));
    CascadeMux I__3704 (
            .O(N__17648),
            .I(N__17644));
    InMux I__3703 (
            .O(N__17647),
            .I(N__17640));
    InMux I__3702 (
            .O(N__17644),
            .I(N__17637));
    InMux I__3701 (
            .O(N__17643),
            .I(N__17634));
    LocalMux I__3700 (
            .O(N__17640),
            .I(\POWERLED.count_clkZ0Z_2 ));
    LocalMux I__3699 (
            .O(N__17637),
            .I(\POWERLED.count_clkZ0Z_2 ));
    LocalMux I__3698 (
            .O(N__17634),
            .I(\POWERLED.count_clkZ0Z_2 ));
    InMux I__3697 (
            .O(N__17627),
            .I(\POWERLED.un1_count_clk_1_cry_1 ));
    InMux I__3696 (
            .O(N__17624),
            .I(N__17621));
    LocalMux I__3695 (
            .O(N__17621),
            .I(N__17618));
    Span4Mux_v I__3694 (
            .O(N__17618),
            .I(N__17615));
    Odrv4 I__3693 (
            .O(N__17615),
            .I(\COUNTER.counter_1_cry_3_THRU_CO ));
    InMux I__3692 (
            .O(N__17612),
            .I(N__17608));
    CascadeMux I__3691 (
            .O(N__17611),
            .I(N__17604));
    LocalMux I__3690 (
            .O(N__17608),
            .I(N__17601));
    InMux I__3689 (
            .O(N__17607),
            .I(N__17596));
    InMux I__3688 (
            .O(N__17604),
            .I(N__17596));
    Odrv12 I__3687 (
            .O(N__17601),
            .I(\COUNTER.counterZ0Z_4 ));
    LocalMux I__3686 (
            .O(N__17596),
            .I(\COUNTER.counterZ0Z_4 ));
    InMux I__3685 (
            .O(N__17591),
            .I(N__17587));
    CascadeMux I__3684 (
            .O(N__17590),
            .I(N__17584));
    LocalMux I__3683 (
            .O(N__17587),
            .I(N__17581));
    InMux I__3682 (
            .O(N__17584),
            .I(N__17578));
    Sp12to4 I__3681 (
            .O(N__17581),
            .I(N__17571));
    LocalMux I__3680 (
            .O(N__17578),
            .I(N__17571));
    InMux I__3679 (
            .O(N__17577),
            .I(N__17566));
    InMux I__3678 (
            .O(N__17576),
            .I(N__17566));
    Odrv12 I__3677 (
            .O(N__17571),
            .I(\COUNTER.counterZ0Z_0 ));
    LocalMux I__3676 (
            .O(N__17566),
            .I(\COUNTER.counterZ0Z_0 ));
    InMux I__3675 (
            .O(N__17561),
            .I(N__17558));
    LocalMux I__3674 (
            .O(N__17558),
            .I(N__17555));
    Odrv12 I__3673 (
            .O(N__17555),
            .I(\COUNTER.counter_1_cry_1_THRU_CO ));
    InMux I__3672 (
            .O(N__17552),
            .I(N__17549));
    LocalMux I__3671 (
            .O(N__17549),
            .I(N__17546));
    Span4Mux_s1_v I__3670 (
            .O(N__17546),
            .I(N__17541));
    InMux I__3669 (
            .O(N__17545),
            .I(N__17536));
    InMux I__3668 (
            .O(N__17544),
            .I(N__17536));
    Odrv4 I__3667 (
            .O(N__17541),
            .I(\COUNTER.counterZ0Z_2 ));
    LocalMux I__3666 (
            .O(N__17536),
            .I(\COUNTER.counterZ0Z_2 ));
    InMux I__3665 (
            .O(N__17531),
            .I(N__17528));
    LocalMux I__3664 (
            .O(N__17528),
            .I(N__17525));
    Odrv12 I__3663 (
            .O(N__17525),
            .I(\COUNTER.counter_1_cry_2_THRU_CO ));
    InMux I__3662 (
            .O(N__17522),
            .I(N__17518));
    CascadeMux I__3661 (
            .O(N__17521),
            .I(N__17515));
    LocalMux I__3660 (
            .O(N__17518),
            .I(N__17511));
    InMux I__3659 (
            .O(N__17515),
            .I(N__17506));
    InMux I__3658 (
            .O(N__17514),
            .I(N__17506));
    Odrv12 I__3657 (
            .O(N__17511),
            .I(\COUNTER.counterZ0Z_3 ));
    LocalMux I__3656 (
            .O(N__17506),
            .I(\COUNTER.counterZ0Z_3 ));
    InMux I__3655 (
            .O(N__17501),
            .I(N__17497));
    InMux I__3654 (
            .O(N__17500),
            .I(N__17494));
    LocalMux I__3653 (
            .O(N__17497),
            .I(\ALL_SYS_PWRGD.countZ0Z_7 ));
    LocalMux I__3652 (
            .O(N__17494),
            .I(\ALL_SYS_PWRGD.countZ0Z_7 ));
    InMux I__3651 (
            .O(N__17489),
            .I(N__17485));
    InMux I__3650 (
            .O(N__17488),
            .I(N__17482));
    LocalMux I__3649 (
            .O(N__17485),
            .I(\ALL_SYS_PWRGD.countZ0Z_8 ));
    LocalMux I__3648 (
            .O(N__17482),
            .I(\ALL_SYS_PWRGD.countZ0Z_8 ));
    CascadeMux I__3647 (
            .O(N__17477),
            .I(N__17473));
    InMux I__3646 (
            .O(N__17476),
            .I(N__17470));
    InMux I__3645 (
            .O(N__17473),
            .I(N__17467));
    LocalMux I__3644 (
            .O(N__17470),
            .I(\ALL_SYS_PWRGD.countZ0Z_6 ));
    LocalMux I__3643 (
            .O(N__17467),
            .I(\ALL_SYS_PWRGD.countZ0Z_6 ));
    InMux I__3642 (
            .O(N__17462),
            .I(N__17458));
    InMux I__3641 (
            .O(N__17461),
            .I(N__17455));
    LocalMux I__3640 (
            .O(N__17458),
            .I(\ALL_SYS_PWRGD.countZ0Z_4 ));
    LocalMux I__3639 (
            .O(N__17455),
            .I(\ALL_SYS_PWRGD.countZ0Z_4 ));
    InMux I__3638 (
            .O(N__17450),
            .I(N__17446));
    InMux I__3637 (
            .O(N__17449),
            .I(N__17443));
    LocalMux I__3636 (
            .O(N__17446),
            .I(\ALL_SYS_PWRGD.countZ0Z_14 ));
    LocalMux I__3635 (
            .O(N__17443),
            .I(\ALL_SYS_PWRGD.countZ0Z_14 ));
    InMux I__3634 (
            .O(N__17438),
            .I(N__17434));
    InMux I__3633 (
            .O(N__17437),
            .I(N__17431));
    LocalMux I__3632 (
            .O(N__17434),
            .I(\ALL_SYS_PWRGD.countZ0Z_15 ));
    LocalMux I__3631 (
            .O(N__17431),
            .I(\ALL_SYS_PWRGD.countZ0Z_15 ));
    CascadeMux I__3630 (
            .O(N__17426),
            .I(N__17422));
    InMux I__3629 (
            .O(N__17425),
            .I(N__17419));
    InMux I__3628 (
            .O(N__17422),
            .I(N__17416));
    LocalMux I__3627 (
            .O(N__17419),
            .I(\ALL_SYS_PWRGD.countZ0Z_13 ));
    LocalMux I__3626 (
            .O(N__17416),
            .I(\ALL_SYS_PWRGD.countZ0Z_13 ));
    InMux I__3625 (
            .O(N__17411),
            .I(N__17407));
    InMux I__3624 (
            .O(N__17410),
            .I(N__17404));
    LocalMux I__3623 (
            .O(N__17407),
            .I(\ALL_SYS_PWRGD.countZ0Z_12 ));
    LocalMux I__3622 (
            .O(N__17404),
            .I(\ALL_SYS_PWRGD.countZ0Z_12 ));
    InMux I__3621 (
            .O(N__17399),
            .I(N__17396));
    LocalMux I__3620 (
            .O(N__17396),
            .I(\ALL_SYS_PWRGD.un4_count_10 ));
    CascadeMux I__3619 (
            .O(N__17393),
            .I(\ALL_SYS_PWRGD.un4_count_11_cascade_ ));
    InMux I__3618 (
            .O(N__17390),
            .I(N__17387));
    LocalMux I__3617 (
            .O(N__17387),
            .I(\ALL_SYS_PWRGD.un4_count_8 ));
    InMux I__3616 (
            .O(N__17384),
            .I(N__17380));
    InMux I__3615 (
            .O(N__17383),
            .I(N__17377));
    LocalMux I__3614 (
            .O(N__17380),
            .I(\ALL_SYS_PWRGD.countZ0Z_1 ));
    LocalMux I__3613 (
            .O(N__17377),
            .I(\ALL_SYS_PWRGD.countZ0Z_1 ));
    InMux I__3612 (
            .O(N__17372),
            .I(N__17368));
    InMux I__3611 (
            .O(N__17371),
            .I(N__17365));
    LocalMux I__3610 (
            .O(N__17368),
            .I(\ALL_SYS_PWRGD.countZ0Z_9 ));
    LocalMux I__3609 (
            .O(N__17365),
            .I(\ALL_SYS_PWRGD.countZ0Z_9 ));
    CascadeMux I__3608 (
            .O(N__17360),
            .I(N__17356));
    InMux I__3607 (
            .O(N__17359),
            .I(N__17353));
    InMux I__3606 (
            .O(N__17356),
            .I(N__17350));
    LocalMux I__3605 (
            .O(N__17353),
            .I(\ALL_SYS_PWRGD.countZ0Z_10 ));
    LocalMux I__3604 (
            .O(N__17350),
            .I(\ALL_SYS_PWRGD.countZ0Z_10 ));
    InMux I__3603 (
            .O(N__17345),
            .I(N__17341));
    InMux I__3602 (
            .O(N__17344),
            .I(N__17338));
    LocalMux I__3601 (
            .O(N__17341),
            .I(\ALL_SYS_PWRGD.countZ0Z_0 ));
    LocalMux I__3600 (
            .O(N__17338),
            .I(\ALL_SYS_PWRGD.countZ0Z_0 ));
    InMux I__3599 (
            .O(N__17333),
            .I(\COUNTER.counter_1_cry_27 ));
    InMux I__3598 (
            .O(N__17330),
            .I(\COUNTER.counter_1_cry_28 ));
    InMux I__3597 (
            .O(N__17327),
            .I(\COUNTER.counter_1_cry_29 ));
    InMux I__3596 (
            .O(N__17324),
            .I(\COUNTER.counter_1_cry_30 ));
    InMux I__3595 (
            .O(N__17321),
            .I(N__17317));
    InMux I__3594 (
            .O(N__17320),
            .I(N__17314));
    LocalMux I__3593 (
            .O(N__17317),
            .I(\COUNTER.counterZ0Z_22 ));
    LocalMux I__3592 (
            .O(N__17314),
            .I(\COUNTER.counterZ0Z_22 ));
    InMux I__3591 (
            .O(N__17309),
            .I(N__17305));
    InMux I__3590 (
            .O(N__17308),
            .I(N__17302));
    LocalMux I__3589 (
            .O(N__17305),
            .I(\COUNTER.counterZ0Z_21 ));
    LocalMux I__3588 (
            .O(N__17302),
            .I(\COUNTER.counterZ0Z_21 ));
    CascadeMux I__3587 (
            .O(N__17297),
            .I(N__17293));
    InMux I__3586 (
            .O(N__17296),
            .I(N__17290));
    InMux I__3585 (
            .O(N__17293),
            .I(N__17287));
    LocalMux I__3584 (
            .O(N__17290),
            .I(\COUNTER.counterZ0Z_23 ));
    LocalMux I__3583 (
            .O(N__17287),
            .I(\COUNTER.counterZ0Z_23 ));
    InMux I__3582 (
            .O(N__17282),
            .I(N__17278));
    InMux I__3581 (
            .O(N__17281),
            .I(N__17275));
    LocalMux I__3580 (
            .O(N__17278),
            .I(\COUNTER.counterZ0Z_20 ));
    LocalMux I__3579 (
            .O(N__17275),
            .I(\COUNTER.counterZ0Z_20 ));
    InMux I__3578 (
            .O(N__17270),
            .I(N__17266));
    InMux I__3577 (
            .O(N__17269),
            .I(N__17263));
    LocalMux I__3576 (
            .O(N__17266),
            .I(\ALL_SYS_PWRGD.countZ0Z_5 ));
    LocalMux I__3575 (
            .O(N__17263),
            .I(\ALL_SYS_PWRGD.countZ0Z_5 ));
    InMux I__3574 (
            .O(N__17258),
            .I(N__17254));
    InMux I__3573 (
            .O(N__17257),
            .I(N__17251));
    LocalMux I__3572 (
            .O(N__17254),
            .I(\ALL_SYS_PWRGD.countZ0Z_3 ));
    LocalMux I__3571 (
            .O(N__17251),
            .I(\ALL_SYS_PWRGD.countZ0Z_3 ));
    CascadeMux I__3570 (
            .O(N__17246),
            .I(N__17242));
    InMux I__3569 (
            .O(N__17245),
            .I(N__17239));
    InMux I__3568 (
            .O(N__17242),
            .I(N__17236));
    LocalMux I__3567 (
            .O(N__17239),
            .I(\ALL_SYS_PWRGD.countZ0Z_11 ));
    LocalMux I__3566 (
            .O(N__17236),
            .I(\ALL_SYS_PWRGD.countZ0Z_11 ));
    InMux I__3565 (
            .O(N__17231),
            .I(N__17227));
    InMux I__3564 (
            .O(N__17230),
            .I(N__17224));
    LocalMux I__3563 (
            .O(N__17227),
            .I(\ALL_SYS_PWRGD.countZ0Z_2 ));
    LocalMux I__3562 (
            .O(N__17224),
            .I(\ALL_SYS_PWRGD.countZ0Z_2 ));
    InMux I__3561 (
            .O(N__17219),
            .I(N__17215));
    InMux I__3560 (
            .O(N__17218),
            .I(N__17212));
    LocalMux I__3559 (
            .O(N__17215),
            .I(\COUNTER.counterZ0Z_26 ));
    LocalMux I__3558 (
            .O(N__17212),
            .I(\COUNTER.counterZ0Z_26 ));
    InMux I__3557 (
            .O(N__17207),
            .I(N__17203));
    InMux I__3556 (
            .O(N__17206),
            .I(N__17200));
    LocalMux I__3555 (
            .O(N__17203),
            .I(\COUNTER.counterZ0Z_25 ));
    LocalMux I__3554 (
            .O(N__17200),
            .I(\COUNTER.counterZ0Z_25 ));
    CascadeMux I__3553 (
            .O(N__17195),
            .I(N__17191));
    InMux I__3552 (
            .O(N__17194),
            .I(N__17188));
    InMux I__3551 (
            .O(N__17191),
            .I(N__17185));
    LocalMux I__3550 (
            .O(N__17188),
            .I(\COUNTER.counterZ0Z_27 ));
    LocalMux I__3549 (
            .O(N__17185),
            .I(\COUNTER.counterZ0Z_27 ));
    InMux I__3548 (
            .O(N__17180),
            .I(N__17176));
    InMux I__3547 (
            .O(N__17179),
            .I(N__17173));
    LocalMux I__3546 (
            .O(N__17176),
            .I(N__17170));
    LocalMux I__3545 (
            .O(N__17173),
            .I(\COUNTER.counterZ0Z_24 ));
    Odrv4 I__3544 (
            .O(N__17170),
            .I(\COUNTER.counterZ0Z_24 ));
    InMux I__3543 (
            .O(N__17165),
            .I(N__17161));
    InMux I__3542 (
            .O(N__17164),
            .I(N__17158));
    LocalMux I__3541 (
            .O(N__17161),
            .I(\COUNTER.counterZ0Z_30 ));
    LocalMux I__3540 (
            .O(N__17158),
            .I(\COUNTER.counterZ0Z_30 ));
    InMux I__3539 (
            .O(N__17153),
            .I(N__17149));
    InMux I__3538 (
            .O(N__17152),
            .I(N__17146));
    LocalMux I__3537 (
            .O(N__17149),
            .I(\COUNTER.counterZ0Z_28 ));
    LocalMux I__3536 (
            .O(N__17146),
            .I(\COUNTER.counterZ0Z_28 ));
    CascadeMux I__3535 (
            .O(N__17141),
            .I(N__17137));
    InMux I__3534 (
            .O(N__17140),
            .I(N__17134));
    InMux I__3533 (
            .O(N__17137),
            .I(N__17131));
    LocalMux I__3532 (
            .O(N__17134),
            .I(\COUNTER.counterZ0Z_29 ));
    LocalMux I__3531 (
            .O(N__17131),
            .I(\COUNTER.counterZ0Z_29 ));
    InMux I__3530 (
            .O(N__17126),
            .I(N__17122));
    InMux I__3529 (
            .O(N__17125),
            .I(N__17119));
    LocalMux I__3528 (
            .O(N__17122),
            .I(\COUNTER.counterZ0Z_31 ));
    LocalMux I__3527 (
            .O(N__17119),
            .I(\COUNTER.counterZ0Z_31 ));
    InMux I__3526 (
            .O(N__17114),
            .I(\COUNTER.counter_1_cry_18 ));
    InMux I__3525 (
            .O(N__17111),
            .I(\COUNTER.counter_1_cry_19 ));
    InMux I__3524 (
            .O(N__17108),
            .I(\COUNTER.counter_1_cry_20 ));
    InMux I__3523 (
            .O(N__17105),
            .I(\COUNTER.counter_1_cry_21 ));
    InMux I__3522 (
            .O(N__17102),
            .I(\COUNTER.counter_1_cry_22 ));
    InMux I__3521 (
            .O(N__17099),
            .I(\COUNTER.counter_1_cry_23 ));
    InMux I__3520 (
            .O(N__17096),
            .I(bfn_9_4_0_));
    InMux I__3519 (
            .O(N__17093),
            .I(\COUNTER.counter_1_cry_25 ));
    InMux I__3518 (
            .O(N__17090),
            .I(\COUNTER.counter_1_cry_26 ));
    InMux I__3517 (
            .O(N__17087),
            .I(\COUNTER.counter_1_cry_9 ));
    InMux I__3516 (
            .O(N__17084),
            .I(\COUNTER.counter_1_cry_10 ));
    InMux I__3515 (
            .O(N__17081),
            .I(\COUNTER.counter_1_cry_11 ));
    InMux I__3514 (
            .O(N__17078),
            .I(\COUNTER.counter_1_cry_12 ));
    InMux I__3513 (
            .O(N__17075),
            .I(\COUNTER.counter_1_cry_13 ));
    InMux I__3512 (
            .O(N__17072),
            .I(\COUNTER.counter_1_cry_14 ));
    InMux I__3511 (
            .O(N__17069),
            .I(\COUNTER.counter_1_cry_15 ));
    InMux I__3510 (
            .O(N__17066),
            .I(bfn_9_3_0_));
    InMux I__3509 (
            .O(N__17063),
            .I(\COUNTER.counter_1_cry_17 ));
    InMux I__3508 (
            .O(N__17060),
            .I(\COUNTER.counter_1_cry_1 ));
    InMux I__3507 (
            .O(N__17057),
            .I(\COUNTER.counter_1_cry_2 ));
    InMux I__3506 (
            .O(N__17054),
            .I(\COUNTER.counter_1_cry_3 ));
    InMux I__3505 (
            .O(N__17051),
            .I(N__17046));
    InMux I__3504 (
            .O(N__17050),
            .I(N__17041));
    InMux I__3503 (
            .O(N__17049),
            .I(N__17041));
    LocalMux I__3502 (
            .O(N__17046),
            .I(\COUNTER.counterZ0Z_5 ));
    LocalMux I__3501 (
            .O(N__17041),
            .I(\COUNTER.counterZ0Z_5 ));
    InMux I__3500 (
            .O(N__17036),
            .I(N__17033));
    LocalMux I__3499 (
            .O(N__17033),
            .I(\COUNTER.counter_1_cry_4_THRU_CO ));
    InMux I__3498 (
            .O(N__17030),
            .I(\COUNTER.counter_1_cry_4 ));
    CascadeMux I__3497 (
            .O(N__17027),
            .I(N__17023));
    InMux I__3496 (
            .O(N__17026),
            .I(N__17019));
    InMux I__3495 (
            .O(N__17023),
            .I(N__17014));
    InMux I__3494 (
            .O(N__17022),
            .I(N__17014));
    LocalMux I__3493 (
            .O(N__17019),
            .I(\COUNTER.counterZ0Z_6 ));
    LocalMux I__3492 (
            .O(N__17014),
            .I(\COUNTER.counterZ0Z_6 ));
    InMux I__3491 (
            .O(N__17009),
            .I(N__17006));
    LocalMux I__3490 (
            .O(N__17006),
            .I(\COUNTER.counter_1_cry_5_THRU_CO ));
    InMux I__3489 (
            .O(N__17003),
            .I(\COUNTER.counter_1_cry_5 ));
    CascadeMux I__3488 (
            .O(N__17000),
            .I(N__16996));
    InMux I__3487 (
            .O(N__16999),
            .I(N__16993));
    InMux I__3486 (
            .O(N__16996),
            .I(N__16990));
    LocalMux I__3485 (
            .O(N__16993),
            .I(\COUNTER.counterZ0Z_7 ));
    LocalMux I__3484 (
            .O(N__16990),
            .I(\COUNTER.counterZ0Z_7 ));
    InMux I__3483 (
            .O(N__16985),
            .I(\COUNTER.counter_1_cry_6 ));
    InMux I__3482 (
            .O(N__16982),
            .I(\COUNTER.counter_1_cry_7 ));
    InMux I__3481 (
            .O(N__16979),
            .I(bfn_9_2_0_));
    InMux I__3480 (
            .O(N__16976),
            .I(\VPP_VDDQ.un1_count_1_cry_8 ));
    InMux I__3479 (
            .O(N__16973),
            .I(\VPP_VDDQ.un1_count_1_cry_9 ));
    InMux I__3478 (
            .O(N__16970),
            .I(\VPP_VDDQ.un1_count_1_cry_10 ));
    InMux I__3477 (
            .O(N__16967),
            .I(\VPP_VDDQ.un1_count_1_cry_11 ));
    InMux I__3476 (
            .O(N__16964),
            .I(\VPP_VDDQ.un1_count_1_cry_12 ));
    InMux I__3475 (
            .O(N__16961),
            .I(\VPP_VDDQ.un1_count_1_cry_13 ));
    InMux I__3474 (
            .O(N__16958),
            .I(bfn_8_16_0_));
    CEMux I__3473 (
            .O(N__16955),
            .I(N__16952));
    LocalMux I__3472 (
            .O(N__16952),
            .I(N__16949));
    Odrv4 I__3471 (
            .O(N__16949),
            .I(\VPP_VDDQ.N_65_1 ));
    SRMux I__3470 (
            .O(N__16946),
            .I(N__16943));
    LocalMux I__3469 (
            .O(N__16943),
            .I(N__16939));
    SRMux I__3468 (
            .O(N__16942),
            .I(N__16936));
    Span4Mux_s1_v I__3467 (
            .O(N__16939),
            .I(N__16931));
    LocalMux I__3466 (
            .O(N__16936),
            .I(N__16931));
    Span4Mux_v I__3465 (
            .O(N__16931),
            .I(N__16927));
    SRMux I__3464 (
            .O(N__16930),
            .I(N__16924));
    Sp12to4 I__3463 (
            .O(N__16927),
            .I(N__16918));
    LocalMux I__3462 (
            .O(N__16924),
            .I(N__16918));
    InMux I__3461 (
            .O(N__16923),
            .I(N__16915));
    Odrv12 I__3460 (
            .O(N__16918),
            .I(\VPP_VDDQ.curr_state_RNIGR9S7Z0Z_0 ));
    LocalMux I__3459 (
            .O(N__16915),
            .I(\VPP_VDDQ.curr_state_RNIGR9S7Z0Z_0 ));
    InMux I__3458 (
            .O(N__16910),
            .I(N__16905));
    InMux I__3457 (
            .O(N__16909),
            .I(N__16900));
    InMux I__3456 (
            .O(N__16908),
            .I(N__16900));
    LocalMux I__3455 (
            .O(N__16905),
            .I(\COUNTER.counterZ0Z_1 ));
    LocalMux I__3454 (
            .O(N__16900),
            .I(\COUNTER.counterZ0Z_1 ));
    InMux I__3453 (
            .O(N__16895),
            .I(N__16891));
    CascadeMux I__3452 (
            .O(N__16894),
            .I(N__16888));
    LocalMux I__3451 (
            .O(N__16891),
            .I(N__16885));
    InMux I__3450 (
            .O(N__16888),
            .I(N__16882));
    Odrv4 I__3449 (
            .O(N__16885),
            .I(\VPP_VDDQ.N_108_i ));
    LocalMux I__3448 (
            .O(N__16882),
            .I(\VPP_VDDQ.N_108_i ));
    InMux I__3447 (
            .O(N__16877),
            .I(\VPP_VDDQ.un1_count_1_cry_0 ));
    InMux I__3446 (
            .O(N__16874),
            .I(\VPP_VDDQ.un1_count_1_cry_1 ));
    InMux I__3445 (
            .O(N__16871),
            .I(\VPP_VDDQ.un1_count_1_cry_2 ));
    InMux I__3444 (
            .O(N__16868),
            .I(\VPP_VDDQ.un1_count_1_cry_3 ));
    InMux I__3443 (
            .O(N__16865),
            .I(\VPP_VDDQ.un1_count_1_cry_4 ));
    InMux I__3442 (
            .O(N__16862),
            .I(\VPP_VDDQ.un1_count_1_cry_5 ));
    InMux I__3441 (
            .O(N__16859),
            .I(\VPP_VDDQ.un1_count_1_cry_6 ));
    InMux I__3440 (
            .O(N__16856),
            .I(bfn_8_15_0_));
    InMux I__3439 (
            .O(N__16853),
            .I(bfn_8_12_0_));
    InMux I__3438 (
            .O(N__16850),
            .I(\RSMRST_PWRGD.un1_count_1_cry_8 ));
    InMux I__3437 (
            .O(N__16847),
            .I(\RSMRST_PWRGD.un1_count_1_cry_9 ));
    InMux I__3436 (
            .O(N__16844),
            .I(\RSMRST_PWRGD.un1_count_1_cry_10 ));
    InMux I__3435 (
            .O(N__16841),
            .I(\RSMRST_PWRGD.un1_count_1_cry_11 ));
    InMux I__3434 (
            .O(N__16838),
            .I(\RSMRST_PWRGD.un1_count_1_cry_12 ));
    InMux I__3433 (
            .O(N__16835),
            .I(\RSMRST_PWRGD.un1_count_1_cry_13 ));
    InMux I__3432 (
            .O(N__16832),
            .I(bfn_8_13_0_));
    CascadeMux I__3431 (
            .O(N__16829),
            .I(\POWERLED.count_off_1_sqmuxa_i_a6_0_1_cascade_ ));
    InMux I__3430 (
            .O(N__16826),
            .I(N__16822));
    InMux I__3429 (
            .O(N__16825),
            .I(N__16819));
    LocalMux I__3428 (
            .O(N__16822),
            .I(\POWERLED.N_136 ));
    LocalMux I__3427 (
            .O(N__16819),
            .I(\POWERLED.N_136 ));
    InMux I__3426 (
            .O(N__16814),
            .I(N__16811));
    LocalMux I__3425 (
            .O(N__16811),
            .I(N__16808));
    Odrv4 I__3424 (
            .O(N__16808),
            .I(\POWERLED.count_off_1_sqmuxa_i_a6_0_3 ));
    InMux I__3423 (
            .O(N__16805),
            .I(\RSMRST_PWRGD.un1_count_1_cry_0 ));
    InMux I__3422 (
            .O(N__16802),
            .I(\RSMRST_PWRGD.un1_count_1_cry_1 ));
    InMux I__3421 (
            .O(N__16799),
            .I(\RSMRST_PWRGD.un1_count_1_cry_2 ));
    InMux I__3420 (
            .O(N__16796),
            .I(\RSMRST_PWRGD.un1_count_1_cry_3 ));
    InMux I__3419 (
            .O(N__16793),
            .I(\RSMRST_PWRGD.un1_count_1_cry_4 ));
    InMux I__3418 (
            .O(N__16790),
            .I(\RSMRST_PWRGD.un1_count_1_cry_5 ));
    InMux I__3417 (
            .O(N__16787),
            .I(\RSMRST_PWRGD.un1_count_1_cry_6 ));
    InMux I__3416 (
            .O(N__16784),
            .I(N__16781));
    LocalMux I__3415 (
            .O(N__16781),
            .I(N__16778));
    Odrv4 I__3414 (
            .O(N__16778),
            .I(\POWERLED.N_366_1 ));
    InMux I__3413 (
            .O(N__16775),
            .I(N__16762));
    InMux I__3412 (
            .O(N__16774),
            .I(N__16762));
    InMux I__3411 (
            .O(N__16773),
            .I(N__16762));
    InMux I__3410 (
            .O(N__16772),
            .I(N__16753));
    InMux I__3409 (
            .O(N__16771),
            .I(N__16746));
    InMux I__3408 (
            .O(N__16770),
            .I(N__16746));
    InMux I__3407 (
            .O(N__16769),
            .I(N__16746));
    LocalMux I__3406 (
            .O(N__16762),
            .I(N__16743));
    InMux I__3405 (
            .O(N__16761),
            .I(N__16740));
    InMux I__3404 (
            .O(N__16760),
            .I(N__16732));
    InMux I__3403 (
            .O(N__16759),
            .I(N__16723));
    InMux I__3402 (
            .O(N__16758),
            .I(N__16723));
    InMux I__3401 (
            .O(N__16757),
            .I(N__16723));
    InMux I__3400 (
            .O(N__16756),
            .I(N__16723));
    LocalMux I__3399 (
            .O(N__16753),
            .I(N__16720));
    LocalMux I__3398 (
            .O(N__16746),
            .I(N__16717));
    Span4Mux_v I__3397 (
            .O(N__16743),
            .I(N__16712));
    LocalMux I__3396 (
            .O(N__16740),
            .I(N__16712));
    InMux I__3395 (
            .O(N__16739),
            .I(N__16709));
    InMux I__3394 (
            .O(N__16738),
            .I(N__16700));
    InMux I__3393 (
            .O(N__16737),
            .I(N__16700));
    InMux I__3392 (
            .O(N__16736),
            .I(N__16700));
    InMux I__3391 (
            .O(N__16735),
            .I(N__16700));
    LocalMux I__3390 (
            .O(N__16732),
            .I(N__16697));
    LocalMux I__3389 (
            .O(N__16723),
            .I(N__16692));
    Span4Mux_h I__3388 (
            .O(N__16720),
            .I(N__16692));
    Span4Mux_h I__3387 (
            .O(N__16717),
            .I(N__16687));
    Span4Mux_h I__3386 (
            .O(N__16712),
            .I(N__16687));
    LocalMux I__3385 (
            .O(N__16709),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    LocalMux I__3384 (
            .O(N__16700),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    Odrv4 I__3383 (
            .O(N__16697),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    Odrv4 I__3382 (
            .O(N__16692),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    Odrv4 I__3381 (
            .O(N__16687),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    InMux I__3380 (
            .O(N__16676),
            .I(N__16673));
    LocalMux I__3379 (
            .O(N__16673),
            .I(N__16669));
    CascadeMux I__3378 (
            .O(N__16672),
            .I(N__16666));
    Span4Mux_h I__3377 (
            .O(N__16669),
            .I(N__16663));
    InMux I__3376 (
            .O(N__16666),
            .I(N__16660));
    Odrv4 I__3375 (
            .O(N__16663),
            .I(\POWERLED.N_177_5 ));
    LocalMux I__3374 (
            .O(N__16660),
            .I(\POWERLED.N_177_5 ));
    CascadeMux I__3373 (
            .O(N__16655),
            .I(\POWERLED.count_clk_0_sqmuxa_5_0_o2_0_0_cascade_ ));
    InMux I__3372 (
            .O(N__16652),
            .I(N__16649));
    LocalMux I__3371 (
            .O(N__16649),
            .I(N__16646));
    Span4Mux_v I__3370 (
            .O(N__16646),
            .I(N__16642));
    InMux I__3369 (
            .O(N__16645),
            .I(N__16639));
    Odrv4 I__3368 (
            .O(N__16642),
            .I(\POWERLED.N_141 ));
    LocalMux I__3367 (
            .O(N__16639),
            .I(\POWERLED.N_141 ));
    CascadeMux I__3366 (
            .O(N__16634),
            .I(\POWERLED.N_136_cascade_ ));
    InMux I__3365 (
            .O(N__16631),
            .I(N__16624));
    InMux I__3364 (
            .O(N__16630),
            .I(N__16624));
    InMux I__3363 (
            .O(N__16629),
            .I(N__16620));
    LocalMux I__3362 (
            .O(N__16624),
            .I(N__16617));
    InMux I__3361 (
            .O(N__16623),
            .I(N__16614));
    LocalMux I__3360 (
            .O(N__16620),
            .I(\POWERLED.N_146 ));
    Odrv4 I__3359 (
            .O(N__16617),
            .I(\POWERLED.N_146 ));
    LocalMux I__3358 (
            .O(N__16614),
            .I(\POWERLED.N_146 ));
    InMux I__3357 (
            .O(N__16607),
            .I(N__16604));
    LocalMux I__3356 (
            .O(N__16604),
            .I(N__16601));
    Odrv4 I__3355 (
            .O(N__16601),
            .I(\POWERLED.count_clk_0_sqmuxa_5_0_a6_1 ));
    InMux I__3354 (
            .O(N__16598),
            .I(N__16595));
    LocalMux I__3353 (
            .O(N__16595),
            .I(\POWERLED.count_clk_0_sqmuxa_5_0_o2_4 ));
    IoInMux I__3352 (
            .O(N__16592),
            .I(N__16587));
    CascadeMux I__3351 (
            .O(N__16591),
            .I(N__16584));
    CascadeMux I__3350 (
            .O(N__16590),
            .I(N__16578));
    LocalMux I__3349 (
            .O(N__16587),
            .I(N__16574));
    InMux I__3348 (
            .O(N__16584),
            .I(N__16567));
    InMux I__3347 (
            .O(N__16583),
            .I(N__16567));
    InMux I__3346 (
            .O(N__16582),
            .I(N__16567));
    InMux I__3345 (
            .O(N__16581),
            .I(N__16564));
    InMux I__3344 (
            .O(N__16578),
            .I(N__16561));
    CascadeMux I__3343 (
            .O(N__16577),
            .I(N__16558));
    IoSpan4Mux I__3342 (
            .O(N__16574),
            .I(N__16553));
    LocalMux I__3341 (
            .O(N__16567),
            .I(N__16546));
    LocalMux I__3340 (
            .O(N__16564),
            .I(N__16546));
    LocalMux I__3339 (
            .O(N__16561),
            .I(N__16546));
    InMux I__3338 (
            .O(N__16558),
            .I(N__16543));
    InMux I__3337 (
            .O(N__16557),
            .I(N__16538));
    InMux I__3336 (
            .O(N__16556),
            .I(N__16538));
    Span4Mux_s2_h I__3335 (
            .O(N__16553),
            .I(N__16534));
    Span4Mux_v I__3334 (
            .O(N__16546),
            .I(N__16531));
    LocalMux I__3333 (
            .O(N__16543),
            .I(N__16528));
    LocalMux I__3332 (
            .O(N__16538),
            .I(N__16525));
    InMux I__3331 (
            .O(N__16537),
            .I(N__16522));
    Span4Mux_h I__3330 (
            .O(N__16534),
            .I(N__16517));
    Span4Mux_v I__3329 (
            .O(N__16531),
            .I(N__16517));
    Sp12to4 I__3328 (
            .O(N__16528),
            .I(N__16510));
    Sp12to4 I__3327 (
            .O(N__16525),
            .I(N__16510));
    LocalMux I__3326 (
            .O(N__16522),
            .I(N__16510));
    Sp12to4 I__3325 (
            .O(N__16517),
            .I(N__16505));
    Span12Mux_v I__3324 (
            .O(N__16510),
            .I(N__16505));
    Odrv12 I__3323 (
            .O(N__16505),
            .I(gpio_fpga_soc_4));
    InMux I__3322 (
            .O(N__16502),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_12 ));
    InMux I__3321 (
            .O(N__16499),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_13 ));
    InMux I__3320 (
            .O(N__16496),
            .I(bfn_8_7_0_));
    CascadeMux I__3319 (
            .O(N__16493),
            .I(N__16490));
    InMux I__3318 (
            .O(N__16490),
            .I(N__16486));
    InMux I__3317 (
            .O(N__16489),
            .I(N__16483));
    LocalMux I__3316 (
            .O(N__16486),
            .I(N__16480));
    LocalMux I__3315 (
            .O(N__16483),
            .I(N__16477));
    Span4Mux_h I__3314 (
            .O(N__16480),
            .I(N__16474));
    Odrv4 I__3313 (
            .O(N__16477),
            .I(\POWERLED.dutycycle_RNIO18NZ0Z_9 ));
    Odrv4 I__3312 (
            .O(N__16474),
            .I(\POWERLED.dutycycle_RNIO18NZ0Z_9 ));
    CascadeMux I__3311 (
            .O(N__16469),
            .I(N__16462));
    InMux I__3310 (
            .O(N__16468),
            .I(N__16453));
    InMux I__3309 (
            .O(N__16467),
            .I(N__16453));
    CascadeMux I__3308 (
            .O(N__16466),
            .I(N__16449));
    InMux I__3307 (
            .O(N__16465),
            .I(N__16445));
    InMux I__3306 (
            .O(N__16462),
            .I(N__16442));
    InMux I__3305 (
            .O(N__16461),
            .I(N__16439));
    InMux I__3304 (
            .O(N__16460),
            .I(N__16434));
    InMux I__3303 (
            .O(N__16459),
            .I(N__16434));
    InMux I__3302 (
            .O(N__16458),
            .I(N__16431));
    LocalMux I__3301 (
            .O(N__16453),
            .I(N__16428));
    InMux I__3300 (
            .O(N__16452),
            .I(N__16425));
    InMux I__3299 (
            .O(N__16449),
            .I(N__16420));
    InMux I__3298 (
            .O(N__16448),
            .I(N__16420));
    LocalMux I__3297 (
            .O(N__16445),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__3296 (
            .O(N__16442),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__3295 (
            .O(N__16439),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__3294 (
            .O(N__16434),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__3293 (
            .O(N__16431),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    Odrv12 I__3292 (
            .O(N__16428),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__3291 (
            .O(N__16425),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__3290 (
            .O(N__16420),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    CascadeMux I__3289 (
            .O(N__16403),
            .I(N__16399));
    CascadeMux I__3288 (
            .O(N__16402),
            .I(N__16390));
    InMux I__3287 (
            .O(N__16399),
            .I(N__16381));
    InMux I__3286 (
            .O(N__16398),
            .I(N__16381));
    InMux I__3285 (
            .O(N__16397),
            .I(N__16381));
    InMux I__3284 (
            .O(N__16396),
            .I(N__16378));
    InMux I__3283 (
            .O(N__16395),
            .I(N__16375));
    InMux I__3282 (
            .O(N__16394),
            .I(N__16372));
    InMux I__3281 (
            .O(N__16393),
            .I(N__16367));
    InMux I__3280 (
            .O(N__16390),
            .I(N__16367));
    InMux I__3279 (
            .O(N__16389),
            .I(N__16362));
    InMux I__3278 (
            .O(N__16388),
            .I(N__16362));
    LocalMux I__3277 (
            .O(N__16381),
            .I(N__16359));
    LocalMux I__3276 (
            .O(N__16378),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__3275 (
            .O(N__16375),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__3274 (
            .O(N__16372),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__3273 (
            .O(N__16367),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__3272 (
            .O(N__16362),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    Odrv4 I__3271 (
            .O(N__16359),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    CascadeMux I__3270 (
            .O(N__16346),
            .I(N__16340));
    CascadeMux I__3269 (
            .O(N__16345),
            .I(N__16336));
    CascadeMux I__3268 (
            .O(N__16344),
            .I(N__16331));
    InMux I__3267 (
            .O(N__16343),
            .I(N__16326));
    InMux I__3266 (
            .O(N__16340),
            .I(N__16323));
    InMux I__3265 (
            .O(N__16339),
            .I(N__16318));
    InMux I__3264 (
            .O(N__16336),
            .I(N__16318));
    InMux I__3263 (
            .O(N__16335),
            .I(N__16315));
    InMux I__3262 (
            .O(N__16334),
            .I(N__16312));
    InMux I__3261 (
            .O(N__16331),
            .I(N__16305));
    InMux I__3260 (
            .O(N__16330),
            .I(N__16305));
    InMux I__3259 (
            .O(N__16329),
            .I(N__16305));
    LocalMux I__3258 (
            .O(N__16326),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__3257 (
            .O(N__16323),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__3256 (
            .O(N__16318),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__3255 (
            .O(N__16315),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__3254 (
            .O(N__16312),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__3253 (
            .O(N__16305),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    CascadeMux I__3252 (
            .O(N__16292),
            .I(N__16289));
    InMux I__3251 (
            .O(N__16289),
            .I(N__16276));
    InMux I__3250 (
            .O(N__16288),
            .I(N__16276));
    InMux I__3249 (
            .O(N__16287),
            .I(N__16273));
    InMux I__3248 (
            .O(N__16286),
            .I(N__16268));
    InMux I__3247 (
            .O(N__16285),
            .I(N__16268));
    InMux I__3246 (
            .O(N__16284),
            .I(N__16265));
    InMux I__3245 (
            .O(N__16283),
            .I(N__16258));
    InMux I__3244 (
            .O(N__16282),
            .I(N__16258));
    InMux I__3243 (
            .O(N__16281),
            .I(N__16258));
    LocalMux I__3242 (
            .O(N__16276),
            .I(N__16255));
    LocalMux I__3241 (
            .O(N__16273),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__3240 (
            .O(N__16268),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__3239 (
            .O(N__16265),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__3238 (
            .O(N__16258),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv4 I__3237 (
            .O(N__16255),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    CascadeMux I__3236 (
            .O(N__16244),
            .I(N__16239));
    InMux I__3235 (
            .O(N__16243),
            .I(N__16232));
    InMux I__3234 (
            .O(N__16242),
            .I(N__16228));
    InMux I__3233 (
            .O(N__16239),
            .I(N__16225));
    InMux I__3232 (
            .O(N__16238),
            .I(N__16222));
    InMux I__3231 (
            .O(N__16237),
            .I(N__16219));
    InMux I__3230 (
            .O(N__16236),
            .I(N__16216));
    InMux I__3229 (
            .O(N__16235),
            .I(N__16213));
    LocalMux I__3228 (
            .O(N__16232),
            .I(N__16210));
    InMux I__3227 (
            .O(N__16231),
            .I(N__16207));
    LocalMux I__3226 (
            .O(N__16228),
            .I(N__16204));
    LocalMux I__3225 (
            .O(N__16225),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__3224 (
            .O(N__16222),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__3223 (
            .O(N__16219),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__3222 (
            .O(N__16216),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__3221 (
            .O(N__16213),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__3220 (
            .O(N__16210),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__3219 (
            .O(N__16207),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__3218 (
            .O(N__16204),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    CascadeMux I__3217 (
            .O(N__16187),
            .I(N__16181));
    InMux I__3216 (
            .O(N__16186),
            .I(N__16177));
    InMux I__3215 (
            .O(N__16185),
            .I(N__16174));
    CascadeMux I__3214 (
            .O(N__16184),
            .I(N__16169));
    InMux I__3213 (
            .O(N__16181),
            .I(N__16164));
    InMux I__3212 (
            .O(N__16180),
            .I(N__16161));
    LocalMux I__3211 (
            .O(N__16177),
            .I(N__16156));
    LocalMux I__3210 (
            .O(N__16174),
            .I(N__16156));
    InMux I__3209 (
            .O(N__16173),
            .I(N__16149));
    InMux I__3208 (
            .O(N__16172),
            .I(N__16149));
    InMux I__3207 (
            .O(N__16169),
            .I(N__16149));
    InMux I__3206 (
            .O(N__16168),
            .I(N__16146));
    InMux I__3205 (
            .O(N__16167),
            .I(N__16143));
    LocalMux I__3204 (
            .O(N__16164),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__3203 (
            .O(N__16161),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv4 I__3202 (
            .O(N__16156),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__3201 (
            .O(N__16149),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__3200 (
            .O(N__16146),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__3199 (
            .O(N__16143),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    CascadeMux I__3198 (
            .O(N__16130),
            .I(N__16125));
    CascadeMux I__3197 (
            .O(N__16129),
            .I(N__16122));
    InMux I__3196 (
            .O(N__16128),
            .I(N__16119));
    InMux I__3195 (
            .O(N__16125),
            .I(N__16112));
    InMux I__3194 (
            .O(N__16122),
            .I(N__16109));
    LocalMux I__3193 (
            .O(N__16119),
            .I(N__16106));
    InMux I__3192 (
            .O(N__16118),
            .I(N__16103));
    InMux I__3191 (
            .O(N__16117),
            .I(N__16098));
    InMux I__3190 (
            .O(N__16116),
            .I(N__16098));
    InMux I__3189 (
            .O(N__16115),
            .I(N__16095));
    LocalMux I__3188 (
            .O(N__16112),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    LocalMux I__3187 (
            .O(N__16109),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    Odrv4 I__3186 (
            .O(N__16106),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    LocalMux I__3185 (
            .O(N__16103),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    LocalMux I__3184 (
            .O(N__16098),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    LocalMux I__3183 (
            .O(N__16095),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    InMux I__3182 (
            .O(N__16082),
            .I(N__16077));
    InMux I__3181 (
            .O(N__16081),
            .I(N__16074));
    InMux I__3180 (
            .O(N__16080),
            .I(N__16069));
    LocalMux I__3179 (
            .O(N__16077),
            .I(N__16062));
    LocalMux I__3178 (
            .O(N__16074),
            .I(N__16059));
    InMux I__3177 (
            .O(N__16073),
            .I(N__16056));
    InMux I__3176 (
            .O(N__16072),
            .I(N__16053));
    LocalMux I__3175 (
            .O(N__16069),
            .I(N__16050));
    InMux I__3174 (
            .O(N__16068),
            .I(N__16043));
    InMux I__3173 (
            .O(N__16067),
            .I(N__16043));
    InMux I__3172 (
            .O(N__16066),
            .I(N__16043));
    InMux I__3171 (
            .O(N__16065),
            .I(N__16040));
    Span4Mux_h I__3170 (
            .O(N__16062),
            .I(N__16035));
    Span4Mux_h I__3169 (
            .O(N__16059),
            .I(N__16035));
    LocalMux I__3168 (
            .O(N__16056),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__3167 (
            .O(N__16053),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__3166 (
            .O(N__16050),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__3165 (
            .O(N__16043),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__3164 (
            .O(N__16040),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__3163 (
            .O(N__16035),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    InMux I__3162 (
            .O(N__16022),
            .I(N__16019));
    LocalMux I__3161 (
            .O(N__16019),
            .I(\POWERLED.un2_slp_s3n_2_0_o2_3_7 ));
    CascadeMux I__3160 (
            .O(N__16016),
            .I(\POWERLED.un2_slp_s3n_2_0_o2_3_8_cascade_ ));
    InMux I__3159 (
            .O(N__16013),
            .I(N__16010));
    LocalMux I__3158 (
            .O(N__16010),
            .I(N__16007));
    Span4Mux_v I__3157 (
            .O(N__16007),
            .I(N__16004));
    Odrv4 I__3156 (
            .O(N__16004),
            .I(\POWERLED.un2_slp_s3n_2_0_o2_3_6 ));
    InMux I__3155 (
            .O(N__16001),
            .I(N__15993));
    InMux I__3154 (
            .O(N__16000),
            .I(N__15990));
    InMux I__3153 (
            .O(N__15999),
            .I(N__15981));
    InMux I__3152 (
            .O(N__15998),
            .I(N__15981));
    InMux I__3151 (
            .O(N__15997),
            .I(N__15981));
    InMux I__3150 (
            .O(N__15996),
            .I(N__15981));
    LocalMux I__3149 (
            .O(N__15993),
            .I(N__15978));
    LocalMux I__3148 (
            .O(N__15990),
            .I(N__15975));
    LocalMux I__3147 (
            .O(N__15981),
            .I(N__15972));
    Span4Mux_h I__3146 (
            .O(N__15978),
            .I(N__15969));
    Span4Mux_h I__3145 (
            .O(N__15975),
            .I(N__15966));
    Span4Mux_h I__3144 (
            .O(N__15972),
            .I(N__15963));
    Odrv4 I__3143 (
            .O(N__15969),
            .I(\POWERLED.N_112 ));
    Odrv4 I__3142 (
            .O(N__15966),
            .I(\POWERLED.N_112 ));
    Odrv4 I__3141 (
            .O(N__15963),
            .I(\POWERLED.N_112 ));
    InMux I__3140 (
            .O(N__15956),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_3 ));
    InMux I__3139 (
            .O(N__15953),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_4 ));
    InMux I__3138 (
            .O(N__15950),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_5 ));
    InMux I__3137 (
            .O(N__15947),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_6 ));
    InMux I__3136 (
            .O(N__15944),
            .I(bfn_8_6_0_));
    InMux I__3135 (
            .O(N__15941),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_8 ));
    InMux I__3134 (
            .O(N__15938),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_9 ));
    InMux I__3133 (
            .O(N__15935),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_10 ));
    InMux I__3132 (
            .O(N__15932),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_11 ));
    InMux I__3131 (
            .O(N__15929),
            .I(N__15926));
    LocalMux I__3130 (
            .O(N__15926),
            .I(N__15923));
    Span4Mux_h I__3129 (
            .O(N__15923),
            .I(N__15920));
    Odrv4 I__3128 (
            .O(N__15920),
            .I(\HDA_STRAP.count_RNO_0Z0Z_6 ));
    CascadeMux I__3127 (
            .O(N__15917),
            .I(N__15911));
    CascadeMux I__3126 (
            .O(N__15916),
            .I(N__15908));
    CascadeMux I__3125 (
            .O(N__15915),
            .I(N__15905));
    InMux I__3124 (
            .O(N__15914),
            .I(N__15896));
    InMux I__3123 (
            .O(N__15911),
            .I(N__15891));
    InMux I__3122 (
            .O(N__15908),
            .I(N__15891));
    InMux I__3121 (
            .O(N__15905),
            .I(N__15886));
    InMux I__3120 (
            .O(N__15904),
            .I(N__15886));
    InMux I__3119 (
            .O(N__15903),
            .I(N__15883));
    InMux I__3118 (
            .O(N__15902),
            .I(N__15880));
    CascadeMux I__3117 (
            .O(N__15901),
            .I(N__15876));
    CascadeMux I__3116 (
            .O(N__15900),
            .I(N__15873));
    CascadeMux I__3115 (
            .O(N__15899),
            .I(N__15869));
    LocalMux I__3114 (
            .O(N__15896),
            .I(N__15864));
    LocalMux I__3113 (
            .O(N__15891),
            .I(N__15855));
    LocalMux I__3112 (
            .O(N__15886),
            .I(N__15855));
    LocalMux I__3111 (
            .O(N__15883),
            .I(N__15855));
    LocalMux I__3110 (
            .O(N__15880),
            .I(N__15855));
    InMux I__3109 (
            .O(N__15879),
            .I(N__15852));
    InMux I__3108 (
            .O(N__15876),
            .I(N__15849));
    InMux I__3107 (
            .O(N__15873),
            .I(N__15846));
    InMux I__3106 (
            .O(N__15872),
            .I(N__15839));
    InMux I__3105 (
            .O(N__15869),
            .I(N__15839));
    InMux I__3104 (
            .O(N__15868),
            .I(N__15839));
    InMux I__3103 (
            .O(N__15867),
            .I(N__15836));
    Span4Mux_v I__3102 (
            .O(N__15864),
            .I(N__15829));
    Span4Mux_v I__3101 (
            .O(N__15855),
            .I(N__15829));
    LocalMux I__3100 (
            .O(N__15852),
            .I(N__15829));
    LocalMux I__3099 (
            .O(N__15849),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    LocalMux I__3098 (
            .O(N__15846),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    LocalMux I__3097 (
            .O(N__15839),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    LocalMux I__3096 (
            .O(N__15836),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    Odrv4 I__3095 (
            .O(N__15829),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    CascadeMux I__3094 (
            .O(N__15818),
            .I(N__15815));
    InMux I__3093 (
            .O(N__15815),
            .I(N__15804));
    InMux I__3092 (
            .O(N__15814),
            .I(N__15795));
    InMux I__3091 (
            .O(N__15813),
            .I(N__15795));
    InMux I__3090 (
            .O(N__15812),
            .I(N__15795));
    InMux I__3089 (
            .O(N__15811),
            .I(N__15795));
    InMux I__3088 (
            .O(N__15810),
            .I(N__15792));
    InMux I__3087 (
            .O(N__15809),
            .I(N__15789));
    InMux I__3086 (
            .O(N__15808),
            .I(N__15782));
    InMux I__3085 (
            .O(N__15807),
            .I(N__15782));
    LocalMux I__3084 (
            .O(N__15804),
            .I(N__15779));
    LocalMux I__3083 (
            .O(N__15795),
            .I(N__15770));
    LocalMux I__3082 (
            .O(N__15792),
            .I(N__15770));
    LocalMux I__3081 (
            .O(N__15789),
            .I(N__15770));
    InMux I__3080 (
            .O(N__15788),
            .I(N__15767));
    InMux I__3079 (
            .O(N__15787),
            .I(N__15764));
    LocalMux I__3078 (
            .O(N__15782),
            .I(N__15761));
    Span4Mux_h I__3077 (
            .O(N__15779),
            .I(N__15758));
    InMux I__3076 (
            .O(N__15778),
            .I(N__15753));
    InMux I__3075 (
            .O(N__15777),
            .I(N__15753));
    Span4Mux_s2_v I__3074 (
            .O(N__15770),
            .I(N__15750));
    LocalMux I__3073 (
            .O(N__15767),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__3072 (
            .O(N__15764),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    Odrv4 I__3071 (
            .O(N__15761),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    Odrv4 I__3070 (
            .O(N__15758),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__3069 (
            .O(N__15753),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    Odrv4 I__3068 (
            .O(N__15750),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    InMux I__3067 (
            .O(N__15737),
            .I(N__15729));
    InMux I__3066 (
            .O(N__15736),
            .I(N__15729));
    InMux I__3065 (
            .O(N__15735),
            .I(N__15726));
    InMux I__3064 (
            .O(N__15734),
            .I(N__15718));
    LocalMux I__3063 (
            .O(N__15729),
            .I(N__15715));
    LocalMux I__3062 (
            .O(N__15726),
            .I(N__15712));
    InMux I__3061 (
            .O(N__15725),
            .I(N__15703));
    InMux I__3060 (
            .O(N__15724),
            .I(N__15703));
    InMux I__3059 (
            .O(N__15723),
            .I(N__15703));
    InMux I__3058 (
            .O(N__15722),
            .I(N__15703));
    InMux I__3057 (
            .O(N__15721),
            .I(N__15700));
    LocalMux I__3056 (
            .O(N__15718),
            .I(N__15693));
    Span4Mux_s1_v I__3055 (
            .O(N__15715),
            .I(N__15693));
    Span4Mux_v I__3054 (
            .O(N__15712),
            .I(N__15693));
    LocalMux I__3053 (
            .O(N__15703),
            .I(\HDA_STRAP.count_RNIB5IA5Z0Z_0 ));
    LocalMux I__3052 (
            .O(N__15700),
            .I(\HDA_STRAP.count_RNIB5IA5Z0Z_0 ));
    Odrv4 I__3051 (
            .O(N__15693),
            .I(\HDA_STRAP.count_RNIB5IA5Z0Z_0 ));
    InMux I__3050 (
            .O(N__15686),
            .I(N__15683));
    LocalMux I__3049 (
            .O(N__15683),
            .I(N__15680));
    Span4Mux_s1_v I__3048 (
            .O(N__15680),
            .I(N__15676));
    InMux I__3047 (
            .O(N__15679),
            .I(N__15673));
    Odrv4 I__3046 (
            .O(N__15676),
            .I(\HDA_STRAP.countZ0Z_6 ));
    LocalMux I__3045 (
            .O(N__15673),
            .I(\HDA_STRAP.countZ0Z_6 ));
    InMux I__3044 (
            .O(N__15668),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_0 ));
    InMux I__3043 (
            .O(N__15665),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_1 ));
    InMux I__3042 (
            .O(N__15662),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_2 ));
    InMux I__3041 (
            .O(N__15659),
            .I(N__15656));
    LocalMux I__3040 (
            .O(N__15656),
            .I(N__15653));
    Span4Mux_v I__3039 (
            .O(N__15653),
            .I(N__15640));
    InMux I__3038 (
            .O(N__15652),
            .I(N__15637));
    InMux I__3037 (
            .O(N__15651),
            .I(N__15632));
    InMux I__3036 (
            .O(N__15650),
            .I(N__15625));
    InMux I__3035 (
            .O(N__15649),
            .I(N__15625));
    InMux I__3034 (
            .O(N__15648),
            .I(N__15625));
    InMux I__3033 (
            .O(N__15647),
            .I(N__15622));
    InMux I__3032 (
            .O(N__15646),
            .I(N__15617));
    InMux I__3031 (
            .O(N__15645),
            .I(N__15617));
    InMux I__3030 (
            .O(N__15644),
            .I(N__15612));
    InMux I__3029 (
            .O(N__15643),
            .I(N__15612));
    Span4Mux_h I__3028 (
            .O(N__15640),
            .I(N__15607));
    LocalMux I__3027 (
            .O(N__15637),
            .I(N__15607));
    InMux I__3026 (
            .O(N__15636),
            .I(N__15602));
    InMux I__3025 (
            .O(N__15635),
            .I(N__15602));
    LocalMux I__3024 (
            .O(N__15632),
            .I(N__15597));
    LocalMux I__3023 (
            .O(N__15625),
            .I(N__15597));
    LocalMux I__3022 (
            .O(N__15622),
            .I(N_55));
    LocalMux I__3021 (
            .O(N__15617),
            .I(N_55));
    LocalMux I__3020 (
            .O(N__15612),
            .I(N_55));
    Odrv4 I__3019 (
            .O(N__15607),
            .I(N_55));
    LocalMux I__3018 (
            .O(N__15602),
            .I(N_55));
    Odrv4 I__3017 (
            .O(N__15597),
            .I(N_55));
    InMux I__3016 (
            .O(N__15584),
            .I(N__15576));
    InMux I__3015 (
            .O(N__15583),
            .I(N__15576));
    InMux I__3014 (
            .O(N__15582),
            .I(N__15571));
    InMux I__3013 (
            .O(N__15581),
            .I(N__15571));
    LocalMux I__3012 (
            .O(N__15576),
            .I(\VPP_VDDQ.N_238 ));
    LocalMux I__3011 (
            .O(N__15571),
            .I(\VPP_VDDQ.N_238 ));
    CascadeMux I__3010 (
            .O(N__15566),
            .I(\VPP_VDDQ.N_238_cascade_ ));
    CascadeMux I__3009 (
            .O(N__15563),
            .I(\VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_ ));
    InMux I__3008 (
            .O(N__15560),
            .I(N__15557));
    LocalMux I__3007 (
            .O(N__15557),
            .I(\VPP_VDDQ.G_127_0 ));
    InMux I__3006 (
            .O(N__15554),
            .I(N__15550));
    InMux I__3005 (
            .O(N__15553),
            .I(N__15547));
    LocalMux I__3004 (
            .O(N__15550),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    LocalMux I__3003 (
            .O(N__15547),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    InMux I__3002 (
            .O(N__15542),
            .I(N__15532));
    InMux I__3001 (
            .O(N__15541),
            .I(N__15532));
    InMux I__3000 (
            .O(N__15540),
            .I(N__15529));
    InMux I__2999 (
            .O(N__15539),
            .I(N__15526));
    InMux I__2998 (
            .O(N__15538),
            .I(N__15521));
    InMux I__2997 (
            .O(N__15537),
            .I(N__15521));
    LocalMux I__2996 (
            .O(N__15532),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    LocalMux I__2995 (
            .O(N__15529),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    LocalMux I__2994 (
            .O(N__15526),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    LocalMux I__2993 (
            .O(N__15521),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    InMux I__2992 (
            .O(N__15512),
            .I(N__15504));
    InMux I__2991 (
            .O(N__15511),
            .I(N__15501));
    InMux I__2990 (
            .O(N__15510),
            .I(N__15498));
    InMux I__2989 (
            .O(N__15509),
            .I(N__15491));
    InMux I__2988 (
            .O(N__15508),
            .I(N__15491));
    InMux I__2987 (
            .O(N__15507),
            .I(N__15491));
    LocalMux I__2986 (
            .O(N__15504),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    LocalMux I__2985 (
            .O(N__15501),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    LocalMux I__2984 (
            .O(N__15498),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    LocalMux I__2983 (
            .O(N__15491),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    CascadeMux I__2982 (
            .O(N__15482),
            .I(N__15479));
    InMux I__2981 (
            .O(N__15479),
            .I(N__15476));
    LocalMux I__2980 (
            .O(N__15476),
            .I(N__15472));
    InMux I__2979 (
            .O(N__15475),
            .I(N__15469));
    Odrv4 I__2978 (
            .O(N__15472),
            .I(\VPP_VDDQ.N_128 ));
    LocalMux I__2977 (
            .O(N__15469),
            .I(\VPP_VDDQ.N_128 ));
    CascadeMux I__2976 (
            .O(N__15464),
            .I(\VPP_VDDQ.N_154_cascade_ ));
    InMux I__2975 (
            .O(N__15461),
            .I(N__15458));
    LocalMux I__2974 (
            .O(N__15458),
            .I(\POWERLED.count_clk_1_sqmuxa_5_0_1 ));
    CascadeMux I__2973 (
            .O(N__15455),
            .I(\POWERLED.N_127_cascade_ ));
    InMux I__2972 (
            .O(N__15452),
            .I(N__15449));
    LocalMux I__2971 (
            .O(N__15449),
            .I(\POWERLED.count_clk_1_sqmuxa_5_0_0 ));
    CascadeMux I__2970 (
            .O(N__15446),
            .I(N__15442));
    CascadeMux I__2969 (
            .O(N__15445),
            .I(N__15439));
    InMux I__2968 (
            .O(N__15442),
            .I(N__15435));
    InMux I__2967 (
            .O(N__15439),
            .I(N__15432));
    InMux I__2966 (
            .O(N__15438),
            .I(N__15429));
    LocalMux I__2965 (
            .O(N__15435),
            .I(\POWERLED.N_88 ));
    LocalMux I__2964 (
            .O(N__15432),
            .I(\POWERLED.N_88 ));
    LocalMux I__2963 (
            .O(N__15429),
            .I(\POWERLED.N_88 ));
    CascadeMux I__2962 (
            .O(N__15422),
            .I(\POWERLED.dutycycle_3_sqmuxa_1_i_0_1_1_cascade_ ));
    InMux I__2961 (
            .O(N__15419),
            .I(N__15415));
    InMux I__2960 (
            .O(N__15418),
            .I(N__15412));
    LocalMux I__2959 (
            .O(N__15415),
            .I(\POWERLED.N_200_2 ));
    LocalMux I__2958 (
            .O(N__15412),
            .I(\POWERLED.N_200_2 ));
    InMux I__2957 (
            .O(N__15407),
            .I(N__15404));
    LocalMux I__2956 (
            .O(N__15404),
            .I(\POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_1 ));
    CascadeMux I__2955 (
            .O(N__15401),
            .I(\POWERLED.N_366_1_cascade_ ));
    InMux I__2954 (
            .O(N__15398),
            .I(N__15395));
    LocalMux I__2953 (
            .O(N__15395),
            .I(\POWERLED.N_251 ));
    CascadeMux I__2952 (
            .O(N__15392),
            .I(N__15389));
    InMux I__2951 (
            .O(N__15389),
            .I(N__15385));
    InMux I__2950 (
            .O(N__15388),
            .I(N__15382));
    LocalMux I__2949 (
            .O(N__15385),
            .I(N__15377));
    LocalMux I__2948 (
            .O(N__15382),
            .I(N__15377));
    Odrv12 I__2947 (
            .O(N__15377),
            .I(\POWERLED.dutycycle ));
    InMux I__2946 (
            .O(N__15374),
            .I(N__15369));
    InMux I__2945 (
            .O(N__15373),
            .I(N__15364));
    InMux I__2944 (
            .O(N__15372),
            .I(N__15364));
    LocalMux I__2943 (
            .O(N__15369),
            .I(\POWERLED.N_243 ));
    LocalMux I__2942 (
            .O(N__15364),
            .I(\POWERLED.N_243 ));
    InMux I__2941 (
            .O(N__15359),
            .I(N__15352));
    InMux I__2940 (
            .O(N__15358),
            .I(N__15347));
    InMux I__2939 (
            .O(N__15357),
            .I(N__15340));
    InMux I__2938 (
            .O(N__15356),
            .I(N__15340));
    InMux I__2937 (
            .O(N__15355),
            .I(N__15340));
    LocalMux I__2936 (
            .O(N__15352),
            .I(N__15337));
    InMux I__2935 (
            .O(N__15351),
            .I(N__15334));
    InMux I__2934 (
            .O(N__15350),
            .I(N__15331));
    LocalMux I__2933 (
            .O(N__15347),
            .I(N__15326));
    LocalMux I__2932 (
            .O(N__15340),
            .I(N__15326));
    Span4Mux_h I__2931 (
            .O(N__15337),
            .I(N__15323));
    LocalMux I__2930 (
            .O(N__15334),
            .I(N__15318));
    LocalMux I__2929 (
            .O(N__15331),
            .I(N__15318));
    Span4Mux_h I__2928 (
            .O(N__15326),
            .I(N__15315));
    Sp12to4 I__2927 (
            .O(N__15323),
            .I(N__15310));
    Span12Mux_s8_h I__2926 (
            .O(N__15318),
            .I(N__15310));
    Span4Mux_v I__2925 (
            .O(N__15315),
            .I(N__15307));
    Odrv12 I__2924 (
            .O(N__15310),
            .I(slp_s4n));
    Odrv4 I__2923 (
            .O(N__15307),
            .I(slp_s4n));
    InMux I__2922 (
            .O(N__15302),
            .I(N__15295));
    InMux I__2921 (
            .O(N__15301),
            .I(N__15290));
    InMux I__2920 (
            .O(N__15300),
            .I(N__15286));
    InMux I__2919 (
            .O(N__15299),
            .I(N__15283));
    InMux I__2918 (
            .O(N__15298),
            .I(N__15279));
    LocalMux I__2917 (
            .O(N__15295),
            .I(N__15276));
    InMux I__2916 (
            .O(N__15294),
            .I(N__15273));
    InMux I__2915 (
            .O(N__15293),
            .I(N__15270));
    LocalMux I__2914 (
            .O(N__15290),
            .I(N__15267));
    InMux I__2913 (
            .O(N__15289),
            .I(N__15264));
    LocalMux I__2912 (
            .O(N__15286),
            .I(N__15259));
    LocalMux I__2911 (
            .O(N__15283),
            .I(N__15259));
    InMux I__2910 (
            .O(N__15282),
            .I(N__15255));
    LocalMux I__2909 (
            .O(N__15279),
            .I(N__15252));
    Span4Mux_v I__2908 (
            .O(N__15276),
            .I(N__15241));
    LocalMux I__2907 (
            .O(N__15273),
            .I(N__15241));
    LocalMux I__2906 (
            .O(N__15270),
            .I(N__15241));
    Span4Mux_v I__2905 (
            .O(N__15267),
            .I(N__15241));
    LocalMux I__2904 (
            .O(N__15264),
            .I(N__15241));
    Span4Mux_h I__2903 (
            .O(N__15259),
            .I(N__15238));
    InMux I__2902 (
            .O(N__15258),
            .I(N__15235));
    LocalMux I__2901 (
            .O(N__15255),
            .I(\POWERLED.func_stateZ0Z_1 ));
    Odrv4 I__2900 (
            .O(N__15252),
            .I(\POWERLED.func_stateZ0Z_1 ));
    Odrv4 I__2899 (
            .O(N__15241),
            .I(\POWERLED.func_stateZ0Z_1 ));
    Odrv4 I__2898 (
            .O(N__15238),
            .I(\POWERLED.func_stateZ0Z_1 ));
    LocalMux I__2897 (
            .O(N__15235),
            .I(\POWERLED.func_stateZ0Z_1 ));
    CascadeMux I__2896 (
            .O(N__15224),
            .I(N__15217));
    CascadeMux I__2895 (
            .O(N__15223),
            .I(N__15213));
    InMux I__2894 (
            .O(N__15222),
            .I(N__15205));
    InMux I__2893 (
            .O(N__15221),
            .I(N__15202));
    InMux I__2892 (
            .O(N__15220),
            .I(N__15199));
    InMux I__2891 (
            .O(N__15217),
            .I(N__15190));
    InMux I__2890 (
            .O(N__15216),
            .I(N__15190));
    InMux I__2889 (
            .O(N__15213),
            .I(N__15190));
    InMux I__2888 (
            .O(N__15212),
            .I(N__15190));
    InMux I__2887 (
            .O(N__15211),
            .I(N__15185));
    InMux I__2886 (
            .O(N__15210),
            .I(N__15185));
    InMux I__2885 (
            .O(N__15209),
            .I(N__15180));
    InMux I__2884 (
            .O(N__15208),
            .I(N__15180));
    LocalMux I__2883 (
            .O(N__15205),
            .I(N__15171));
    LocalMux I__2882 (
            .O(N__15202),
            .I(N__15171));
    LocalMux I__2881 (
            .O(N__15199),
            .I(N__15171));
    LocalMux I__2880 (
            .O(N__15190),
            .I(N__15171));
    LocalMux I__2879 (
            .O(N__15185),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__2878 (
            .O(N__15180),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv4 I__2877 (
            .O(N__15171),
            .I(\POWERLED.func_stateZ0Z_0 ));
    InMux I__2876 (
            .O(N__15164),
            .I(N__15158));
    InMux I__2875 (
            .O(N__15163),
            .I(N__15152));
    InMux I__2874 (
            .O(N__15162),
            .I(N__15152));
    CascadeMux I__2873 (
            .O(N__15161),
            .I(N__15149));
    LocalMux I__2872 (
            .O(N__15158),
            .I(N__15144));
    InMux I__2871 (
            .O(N__15157),
            .I(N__15141));
    LocalMux I__2870 (
            .O(N__15152),
            .I(N__15138));
    InMux I__2869 (
            .O(N__15149),
            .I(N__15134));
    InMux I__2868 (
            .O(N__15148),
            .I(N__15131));
    InMux I__2867 (
            .O(N__15147),
            .I(N__15128));
    Span4Mux_v I__2866 (
            .O(N__15144),
            .I(N__15123));
    LocalMux I__2865 (
            .O(N__15141),
            .I(N__15123));
    Span4Mux_h I__2864 (
            .O(N__15138),
            .I(N__15120));
    InMux I__2863 (
            .O(N__15137),
            .I(N__15117));
    LocalMux I__2862 (
            .O(N__15134),
            .I(\POWERLED.count_off_RNIIKVR3Z0Z_10 ));
    LocalMux I__2861 (
            .O(N__15131),
            .I(\POWERLED.count_off_RNIIKVR3Z0Z_10 ));
    LocalMux I__2860 (
            .O(N__15128),
            .I(\POWERLED.count_off_RNIIKVR3Z0Z_10 ));
    Odrv4 I__2859 (
            .O(N__15123),
            .I(\POWERLED.count_off_RNIIKVR3Z0Z_10 ));
    Odrv4 I__2858 (
            .O(N__15120),
            .I(\POWERLED.count_off_RNIIKVR3Z0Z_10 ));
    LocalMux I__2857 (
            .O(N__15117),
            .I(\POWERLED.count_off_RNIIKVR3Z0Z_10 ));
    InMux I__2856 (
            .O(N__15104),
            .I(N__15101));
    LocalMux I__2855 (
            .O(N__15101),
            .I(\POWERLED.N_148 ));
    InMux I__2854 (
            .O(N__15098),
            .I(N__15094));
    CascadeMux I__2853 (
            .O(N__15097),
            .I(N__15087));
    LocalMux I__2852 (
            .O(N__15094),
            .I(N__15080));
    InMux I__2851 (
            .O(N__15093),
            .I(N__15077));
    InMux I__2850 (
            .O(N__15092),
            .I(N__15070));
    InMux I__2849 (
            .O(N__15091),
            .I(N__15070));
    InMux I__2848 (
            .O(N__15090),
            .I(N__15070));
    InMux I__2847 (
            .O(N__15087),
            .I(N__15065));
    InMux I__2846 (
            .O(N__15086),
            .I(N__15065));
    InMux I__2845 (
            .O(N__15085),
            .I(N__15058));
    InMux I__2844 (
            .O(N__15084),
            .I(N__15058));
    InMux I__2843 (
            .O(N__15083),
            .I(N__15058));
    Span4Mux_h I__2842 (
            .O(N__15080),
            .I(N__15050));
    LocalMux I__2841 (
            .O(N__15077),
            .I(N__15050));
    LocalMux I__2840 (
            .O(N__15070),
            .I(N__15050));
    LocalMux I__2839 (
            .O(N__15065),
            .I(N__15047));
    LocalMux I__2838 (
            .O(N__15058),
            .I(N__15044));
    InMux I__2837 (
            .O(N__15057),
            .I(N__15041));
    Span4Mux_v I__2836 (
            .O(N__15050),
            .I(N__15038));
    Span4Mux_v I__2835 (
            .O(N__15047),
            .I(N__15031));
    Span4Mux_v I__2834 (
            .O(N__15044),
            .I(N__15031));
    LocalMux I__2833 (
            .O(N__15041),
            .I(N__15031));
    Span4Mux_h I__2832 (
            .O(N__15038),
            .I(N__15026));
    Span4Mux_h I__2831 (
            .O(N__15031),
            .I(N__15026));
    Odrv4 I__2830 (
            .O(N__15026),
            .I(slp_s3n));
    IoInMux I__2829 (
            .O(N__15023),
            .I(N__15020));
    LocalMux I__2828 (
            .O(N__15020),
            .I(N__15016));
    InMux I__2827 (
            .O(N__15019),
            .I(N__15013));
    Span4Mux_s2_h I__2826 (
            .O(N__15016),
            .I(N__15007));
    LocalMux I__2825 (
            .O(N__15013),
            .I(N__15004));
    InMux I__2824 (
            .O(N__15012),
            .I(N__14999));
    InMux I__2823 (
            .O(N__15011),
            .I(N__14994));
    InMux I__2822 (
            .O(N__15010),
            .I(N__14994));
    Span4Mux_h I__2821 (
            .O(N__15007),
            .I(N__14991));
    Span4Mux_v I__2820 (
            .O(N__15004),
            .I(N__14988));
    InMux I__2819 (
            .O(N__15003),
            .I(N__14983));
    InMux I__2818 (
            .O(N__15002),
            .I(N__14983));
    LocalMux I__2817 (
            .O(N__14999),
            .I(N__14978));
    LocalMux I__2816 (
            .O(N__14994),
            .I(N__14978));
    Odrv4 I__2815 (
            .O(N__14991),
            .I(vccst_en));
    Odrv4 I__2814 (
            .O(N__14988),
            .I(vccst_en));
    LocalMux I__2813 (
            .O(N__14983),
            .I(vccst_en));
    Odrv4 I__2812 (
            .O(N__14978),
            .I(vccst_en));
    IoInMux I__2811 (
            .O(N__14969),
            .I(N__14966));
    LocalMux I__2810 (
            .O(N__14966),
            .I(N__14963));
    Odrv12 I__2809 (
            .O(N__14963),
            .I(vpp_en));
    CascadeMux I__2808 (
            .O(N__14960),
            .I(\POWERLED.N_203_cascade_ ));
    CascadeMux I__2807 (
            .O(N__14957),
            .I(\POWERLED.N_251_cascade_ ));
    InMux I__2806 (
            .O(N__14954),
            .I(N__14951));
    LocalMux I__2805 (
            .O(N__14951),
            .I(\POWERLED.un2_slp_s3n_2_0_1_0 ));
    InMux I__2804 (
            .O(N__14948),
            .I(N__14945));
    LocalMux I__2803 (
            .O(N__14945),
            .I(\POWERLED.count_clk_139_tz_0 ));
    CascadeMux I__2802 (
            .O(N__14942),
            .I(\POWERLED.un2_slp_s3n_2_0_cascade_ ));
    InMux I__2801 (
            .O(N__14939),
            .I(N__14936));
    LocalMux I__2800 (
            .O(N__14936),
            .I(\POWERLED.N_246 ));
    InMux I__2799 (
            .O(N__14933),
            .I(N__14930));
    LocalMux I__2798 (
            .O(N__14930),
            .I(N__14927));
    Span4Mux_h I__2797 (
            .O(N__14927),
            .I(N__14923));
    InMux I__2796 (
            .O(N__14926),
            .I(N__14920));
    Odrv4 I__2795 (
            .O(N__14923),
            .I(\POWERLED.N_205 ));
    LocalMux I__2794 (
            .O(N__14920),
            .I(\POWERLED.N_205 ));
    CascadeMux I__2793 (
            .O(N__14915),
            .I(\POWERLED.un2_slp_s3n_2_0_a6_3_0_cascade_ ));
    InMux I__2792 (
            .O(N__14912),
            .I(N__14909));
    LocalMux I__2791 (
            .O(N__14909),
            .I(\POWERLED.un2_slp_s3n_2_0_1 ));
    InMux I__2790 (
            .O(N__14906),
            .I(N__14903));
    LocalMux I__2789 (
            .O(N__14903),
            .I(N__14898));
    CascadeMux I__2788 (
            .O(N__14902),
            .I(N__14894));
    InMux I__2787 (
            .O(N__14901),
            .I(N__14891));
    Span4Mux_h I__2786 (
            .O(N__14898),
            .I(N__14888));
    InMux I__2785 (
            .O(N__14897),
            .I(N__14885));
    InMux I__2784 (
            .O(N__14894),
            .I(N__14882));
    LocalMux I__2783 (
            .O(N__14891),
            .I(N__14879));
    Odrv4 I__2782 (
            .O(N__14888),
            .I(\POWERLED.N_127 ));
    LocalMux I__2781 (
            .O(N__14885),
            .I(\POWERLED.N_127 ));
    LocalMux I__2780 (
            .O(N__14882),
            .I(\POWERLED.N_127 ));
    Odrv4 I__2779 (
            .O(N__14879),
            .I(\POWERLED.N_127 ));
    InMux I__2778 (
            .O(N__14870),
            .I(\POWERLED.dutycycle_cry_9 ));
    InMux I__2777 (
            .O(N__14867),
            .I(\POWERLED.dutycycle_cry_10 ));
    InMux I__2776 (
            .O(N__14864),
            .I(\POWERLED.dutycycle_cry_11 ));
    InMux I__2775 (
            .O(N__14861),
            .I(\POWERLED.dutycycle_cry_12 ));
    InMux I__2774 (
            .O(N__14858),
            .I(\POWERLED.dutycycle_cry_13 ));
    CascadeMux I__2773 (
            .O(N__14855),
            .I(N__14845));
    CascadeMux I__2772 (
            .O(N__14854),
            .I(N__14841));
    CascadeMux I__2771 (
            .O(N__14853),
            .I(N__14837));
    CascadeMux I__2770 (
            .O(N__14852),
            .I(N__14833));
    CascadeMux I__2769 (
            .O(N__14851),
            .I(N__14829));
    CascadeMux I__2768 (
            .O(N__14850),
            .I(N__14825));
    CascadeMux I__2767 (
            .O(N__14849),
            .I(N__14821));
    InMux I__2766 (
            .O(N__14848),
            .I(N__14805));
    InMux I__2765 (
            .O(N__14845),
            .I(N__14805));
    InMux I__2764 (
            .O(N__14844),
            .I(N__14805));
    InMux I__2763 (
            .O(N__14841),
            .I(N__14805));
    InMux I__2762 (
            .O(N__14840),
            .I(N__14805));
    InMux I__2761 (
            .O(N__14837),
            .I(N__14805));
    InMux I__2760 (
            .O(N__14836),
            .I(N__14805));
    InMux I__2759 (
            .O(N__14833),
            .I(N__14787));
    InMux I__2758 (
            .O(N__14832),
            .I(N__14787));
    InMux I__2757 (
            .O(N__14829),
            .I(N__14787));
    InMux I__2756 (
            .O(N__14828),
            .I(N__14787));
    InMux I__2755 (
            .O(N__14825),
            .I(N__14787));
    InMux I__2754 (
            .O(N__14824),
            .I(N__14787));
    InMux I__2753 (
            .O(N__14821),
            .I(N__14787));
    InMux I__2752 (
            .O(N__14820),
            .I(N__14787));
    LocalMux I__2751 (
            .O(N__14805),
            .I(N__14784));
    InMux I__2750 (
            .O(N__14804),
            .I(N__14781));
    LocalMux I__2749 (
            .O(N__14787),
            .I(N__14778));
    Span4Mux_h I__2748 (
            .O(N__14784),
            .I(N__14775));
    LocalMux I__2747 (
            .O(N__14781),
            .I(\POWERLED.N_177 ));
    Odrv4 I__2746 (
            .O(N__14778),
            .I(\POWERLED.N_177 ));
    Odrv4 I__2745 (
            .O(N__14775),
            .I(\POWERLED.N_177 ));
    InMux I__2744 (
            .O(N__14768),
            .I(bfn_7_9_0_));
    CascadeMux I__2743 (
            .O(N__14765),
            .I(\POWERLED.N_246_cascade_ ));
    InMux I__2742 (
            .O(N__14762),
            .I(N__14759));
    LocalMux I__2741 (
            .O(N__14759),
            .I(\POWERLED.N_203_4 ));
    CascadeMux I__2740 (
            .O(N__14756),
            .I(\POWERLED.N_203_4_cascade_ ));
    InMux I__2739 (
            .O(N__14753),
            .I(N__14748));
    InMux I__2738 (
            .O(N__14752),
            .I(N__14745));
    CascadeMux I__2737 (
            .O(N__14751),
            .I(N__14742));
    LocalMux I__2736 (
            .O(N__14748),
            .I(N__14737));
    LocalMux I__2735 (
            .O(N__14745),
            .I(N__14733));
    InMux I__2734 (
            .O(N__14742),
            .I(N__14730));
    CascadeMux I__2733 (
            .O(N__14741),
            .I(N__14727));
    CascadeMux I__2732 (
            .O(N__14740),
            .I(N__14723));
    Span4Mux_v I__2731 (
            .O(N__14737),
            .I(N__14719));
    InMux I__2730 (
            .O(N__14736),
            .I(N__14716));
    Span4Mux_v I__2729 (
            .O(N__14733),
            .I(N__14713));
    LocalMux I__2728 (
            .O(N__14730),
            .I(N__14710));
    InMux I__2727 (
            .O(N__14727),
            .I(N__14707));
    InMux I__2726 (
            .O(N__14726),
            .I(N__14704));
    InMux I__2725 (
            .O(N__14723),
            .I(N__14701));
    InMux I__2724 (
            .O(N__14722),
            .I(N__14698));
    Span4Mux_v I__2723 (
            .O(N__14719),
            .I(N__14693));
    LocalMux I__2722 (
            .O(N__14716),
            .I(N__14693));
    Span4Mux_h I__2721 (
            .O(N__14713),
            .I(N__14688));
    Span4Mux_h I__2720 (
            .O(N__14710),
            .I(N__14688));
    LocalMux I__2719 (
            .O(N__14707),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__2718 (
            .O(N__14704),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__2717 (
            .O(N__14701),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__2716 (
            .O(N__14698),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__2715 (
            .O(N__14693),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__2714 (
            .O(N__14688),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    InMux I__2713 (
            .O(N__14675),
            .I(N__14672));
    LocalMux I__2712 (
            .O(N__14672),
            .I(\POWERLED.dutycycle_s_2 ));
    InMux I__2711 (
            .O(N__14669),
            .I(\POWERLED.dutycycle_cry_1 ));
    InMux I__2710 (
            .O(N__14666),
            .I(N__14662));
    CascadeMux I__2709 (
            .O(N__14665),
            .I(N__14659));
    LocalMux I__2708 (
            .O(N__14662),
            .I(N__14655));
    InMux I__2707 (
            .O(N__14659),
            .I(N__14651));
    InMux I__2706 (
            .O(N__14658),
            .I(N__14648));
    Span4Mux_v I__2705 (
            .O(N__14655),
            .I(N__14641));
    InMux I__2704 (
            .O(N__14654),
            .I(N__14638));
    LocalMux I__2703 (
            .O(N__14651),
            .I(N__14633));
    LocalMux I__2702 (
            .O(N__14648),
            .I(N__14633));
    InMux I__2701 (
            .O(N__14647),
            .I(N__14630));
    InMux I__2700 (
            .O(N__14646),
            .I(N__14625));
    InMux I__2699 (
            .O(N__14645),
            .I(N__14625));
    InMux I__2698 (
            .O(N__14644),
            .I(N__14622));
    Odrv4 I__2697 (
            .O(N__14641),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__2696 (
            .O(N__14638),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__2695 (
            .O(N__14633),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__2694 (
            .O(N__14630),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__2693 (
            .O(N__14625),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__2692 (
            .O(N__14622),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    InMux I__2691 (
            .O(N__14609),
            .I(\POWERLED.dutycycle_cry_2 ));
    InMux I__2690 (
            .O(N__14606),
            .I(N__14598));
    InMux I__2689 (
            .O(N__14605),
            .I(N__14593));
    InMux I__2688 (
            .O(N__14604),
            .I(N__14593));
    CascadeMux I__2687 (
            .O(N__14603),
            .I(N__14590));
    InMux I__2686 (
            .O(N__14602),
            .I(N__14587));
    InMux I__2685 (
            .O(N__14601),
            .I(N__14582));
    LocalMux I__2684 (
            .O(N__14598),
            .I(N__14579));
    LocalMux I__2683 (
            .O(N__14593),
            .I(N__14576));
    InMux I__2682 (
            .O(N__14590),
            .I(N__14573));
    LocalMux I__2681 (
            .O(N__14587),
            .I(N__14570));
    InMux I__2680 (
            .O(N__14586),
            .I(N__14565));
    InMux I__2679 (
            .O(N__14585),
            .I(N__14565));
    LocalMux I__2678 (
            .O(N__14582),
            .I(N__14560));
    Span4Mux_h I__2677 (
            .O(N__14579),
            .I(N__14560));
    Span4Mux_h I__2676 (
            .O(N__14576),
            .I(N__14557));
    LocalMux I__2675 (
            .O(N__14573),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__2674 (
            .O(N__14570),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__2673 (
            .O(N__14565),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__2672 (
            .O(N__14560),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__2671 (
            .O(N__14557),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    InMux I__2670 (
            .O(N__14546),
            .I(\POWERLED.dutycycle_cry_3 ));
    CascadeMux I__2669 (
            .O(N__14543),
            .I(N__14539));
    InMux I__2668 (
            .O(N__14542),
            .I(N__14536));
    InMux I__2667 (
            .O(N__14539),
            .I(N__14533));
    LocalMux I__2666 (
            .O(N__14536),
            .I(N__14527));
    LocalMux I__2665 (
            .O(N__14533),
            .I(N__14524));
    CascadeMux I__2664 (
            .O(N__14532),
            .I(N__14520));
    CascadeMux I__2663 (
            .O(N__14531),
            .I(N__14517));
    InMux I__2662 (
            .O(N__14530),
            .I(N__14514));
    Span4Mux_v I__2661 (
            .O(N__14527),
            .I(N__14511));
    Span4Mux_h I__2660 (
            .O(N__14524),
            .I(N__14508));
    InMux I__2659 (
            .O(N__14523),
            .I(N__14505));
    InMux I__2658 (
            .O(N__14520),
            .I(N__14500));
    InMux I__2657 (
            .O(N__14517),
            .I(N__14500));
    LocalMux I__2656 (
            .O(N__14514),
            .I(N__14497));
    Odrv4 I__2655 (
            .O(N__14511),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__2654 (
            .O(N__14508),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__2653 (
            .O(N__14505),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__2652 (
            .O(N__14500),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__2651 (
            .O(N__14497),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    InMux I__2650 (
            .O(N__14486),
            .I(N__14482));
    InMux I__2649 (
            .O(N__14485),
            .I(N__14479));
    LocalMux I__2648 (
            .O(N__14482),
            .I(N__14476));
    LocalMux I__2647 (
            .O(N__14479),
            .I(N__14473));
    Span4Mux_h I__2646 (
            .O(N__14476),
            .I(N__14470));
    Span4Mux_h I__2645 (
            .O(N__14473),
            .I(N__14467));
    Odrv4 I__2644 (
            .O(N__14470),
            .I(\POWERLED.dutycycle_s_5 ));
    Odrv4 I__2643 (
            .O(N__14467),
            .I(\POWERLED.dutycycle_s_5 ));
    InMux I__2642 (
            .O(N__14462),
            .I(\POWERLED.dutycycle_cry_4 ));
    CascadeMux I__2641 (
            .O(N__14459),
            .I(N__14456));
    InMux I__2640 (
            .O(N__14456),
            .I(N__14451));
    InMux I__2639 (
            .O(N__14455),
            .I(N__14446));
    InMux I__2638 (
            .O(N__14454),
            .I(N__14446));
    LocalMux I__2637 (
            .O(N__14451),
            .I(N__14437));
    LocalMux I__2636 (
            .O(N__14446),
            .I(N__14437));
    InMux I__2635 (
            .O(N__14445),
            .I(N__14434));
    InMux I__2634 (
            .O(N__14444),
            .I(N__14427));
    InMux I__2633 (
            .O(N__14443),
            .I(N__14427));
    InMux I__2632 (
            .O(N__14442),
            .I(N__14427));
    Span4Mux_v I__2631 (
            .O(N__14437),
            .I(N__14424));
    LocalMux I__2630 (
            .O(N__14434),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__2629 (
            .O(N__14427),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__2628 (
            .O(N__14424),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    InMux I__2627 (
            .O(N__14417),
            .I(N__14411));
    InMux I__2626 (
            .O(N__14416),
            .I(N__14411));
    LocalMux I__2625 (
            .O(N__14411),
            .I(N__14408));
    Span4Mux_h I__2624 (
            .O(N__14408),
            .I(N__14405));
    Odrv4 I__2623 (
            .O(N__14405),
            .I(\POWERLED.dutycycle_s_6 ));
    InMux I__2622 (
            .O(N__14402),
            .I(\POWERLED.dutycycle_cry_5 ));
    CascadeMux I__2621 (
            .O(N__14399),
            .I(N__14389));
    InMux I__2620 (
            .O(N__14398),
            .I(N__14386));
    CascadeMux I__2619 (
            .O(N__14397),
            .I(N__14382));
    CascadeMux I__2618 (
            .O(N__14396),
            .I(N__14379));
    InMux I__2617 (
            .O(N__14395),
            .I(N__14374));
    InMux I__2616 (
            .O(N__14394),
            .I(N__14374));
    InMux I__2615 (
            .O(N__14393),
            .I(N__14370));
    InMux I__2614 (
            .O(N__14392),
            .I(N__14365));
    InMux I__2613 (
            .O(N__14389),
            .I(N__14365));
    LocalMux I__2612 (
            .O(N__14386),
            .I(N__14362));
    InMux I__2611 (
            .O(N__14385),
            .I(N__14357));
    InMux I__2610 (
            .O(N__14382),
            .I(N__14357));
    InMux I__2609 (
            .O(N__14379),
            .I(N__14354));
    LocalMux I__2608 (
            .O(N__14374),
            .I(N__14351));
    InMux I__2607 (
            .O(N__14373),
            .I(N__14348));
    LocalMux I__2606 (
            .O(N__14370),
            .I(N__14343));
    LocalMux I__2605 (
            .O(N__14365),
            .I(N__14343));
    Span4Mux_v I__2604 (
            .O(N__14362),
            .I(N__14338));
    LocalMux I__2603 (
            .O(N__14357),
            .I(N__14338));
    LocalMux I__2602 (
            .O(N__14354),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__2601 (
            .O(N__14351),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__2600 (
            .O(N__14348),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__2599 (
            .O(N__14343),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__2598 (
            .O(N__14338),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    InMux I__2597 (
            .O(N__14327),
            .I(bfn_7_8_0_));
    InMux I__2596 (
            .O(N__14324),
            .I(\POWERLED.dutycycle_cry_7 ));
    InMux I__2595 (
            .O(N__14321),
            .I(\POWERLED.dutycycle_cry_8 ));
    CascadeMux I__2594 (
            .O(N__14318),
            .I(\POWERLED.un1_dutycycle_1_39_0_cascade_ ));
    CascadeMux I__2593 (
            .O(N__14315),
            .I(N__14312));
    InMux I__2592 (
            .O(N__14312),
            .I(N__14309));
    LocalMux I__2591 (
            .O(N__14309),
            .I(\POWERLED.dutycycle_RNI34C41Z0Z_8 ));
    CascadeMux I__2590 (
            .O(N__14306),
            .I(N__14301));
    InMux I__2589 (
            .O(N__14305),
            .I(N__14296));
    InMux I__2588 (
            .O(N__14304),
            .I(N__14296));
    InMux I__2587 (
            .O(N__14301),
            .I(N__14293));
    LocalMux I__2586 (
            .O(N__14296),
            .I(N__14290));
    LocalMux I__2585 (
            .O(N__14293),
            .I(N__14285));
    Span4Mux_h I__2584 (
            .O(N__14290),
            .I(N__14285));
    Span4Mux_v I__2583 (
            .O(N__14285),
            .I(N__14282));
    Odrv4 I__2582 (
            .O(N__14282),
            .I(\POWERLED.N_117 ));
    InMux I__2581 (
            .O(N__14279),
            .I(N__14275));
    CascadeMux I__2580 (
            .O(N__14278),
            .I(N__14272));
    LocalMux I__2579 (
            .O(N__14275),
            .I(N__14269));
    InMux I__2578 (
            .O(N__14272),
            .I(N__14266));
    Odrv12 I__2577 (
            .O(N__14269),
            .I(\POWERLED.dutycycle_fast_RNIVCSKZ0Z_5 ));
    LocalMux I__2576 (
            .O(N__14266),
            .I(\POWERLED.dutycycle_fast_RNIVCSKZ0Z_5 ));
    InMux I__2575 (
            .O(N__14261),
            .I(N__14258));
    LocalMux I__2574 (
            .O(N__14258),
            .I(\POWERLED.dutycycle_RNIK4I81Z0Z_6 ));
    CascadeMux I__2573 (
            .O(N__14255),
            .I(N__14252));
    InMux I__2572 (
            .O(N__14252),
            .I(N__14249));
    LocalMux I__2571 (
            .O(N__14249),
            .I(N__14246));
    Odrv4 I__2570 (
            .O(N__14246),
            .I(\POWERLED.dutycycle_lm_0_1_2 ));
    CascadeMux I__2569 (
            .O(N__14243),
            .I(N__14240));
    InMux I__2568 (
            .O(N__14240),
            .I(N__14236));
    InMux I__2567 (
            .O(N__14239),
            .I(N__14233));
    LocalMux I__2566 (
            .O(N__14236),
            .I(N__14230));
    LocalMux I__2565 (
            .O(N__14233),
            .I(\POWERLED.dutycycle_fast_RNI2GSKZ0Z_6 ));
    Odrv4 I__2564 (
            .O(N__14230),
            .I(\POWERLED.dutycycle_fast_RNI2GSKZ0Z_6 ));
    InMux I__2563 (
            .O(N__14225),
            .I(N__14222));
    LocalMux I__2562 (
            .O(N__14222),
            .I(\POWERLED.dutycycle_RNIQAI81Z0Z_4 ));
    InMux I__2561 (
            .O(N__14219),
            .I(N__14216));
    LocalMux I__2560 (
            .O(N__14216),
            .I(\POWERLED.dutycycle_RNIOQLJZ0Z_4 ));
    CascadeMux I__2559 (
            .O(N__14213),
            .I(N__14210));
    InMux I__2558 (
            .O(N__14210),
            .I(N__14206));
    InMux I__2557 (
            .O(N__14209),
            .I(N__14203));
    LocalMux I__2556 (
            .O(N__14206),
            .I(N__14200));
    LocalMux I__2555 (
            .O(N__14203),
            .I(N__14197));
    Span4Mux_v I__2554 (
            .O(N__14200),
            .I(N__14191));
    Span4Mux_h I__2553 (
            .O(N__14197),
            .I(N__14188));
    InMux I__2552 (
            .O(N__14196),
            .I(N__14185));
    InMux I__2551 (
            .O(N__14195),
            .I(N__14182));
    CascadeMux I__2550 (
            .O(N__14194),
            .I(N__14179));
    Span4Mux_h I__2549 (
            .O(N__14191),
            .I(N__14174));
    Span4Mux_v I__2548 (
            .O(N__14188),
            .I(N__14169));
    LocalMux I__2547 (
            .O(N__14185),
            .I(N__14169));
    LocalMux I__2546 (
            .O(N__14182),
            .I(N__14166));
    InMux I__2545 (
            .O(N__14179),
            .I(N__14163));
    InMux I__2544 (
            .O(N__14178),
            .I(N__14160));
    InMux I__2543 (
            .O(N__14177),
            .I(N__14157));
    Odrv4 I__2542 (
            .O(N__14174),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__2541 (
            .O(N__14169),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__2540 (
            .O(N__14166),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__2539 (
            .O(N__14163),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__2538 (
            .O(N__14160),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__2537 (
            .O(N__14157),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    InMux I__2536 (
            .O(N__14144),
            .I(N__14141));
    LocalMux I__2535 (
            .O(N__14141),
            .I(N__14138));
    Span4Mux_v I__2534 (
            .O(N__14138),
            .I(N__14135));
    Odrv4 I__2533 (
            .O(N__14135),
            .I(\POWERLED.dutycycle_s_0 ));
    InMux I__2532 (
            .O(N__14132),
            .I(\POWERLED.dutycycle_cry_c_0_THRU_CO ));
    InMux I__2531 (
            .O(N__14129),
            .I(N__14124));
    InMux I__2530 (
            .O(N__14128),
            .I(N__14120));
    InMux I__2529 (
            .O(N__14127),
            .I(N__14116));
    LocalMux I__2528 (
            .O(N__14124),
            .I(N__14113));
    InMux I__2527 (
            .O(N__14123),
            .I(N__14107));
    LocalMux I__2526 (
            .O(N__14120),
            .I(N__14104));
    InMux I__2525 (
            .O(N__14119),
            .I(N__14101));
    LocalMux I__2524 (
            .O(N__14116),
            .I(N__14098));
    Span4Mux_v I__2523 (
            .O(N__14113),
            .I(N__14095));
    CascadeMux I__2522 (
            .O(N__14112),
            .I(N__14092));
    CascadeMux I__2521 (
            .O(N__14111),
            .I(N__14089));
    CascadeMux I__2520 (
            .O(N__14110),
            .I(N__14085));
    LocalMux I__2519 (
            .O(N__14107),
            .I(N__14082));
    Span4Mux_v I__2518 (
            .O(N__14104),
            .I(N__14077));
    LocalMux I__2517 (
            .O(N__14101),
            .I(N__14077));
    Span4Mux_v I__2516 (
            .O(N__14098),
            .I(N__14072));
    Span4Mux_h I__2515 (
            .O(N__14095),
            .I(N__14072));
    InMux I__2514 (
            .O(N__14092),
            .I(N__14067));
    InMux I__2513 (
            .O(N__14089),
            .I(N__14067));
    InMux I__2512 (
            .O(N__14088),
            .I(N__14062));
    InMux I__2511 (
            .O(N__14085),
            .I(N__14062));
    Odrv12 I__2510 (
            .O(N__14082),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__2509 (
            .O(N__14077),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__2508 (
            .O(N__14072),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__2507 (
            .O(N__14067),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__2506 (
            .O(N__14062),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    InMux I__2505 (
            .O(N__14051),
            .I(N__14048));
    LocalMux I__2504 (
            .O(N__14048),
            .I(N__14045));
    Span4Mux_h I__2503 (
            .O(N__14045),
            .I(N__14042));
    Odrv4 I__2502 (
            .O(N__14042),
            .I(\POWERLED.dutycycle_s_1 ));
    InMux I__2501 (
            .O(N__14039),
            .I(\POWERLED.dutycycle_cry_0 ));
    CascadeMux I__2500 (
            .O(N__14036),
            .I(N__14033));
    InMux I__2499 (
            .O(N__14033),
            .I(N__14030));
    LocalMux I__2498 (
            .O(N__14030),
            .I(N__14027));
    Odrv12 I__2497 (
            .O(N__14027),
            .I(\HDA_STRAP.curr_state_RNO_0Z0Z_2 ));
    CascadeMux I__2496 (
            .O(N__14024),
            .I(N__14021));
    InMux I__2495 (
            .O(N__14021),
            .I(N__14018));
    LocalMux I__2494 (
            .O(N__14018),
            .I(\HDA_STRAP.count_RNO_0Z0Z_10 ));
    CascadeMux I__2493 (
            .O(N__14015),
            .I(N__14012));
    InMux I__2492 (
            .O(N__14012),
            .I(N__14008));
    InMux I__2491 (
            .O(N__14011),
            .I(N__14005));
    LocalMux I__2490 (
            .O(N__14008),
            .I(\HDA_STRAP.countZ0Z_10 ));
    LocalMux I__2489 (
            .O(N__14005),
            .I(\HDA_STRAP.countZ0Z_10 ));
    InMux I__2488 (
            .O(N__14000),
            .I(N__13997));
    LocalMux I__2487 (
            .O(N__13997),
            .I(\HDA_STRAP.count_RNO_0Z0Z_16 ));
    InMux I__2486 (
            .O(N__13994),
            .I(N__13990));
    InMux I__2485 (
            .O(N__13993),
            .I(N__13987));
    LocalMux I__2484 (
            .O(N__13990),
            .I(\HDA_STRAP.countZ0Z_16 ));
    LocalMux I__2483 (
            .O(N__13987),
            .I(\HDA_STRAP.countZ0Z_16 ));
    InMux I__2482 (
            .O(N__13982),
            .I(N__13979));
    LocalMux I__2481 (
            .O(N__13979),
            .I(\HDA_STRAP.count_RNO_0Z0Z_17 ));
    InMux I__2480 (
            .O(N__13976),
            .I(N__13972));
    InMux I__2479 (
            .O(N__13975),
            .I(N__13969));
    LocalMux I__2478 (
            .O(N__13972),
            .I(\HDA_STRAP.countZ0Z_17 ));
    LocalMux I__2477 (
            .O(N__13969),
            .I(\HDA_STRAP.countZ0Z_17 ));
    InMux I__2476 (
            .O(N__13964),
            .I(N__13961));
    LocalMux I__2475 (
            .O(N__13961),
            .I(\HDA_STRAP.count_RNO_0Z0Z_8 ));
    InMux I__2474 (
            .O(N__13958),
            .I(N__13954));
    InMux I__2473 (
            .O(N__13957),
            .I(N__13951));
    LocalMux I__2472 (
            .O(N__13954),
            .I(\HDA_STRAP.countZ0Z_8 ));
    LocalMux I__2471 (
            .O(N__13951),
            .I(\HDA_STRAP.countZ0Z_8 ));
    CascadeMux I__2470 (
            .O(N__13946),
            .I(N__13943));
    InMux I__2469 (
            .O(N__13943),
            .I(N__13940));
    LocalMux I__2468 (
            .O(N__13940),
            .I(\POWERLED.dutycycle_RNI31MG_0Z0Z_12 ));
    CascadeMux I__2467 (
            .O(N__13937),
            .I(N__13934));
    InMux I__2466 (
            .O(N__13934),
            .I(N__13931));
    LocalMux I__2465 (
            .O(N__13931),
            .I(\POWERLED.dutycycle_RNI31MGZ0Z_12 ));
    CascadeMux I__2464 (
            .O(N__13928),
            .I(N__13924));
    InMux I__2463 (
            .O(N__13927),
            .I(N__13921));
    InMux I__2462 (
            .O(N__13924),
            .I(N__13918));
    LocalMux I__2461 (
            .O(N__13921),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ));
    LocalMux I__2460 (
            .O(N__13918),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ));
    InMux I__2459 (
            .O(N__13913),
            .I(N__13909));
    InMux I__2458 (
            .O(N__13912),
            .I(N__13906));
    LocalMux I__2457 (
            .O(N__13909),
            .I(\HDA_STRAP.countZ0Z_2 ));
    LocalMux I__2456 (
            .O(N__13906),
            .I(\HDA_STRAP.countZ0Z_2 ));
    InMux I__2455 (
            .O(N__13901),
            .I(N__13897));
    InMux I__2454 (
            .O(N__13900),
            .I(N__13894));
    LocalMux I__2453 (
            .O(N__13897),
            .I(\HDA_STRAP.countZ0Z_1 ));
    LocalMux I__2452 (
            .O(N__13894),
            .I(\HDA_STRAP.countZ0Z_1 ));
    CascadeMux I__2451 (
            .O(N__13889),
            .I(N__13885));
    InMux I__2450 (
            .O(N__13888),
            .I(N__13882));
    InMux I__2449 (
            .O(N__13885),
            .I(N__13879));
    LocalMux I__2448 (
            .O(N__13882),
            .I(\HDA_STRAP.countZ0Z_3 ));
    LocalMux I__2447 (
            .O(N__13879),
            .I(\HDA_STRAP.countZ0Z_3 ));
    InMux I__2446 (
            .O(N__13874),
            .I(N__13870));
    InMux I__2445 (
            .O(N__13873),
            .I(N__13867));
    LocalMux I__2444 (
            .O(N__13870),
            .I(N__13862));
    LocalMux I__2443 (
            .O(N__13867),
            .I(N__13862));
    Odrv4 I__2442 (
            .O(N__13862),
            .I(\HDA_STRAP.countZ0Z_0 ));
    InMux I__2441 (
            .O(N__13859),
            .I(N__13855));
    InMux I__2440 (
            .O(N__13858),
            .I(N__13852));
    LocalMux I__2439 (
            .O(N__13855),
            .I(\HDA_STRAP.countZ0Z_14 ));
    LocalMux I__2438 (
            .O(N__13852),
            .I(\HDA_STRAP.countZ0Z_14 ));
    CascadeMux I__2437 (
            .O(N__13847),
            .I(N__13843));
    InMux I__2436 (
            .O(N__13846),
            .I(N__13840));
    InMux I__2435 (
            .O(N__13843),
            .I(N__13837));
    LocalMux I__2434 (
            .O(N__13840),
            .I(\HDA_STRAP.countZ0Z_15 ));
    LocalMux I__2433 (
            .O(N__13837),
            .I(\HDA_STRAP.countZ0Z_15 ));
    InMux I__2432 (
            .O(N__13832),
            .I(N__13828));
    InMux I__2431 (
            .O(N__13831),
            .I(N__13825));
    LocalMux I__2430 (
            .O(N__13828),
            .I(\HDA_STRAP.countZ0Z_12 ));
    LocalMux I__2429 (
            .O(N__13825),
            .I(\HDA_STRAP.countZ0Z_12 ));
    CascadeMux I__2428 (
            .O(N__13820),
            .I(\HDA_STRAP.un4_count_9_cascade_ ));
    InMux I__2427 (
            .O(N__13817),
            .I(N__13813));
    InMux I__2426 (
            .O(N__13816),
            .I(N__13810));
    LocalMux I__2425 (
            .O(N__13813),
            .I(\HDA_STRAP.countZ0Z_13 ));
    LocalMux I__2424 (
            .O(N__13810),
            .I(\HDA_STRAP.countZ0Z_13 ));
    InMux I__2423 (
            .O(N__13805),
            .I(N__13801));
    InMux I__2422 (
            .O(N__13804),
            .I(N__13798));
    LocalMux I__2421 (
            .O(N__13801),
            .I(\HDA_STRAP.countZ0Z_7 ));
    LocalMux I__2420 (
            .O(N__13798),
            .I(\HDA_STRAP.countZ0Z_7 ));
    InMux I__2419 (
            .O(N__13793),
            .I(N__13789));
    InMux I__2418 (
            .O(N__13792),
            .I(N__13786));
    LocalMux I__2417 (
            .O(N__13789),
            .I(\HDA_STRAP.countZ0Z_5 ));
    LocalMux I__2416 (
            .O(N__13786),
            .I(\HDA_STRAP.countZ0Z_5 ));
    CascadeMux I__2415 (
            .O(N__13781),
            .I(N__13777));
    InMux I__2414 (
            .O(N__13780),
            .I(N__13774));
    InMux I__2413 (
            .O(N__13777),
            .I(N__13771));
    LocalMux I__2412 (
            .O(N__13774),
            .I(\HDA_STRAP.countZ0Z_9 ));
    LocalMux I__2411 (
            .O(N__13771),
            .I(\HDA_STRAP.countZ0Z_9 ));
    InMux I__2410 (
            .O(N__13766),
            .I(N__13762));
    InMux I__2409 (
            .O(N__13765),
            .I(N__13759));
    LocalMux I__2408 (
            .O(N__13762),
            .I(\HDA_STRAP.countZ0Z_4 ));
    LocalMux I__2407 (
            .O(N__13759),
            .I(\HDA_STRAP.countZ0Z_4 ));
    InMux I__2406 (
            .O(N__13754),
            .I(N__13750));
    InMux I__2405 (
            .O(N__13753),
            .I(N__13747));
    LocalMux I__2404 (
            .O(N__13750),
            .I(N__13744));
    LocalMux I__2403 (
            .O(N__13747),
            .I(\HDA_STRAP.countZ0Z_11 ));
    Odrv4 I__2402 (
            .O(N__13744),
            .I(\HDA_STRAP.countZ0Z_11 ));
    InMux I__2401 (
            .O(N__13739),
            .I(N__13736));
    LocalMux I__2400 (
            .O(N__13736),
            .I(\HDA_STRAP.un4_count_12 ));
    InMux I__2399 (
            .O(N__13733),
            .I(N__13730));
    LocalMux I__2398 (
            .O(N__13730),
            .I(\HDA_STRAP.un4_count_11 ));
    CascadeMux I__2397 (
            .O(N__13727),
            .I(\HDA_STRAP.un4_count_10_cascade_ ));
    InMux I__2396 (
            .O(N__13724),
            .I(N__13721));
    LocalMux I__2395 (
            .O(N__13721),
            .I(\HDA_STRAP.un4_count_13 ));
    CascadeMux I__2394 (
            .O(N__13718),
            .I(\HDA_STRAP.count_RNIB5IA5Z0Z_0_cascade_ ));
    CascadeMux I__2393 (
            .O(N__13715),
            .I(\POWERLED.N_208_cascade_ ));
    InMux I__2392 (
            .O(N__13712),
            .I(N__13709));
    LocalMux I__2391 (
            .O(N__13709),
            .I(\POWERLED.func_state_ns_i_0_1_1 ));
    InMux I__2390 (
            .O(N__13706),
            .I(N__13703));
    LocalMux I__2389 (
            .O(N__13703),
            .I(N__13695));
    InMux I__2388 (
            .O(N__13702),
            .I(N__13690));
    InMux I__2387 (
            .O(N__13701),
            .I(N__13690));
    CascadeMux I__2386 (
            .O(N__13700),
            .I(N__13687));
    CascadeMux I__2385 (
            .O(N__13699),
            .I(N__13684));
    InMux I__2384 (
            .O(N__13698),
            .I(N__13680));
    Span4Mux_h I__2383 (
            .O(N__13695),
            .I(N__13677));
    LocalMux I__2382 (
            .O(N__13690),
            .I(N__13674));
    InMux I__2381 (
            .O(N__13687),
            .I(N__13667));
    InMux I__2380 (
            .O(N__13684),
            .I(N__13667));
    InMux I__2379 (
            .O(N__13683),
            .I(N__13667));
    LocalMux I__2378 (
            .O(N__13680),
            .I(\POWERLED.N_222 ));
    Odrv4 I__2377 (
            .O(N__13677),
            .I(\POWERLED.N_222 ));
    Odrv4 I__2376 (
            .O(N__13674),
            .I(\POWERLED.N_222 ));
    LocalMux I__2375 (
            .O(N__13667),
            .I(\POWERLED.N_222 ));
    CascadeMux I__2374 (
            .O(N__13658),
            .I(\POWERLED.N_222_cascade_ ));
    InMux I__2373 (
            .O(N__13655),
            .I(N__13649));
    InMux I__2372 (
            .O(N__13654),
            .I(N__13649));
    LocalMux I__2371 (
            .O(N__13649),
            .I(\POWERLED.N_228 ));
    CascadeMux I__2370 (
            .O(N__13646),
            .I(\POWERLED.N_211_cascade_ ));
    CascadeMux I__2369 (
            .O(N__13643),
            .I(N__13640));
    InMux I__2368 (
            .O(N__13640),
            .I(N__13637));
    LocalMux I__2367 (
            .O(N__13637),
            .I(\POWERLED.func_state_ns_i_0_0_1 ));
    InMux I__2366 (
            .O(N__13634),
            .I(N__13631));
    LocalMux I__2365 (
            .O(N__13631),
            .I(\POWERLED.N_179 ));
    InMux I__2364 (
            .O(N__13628),
            .I(N__13625));
    LocalMux I__2363 (
            .O(N__13625),
            .I(\POWERLED.N_178 ));
    CascadeMux I__2362 (
            .O(N__13622),
            .I(N__13619));
    InMux I__2361 (
            .O(N__13619),
            .I(N__13616));
    LocalMux I__2360 (
            .O(N__13616),
            .I(N__13613));
    Odrv4 I__2359 (
            .O(N__13613),
            .I(\POWERLED.N_180 ));
    InMux I__2358 (
            .O(N__13610),
            .I(N__13607));
    LocalMux I__2357 (
            .O(N__13607),
            .I(N__13603));
    InMux I__2356 (
            .O(N__13606),
            .I(N__13600));
    Odrv4 I__2355 (
            .O(N__13603),
            .I(\POWERLED.N_250 ));
    LocalMux I__2354 (
            .O(N__13600),
            .I(\POWERLED.N_250 ));
    CascadeMux I__2353 (
            .O(N__13595),
            .I(N__13590));
    CascadeMux I__2352 (
            .O(N__13594),
            .I(N__13587));
    CascadeMux I__2351 (
            .O(N__13593),
            .I(N__13583));
    InMux I__2350 (
            .O(N__13590),
            .I(N__13576));
    InMux I__2349 (
            .O(N__13587),
            .I(N__13576));
    InMux I__2348 (
            .O(N__13586),
            .I(N__13576));
    InMux I__2347 (
            .O(N__13583),
            .I(N__13573));
    LocalMux I__2346 (
            .O(N__13576),
            .I(N__13570));
    LocalMux I__2345 (
            .O(N__13573),
            .I(N__13567));
    Span4Mux_h I__2344 (
            .O(N__13570),
            .I(N__13564));
    Span4Mux_v I__2343 (
            .O(N__13567),
            .I(N__13561));
    Odrv4 I__2342 (
            .O(N__13564),
            .I(\POWERLED.N_213 ));
    Odrv4 I__2341 (
            .O(N__13561),
            .I(\POWERLED.N_213 ));
    InMux I__2340 (
            .O(N__13556),
            .I(N__13550));
    InMux I__2339 (
            .O(N__13555),
            .I(N__13550));
    LocalMux I__2338 (
            .O(N__13550),
            .I(N__13545));
    InMux I__2337 (
            .O(N__13549),
            .I(N__13540));
    InMux I__2336 (
            .O(N__13548),
            .I(N__13540));
    Span4Mux_v I__2335 (
            .O(N__13545),
            .I(N__13535));
    LocalMux I__2334 (
            .O(N__13540),
            .I(N__13535));
    Odrv4 I__2333 (
            .O(N__13535),
            .I(\POWERLED.N_234 ));
    CascadeMux I__2332 (
            .O(N__13532),
            .I(\POWERLED.N_218_cascade_ ));
    InMux I__2331 (
            .O(N__13529),
            .I(N__13525));
    InMux I__2330 (
            .O(N__13528),
            .I(N__13522));
    LocalMux I__2329 (
            .O(N__13525),
            .I(N__13518));
    LocalMux I__2328 (
            .O(N__13522),
            .I(N__13514));
    InMux I__2327 (
            .O(N__13521),
            .I(N__13511));
    Span4Mux_v I__2326 (
            .O(N__13518),
            .I(N__13508));
    InMux I__2325 (
            .O(N__13517),
            .I(N__13505));
    Odrv4 I__2324 (
            .O(N__13514),
            .I(\POWERLED.N_248 ));
    LocalMux I__2323 (
            .O(N__13511),
            .I(\POWERLED.N_248 ));
    Odrv4 I__2322 (
            .O(N__13508),
            .I(\POWERLED.N_248 ));
    LocalMux I__2321 (
            .O(N__13505),
            .I(\POWERLED.N_248 ));
    CascadeMux I__2320 (
            .O(N__13496),
            .I(\POWERLED.N_88_cascade_ ));
    CascadeMux I__2319 (
            .O(N__13493),
            .I(N__13490));
    InMux I__2318 (
            .O(N__13490),
            .I(N__13487));
    LocalMux I__2317 (
            .O(N__13487),
            .I(N__13484));
    Odrv12 I__2316 (
            .O(N__13484),
            .I(\POWERLED.dutycycle_RNIC8C11Z0Z_15 ));
    InMux I__2315 (
            .O(N__13481),
            .I(N__13478));
    LocalMux I__2314 (
            .O(N__13478),
            .I(N__13475));
    Span4Mux_h I__2313 (
            .O(N__13475),
            .I(N__13472));
    Odrv4 I__2312 (
            .O(N__13472),
            .I(\POWERLED.dutycycle_RNI73C11Z0Z_15 ));
    CascadeMux I__2311 (
            .O(N__13469),
            .I(N__13466));
    InMux I__2310 (
            .O(N__13466),
            .I(N__13463));
    LocalMux I__2309 (
            .O(N__13463),
            .I(\POWERLED.N_368_0_i_i_a6_0 ));
    CascadeMux I__2308 (
            .O(N__13460),
            .I(\POWERLED.N_207_cascade_ ));
    CascadeMux I__2307 (
            .O(N__13457),
            .I(N__13453));
    InMux I__2306 (
            .O(N__13456),
            .I(N__13450));
    InMux I__2305 (
            .O(N__13453),
            .I(N__13447));
    LocalMux I__2304 (
            .O(N__13450),
            .I(\POWERLED.N_48 ));
    LocalMux I__2303 (
            .O(N__13447),
            .I(\POWERLED.N_48 ));
    CascadeMux I__2302 (
            .O(N__13442),
            .I(N__13439));
    InMux I__2301 (
            .O(N__13439),
            .I(N__13436));
    LocalMux I__2300 (
            .O(N__13436),
            .I(\POWERLED.N_149 ));
    CascadeMux I__2299 (
            .O(N__13433),
            .I(\POWERLED.N_149_cascade_ ));
    InMux I__2298 (
            .O(N__13430),
            .I(N__13426));
    CascadeMux I__2297 (
            .O(N__13429),
            .I(N__13423));
    LocalMux I__2296 (
            .O(N__13426),
            .I(N__13418));
    InMux I__2295 (
            .O(N__13423),
            .I(N__13411));
    InMux I__2294 (
            .O(N__13422),
            .I(N__13411));
    InMux I__2293 (
            .O(N__13421),
            .I(N__13411));
    Span4Mux_v I__2292 (
            .O(N__13418),
            .I(N__13406));
    LocalMux I__2291 (
            .O(N__13411),
            .I(N__13406));
    Span4Mux_h I__2290 (
            .O(N__13406),
            .I(N__13403));
    Odrv4 I__2289 (
            .O(N__13403),
            .I(\POWERLED.N_214 ));
    CascadeMux I__2288 (
            .O(N__13400),
            .I(N__13397));
    InMux I__2287 (
            .O(N__13397),
            .I(N__13394));
    LocalMux I__2286 (
            .O(N__13394),
            .I(N__13391));
    Odrv4 I__2285 (
            .O(N__13391),
            .I(\POWERLED.dutycycle_RNI2V0PZ0Z_10 ));
    CascadeMux I__2284 (
            .O(N__13388),
            .I(\POWERLED.dutycycle_RNI2V0PZ0Z_10_cascade_ ));
    InMux I__2283 (
            .O(N__13385),
            .I(N__13382));
    LocalMux I__2282 (
            .O(N__13382),
            .I(N__13379));
    Odrv4 I__2281 (
            .O(N__13379),
            .I(\POWERLED.dutycycle_RNI712I1Z0Z_15 ));
    InMux I__2280 (
            .O(N__13376),
            .I(N__13373));
    LocalMux I__2279 (
            .O(N__13373),
            .I(N__13370));
    Odrv4 I__2278 (
            .O(N__13370),
            .I(\POWERLED.dutycycle_RNIQ09G1Z0Z_10 ));
    InMux I__2277 (
            .O(N__13367),
            .I(N__13363));
    InMux I__2276 (
            .O(N__13366),
            .I(N__13360));
    LocalMux I__2275 (
            .O(N__13363),
            .I(\POWERLED.count_offZ0Z_3 ));
    LocalMux I__2274 (
            .O(N__13360),
            .I(\POWERLED.count_offZ0Z_3 ));
    InMux I__2273 (
            .O(N__13355),
            .I(N__13351));
    InMux I__2272 (
            .O(N__13354),
            .I(N__13348));
    LocalMux I__2271 (
            .O(N__13351),
            .I(N__13345));
    LocalMux I__2270 (
            .O(N__13348),
            .I(\POWERLED.count_offZ0Z_7 ));
    Odrv4 I__2269 (
            .O(N__13345),
            .I(\POWERLED.count_offZ0Z_7 ));
    CascadeMux I__2268 (
            .O(N__13340),
            .I(N__13336));
    InMux I__2267 (
            .O(N__13339),
            .I(N__13333));
    InMux I__2266 (
            .O(N__13336),
            .I(N__13330));
    LocalMux I__2265 (
            .O(N__13333),
            .I(\POWERLED.count_offZ0Z_4 ));
    LocalMux I__2264 (
            .O(N__13330),
            .I(\POWERLED.count_offZ0Z_4 ));
    InMux I__2263 (
            .O(N__13325),
            .I(N__13321));
    InMux I__2262 (
            .O(N__13324),
            .I(N__13318));
    LocalMux I__2261 (
            .O(N__13321),
            .I(\POWERLED.count_offZ0Z_2 ));
    LocalMux I__2260 (
            .O(N__13318),
            .I(\POWERLED.count_offZ0Z_2 ));
    InMux I__2259 (
            .O(N__13313),
            .I(N__13310));
    LocalMux I__2258 (
            .O(N__13310),
            .I(N__13307));
    Odrv4 I__2257 (
            .O(N__13307),
            .I(\POWERLED.func_state_ns_0_a2_8_0 ));
    CascadeMux I__2256 (
            .O(N__13304),
            .I(\POWERLED.un1_dutycycle_1_44_0_cascade_ ));
    CascadeMux I__2255 (
            .O(N__13301),
            .I(N__13298));
    InMux I__2254 (
            .O(N__13298),
            .I(N__13295));
    LocalMux I__2253 (
            .O(N__13295),
            .I(N__13292));
    Odrv4 I__2252 (
            .O(N__13292),
            .I(\POWERLED.dutycycle_RNIF3561Z0Z_9 ));
    InMux I__2251 (
            .O(N__13289),
            .I(N__13286));
    LocalMux I__2250 (
            .O(N__13286),
            .I(\POWERLED.dutycycle_RNIE4FLZ0Z_9 ));
    InMux I__2249 (
            .O(N__13283),
            .I(N__13280));
    LocalMux I__2248 (
            .O(N__13280),
            .I(\POWERLED.dutycycle_RNI53MGZ0Z_14 ));
    InMux I__2247 (
            .O(N__13277),
            .I(N__13274));
    LocalMux I__2246 (
            .O(N__13274),
            .I(\POWERLED.dutycycle_RNI84C11Z0Z_14 ));
    InMux I__2245 (
            .O(N__13271),
            .I(N__13268));
    LocalMux I__2244 (
            .O(N__13268),
            .I(\POWERLED.dutycycle_RNIB1FLZ0Z_8 ));
    CascadeMux I__2243 (
            .O(N__13265),
            .I(N__13262));
    InMux I__2242 (
            .O(N__13262),
            .I(N__13259));
    LocalMux I__2241 (
            .O(N__13259),
            .I(\POWERLED.dutycycle_RNI75MGZ0Z_15 ));
    CascadeMux I__2240 (
            .O(N__13256),
            .I(\POWERLED.un1_dutycycle_1_34_0_cascade_ ));
    CascadeMux I__2239 (
            .O(N__13253),
            .I(\POWERLED.un1_dutycycle_1_axb_8_cascade_ ));
    InMux I__2238 (
            .O(N__13250),
            .I(N__13247));
    LocalMux I__2237 (
            .O(N__13247),
            .I(N__13243));
    InMux I__2236 (
            .O(N__13246),
            .I(N__13240));
    Odrv4 I__2235 (
            .O(N__13243),
            .I(\POWERLED.dutycycle_fast_RNILMLMZ0Z_6 ));
    LocalMux I__2234 (
            .O(N__13240),
            .I(\POWERLED.dutycycle_fast_RNILMLMZ0Z_6 ));
    CascadeMux I__2233 (
            .O(N__13235),
            .I(N__13232));
    InMux I__2232 (
            .O(N__13232),
            .I(N__13229));
    LocalMux I__2231 (
            .O(N__13229),
            .I(N__13226));
    Odrv4 I__2230 (
            .O(N__13226),
            .I(\POWERLED.dutycycle_RNIJL1R1Z0Z_6 ));
    CascadeMux I__2229 (
            .O(N__13223),
            .I(N__13219));
    InMux I__2228 (
            .O(N__13222),
            .I(N__13215));
    InMux I__2227 (
            .O(N__13219),
            .I(N__13212));
    InMux I__2226 (
            .O(N__13218),
            .I(N__13209));
    LocalMux I__2225 (
            .O(N__13215),
            .I(\POWERLED.dutycycle_fastZ0Z_6 ));
    LocalMux I__2224 (
            .O(N__13212),
            .I(\POWERLED.dutycycle_fastZ0Z_6 ));
    LocalMux I__2223 (
            .O(N__13209),
            .I(\POWERLED.dutycycle_fastZ0Z_6 ));
    CascadeMux I__2222 (
            .O(N__13202),
            .I(N__13199));
    InMux I__2221 (
            .O(N__13199),
            .I(N__13195));
    InMux I__2220 (
            .O(N__13198),
            .I(N__13192));
    LocalMux I__2219 (
            .O(N__13195),
            .I(N__13189));
    LocalMux I__2218 (
            .O(N__13192),
            .I(\POWERLED.dutycycle_fast_RNIBPSKZ0Z_6 ));
    Odrv4 I__2217 (
            .O(N__13189),
            .I(\POWERLED.dutycycle_fast_RNIBPSKZ0Z_6 ));
    InMux I__2216 (
            .O(N__13184),
            .I(N__13180));
    InMux I__2215 (
            .O(N__13183),
            .I(N__13177));
    LocalMux I__2214 (
            .O(N__13180),
            .I(N__13174));
    LocalMux I__2213 (
            .O(N__13177),
            .I(N__13171));
    Span4Mux_h I__2212 (
            .O(N__13174),
            .I(N__13168));
    Odrv4 I__2211 (
            .O(N__13171),
            .I(\POWERLED.mult1_un68_sum ));
    Odrv4 I__2210 (
            .O(N__13168),
            .I(\POWERLED.mult1_un68_sum ));
    InMux I__2209 (
            .O(N__13163),
            .I(\POWERLED.un1_dutycycle_1_cry_10 ));
    InMux I__2208 (
            .O(N__13160),
            .I(N__13157));
    LocalMux I__2207 (
            .O(N__13157),
            .I(N__13153));
    InMux I__2206 (
            .O(N__13156),
            .I(N__13150));
    Span4Mux_v I__2205 (
            .O(N__13153),
            .I(N__13147));
    LocalMux I__2204 (
            .O(N__13150),
            .I(\POWERLED.mult1_un61_sum ));
    Odrv4 I__2203 (
            .O(N__13147),
            .I(\POWERLED.mult1_un61_sum ));
    InMux I__2202 (
            .O(N__13142),
            .I(\POWERLED.un1_dutycycle_1_cry_11 ));
    InMux I__2201 (
            .O(N__13139),
            .I(N__13136));
    LocalMux I__2200 (
            .O(N__13136),
            .I(N__13132));
    InMux I__2199 (
            .O(N__13135),
            .I(N__13129));
    Span4Mux_h I__2198 (
            .O(N__13132),
            .I(N__13126));
    LocalMux I__2197 (
            .O(N__13129),
            .I(\POWERLED.mult1_un54_sum ));
    Odrv4 I__2196 (
            .O(N__13126),
            .I(\POWERLED.mult1_un54_sum ));
    InMux I__2195 (
            .O(N__13121),
            .I(\POWERLED.un1_dutycycle_1_cry_12 ));
    CascadeMux I__2194 (
            .O(N__13118),
            .I(N__13115));
    InMux I__2193 (
            .O(N__13115),
            .I(N__13111));
    InMux I__2192 (
            .O(N__13114),
            .I(N__13108));
    LocalMux I__2191 (
            .O(N__13111),
            .I(N__13105));
    LocalMux I__2190 (
            .O(N__13108),
            .I(\POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1 ));
    Odrv4 I__2189 (
            .O(N__13105),
            .I(\POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1 ));
    InMux I__2188 (
            .O(N__13100),
            .I(\POWERLED.un1_dutycycle_1_cry_13 ));
    CascadeMux I__2187 (
            .O(N__13097),
            .I(N__13092));
    CascadeMux I__2186 (
            .O(N__13096),
            .I(N__13089));
    InMux I__2185 (
            .O(N__13095),
            .I(N__13079));
    InMux I__2184 (
            .O(N__13092),
            .I(N__13079));
    InMux I__2183 (
            .O(N__13089),
            .I(N__13079));
    InMux I__2182 (
            .O(N__13088),
            .I(N__13079));
    LocalMux I__2181 (
            .O(N__13079),
            .I(\POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1 ));
    InMux I__2180 (
            .O(N__13076),
            .I(\POWERLED.un1_dutycycle_1_cry_14 ));
    CascadeMux I__2179 (
            .O(N__13073),
            .I(N__13070));
    InMux I__2178 (
            .O(N__13070),
            .I(N__13061));
    InMux I__2177 (
            .O(N__13069),
            .I(N__13061));
    InMux I__2176 (
            .O(N__13068),
            .I(N__13061));
    LocalMux I__2175 (
            .O(N__13061),
            .I(\POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71 ));
    InMux I__2174 (
            .O(N__13058),
            .I(bfn_6_7_0_));
    InMux I__2173 (
            .O(N__13055),
            .I(\POWERLED.CO2 ));
    InMux I__2172 (
            .O(N__13052),
            .I(N__13046));
    InMux I__2171 (
            .O(N__13051),
            .I(N__13046));
    LocalMux I__2170 (
            .O(N__13046),
            .I(\POWERLED.CO2_THRU_CO ));
    InMux I__2169 (
            .O(N__13043),
            .I(N__13038));
    InMux I__2168 (
            .O(N__13042),
            .I(N__13035));
    InMux I__2167 (
            .O(N__13041),
            .I(N__13032));
    LocalMux I__2166 (
            .O(N__13038),
            .I(\POWERLED.dutycycle_fastZ0Z_5 ));
    LocalMux I__2165 (
            .O(N__13035),
            .I(\POWERLED.dutycycle_fastZ0Z_5 ));
    LocalMux I__2164 (
            .O(N__13032),
            .I(\POWERLED.dutycycle_fastZ0Z_5 ));
    CascadeMux I__2163 (
            .O(N__13025),
            .I(N__13022));
    InMux I__2162 (
            .O(N__13022),
            .I(N__13018));
    InMux I__2161 (
            .O(N__13021),
            .I(N__13015));
    LocalMux I__2160 (
            .O(N__13018),
            .I(N__13012));
    LocalMux I__2159 (
            .O(N__13015),
            .I(\POWERLED.dutycycle_fast_RNI8MSKZ0Z_5 ));
    Odrv4 I__2158 (
            .O(N__13012),
            .I(\POWERLED.dutycycle_fast_RNI8MSKZ0Z_5 ));
    InMux I__2157 (
            .O(N__13007),
            .I(N__13003));
    InMux I__2156 (
            .O(N__13006),
            .I(N__13000));
    LocalMux I__2155 (
            .O(N__13003),
            .I(N__12997));
    LocalMux I__2154 (
            .O(N__13000),
            .I(N__12992));
    Span4Mux_h I__2153 (
            .O(N__12997),
            .I(N__12992));
    Span4Mux_v I__2152 (
            .O(N__12992),
            .I(N__12989));
    Odrv4 I__2151 (
            .O(N__12989),
            .I(\POWERLED.mult1_un124_sum ));
    InMux I__2150 (
            .O(N__12986),
            .I(\POWERLED.un1_dutycycle_1_cry_2 ));
    InMux I__2149 (
            .O(N__12983),
            .I(N__12980));
    LocalMux I__2148 (
            .O(N__12980),
            .I(N__12976));
    InMux I__2147 (
            .O(N__12979),
            .I(N__12973));
    Span4Mux_h I__2146 (
            .O(N__12976),
            .I(N__12968));
    LocalMux I__2145 (
            .O(N__12973),
            .I(N__12968));
    Span4Mux_v I__2144 (
            .O(N__12968),
            .I(N__12965));
    Odrv4 I__2143 (
            .O(N__12965),
            .I(\POWERLED.mult1_un117_sum ));
    InMux I__2142 (
            .O(N__12962),
            .I(\POWERLED.un1_dutycycle_1_cry_3 ));
    CascadeMux I__2141 (
            .O(N__12959),
            .I(N__12956));
    InMux I__2140 (
            .O(N__12956),
            .I(N__12953));
    LocalMux I__2139 (
            .O(N__12953),
            .I(\POWERLED.dutycycle_RNIEJ021Z0Z_4 ));
    InMux I__2138 (
            .O(N__12950),
            .I(N__12946));
    InMux I__2137 (
            .O(N__12949),
            .I(N__12943));
    LocalMux I__2136 (
            .O(N__12946),
            .I(N__12940));
    LocalMux I__2135 (
            .O(N__12943),
            .I(N__12935));
    Span4Mux_s1_h I__2134 (
            .O(N__12940),
            .I(N__12935));
    Span4Mux_h I__2133 (
            .O(N__12935),
            .I(N__12932));
    Odrv4 I__2132 (
            .O(N__12932),
            .I(\POWERLED.mult1_un110_sum ));
    InMux I__2131 (
            .O(N__12929),
            .I(\POWERLED.un1_dutycycle_1_cry_4 ));
    InMux I__2130 (
            .O(N__12926),
            .I(N__12923));
    LocalMux I__2129 (
            .O(N__12923),
            .I(N__12920));
    Odrv4 I__2128 (
            .O(N__12920),
            .I(\POWERLED.dutycycle_RNI6NI81Z0Z_5 ));
    InMux I__2127 (
            .O(N__12917),
            .I(N__12913));
    InMux I__2126 (
            .O(N__12916),
            .I(N__12910));
    LocalMux I__2125 (
            .O(N__12913),
            .I(N__12907));
    LocalMux I__2124 (
            .O(N__12910),
            .I(N__12904));
    Span4Mux_v I__2123 (
            .O(N__12907),
            .I(N__12899));
    Span4Mux_s1_h I__2122 (
            .O(N__12904),
            .I(N__12899));
    Span4Mux_h I__2121 (
            .O(N__12899),
            .I(N__12896));
    Odrv4 I__2120 (
            .O(N__12896),
            .I(\POWERLED.mult1_un103_sum ));
    InMux I__2119 (
            .O(N__12893),
            .I(\POWERLED.un1_dutycycle_1_cry_5 ));
    InMux I__2118 (
            .O(N__12890),
            .I(N__12887));
    LocalMux I__2117 (
            .O(N__12887),
            .I(N__12884));
    Span4Mux_h I__2116 (
            .O(N__12884),
            .I(N__12881));
    Odrv4 I__2115 (
            .O(N__12881),
            .I(\POWERLED.dutycycle_RNIJNBA1Z0Z_6 ));
    InMux I__2114 (
            .O(N__12878),
            .I(N__12875));
    LocalMux I__2113 (
            .O(N__12875),
            .I(N__12871));
    InMux I__2112 (
            .O(N__12874),
            .I(N__12868));
    Span4Mux_v I__2111 (
            .O(N__12871),
            .I(N__12865));
    LocalMux I__2110 (
            .O(N__12868),
            .I(N__12862));
    Span4Mux_v I__2109 (
            .O(N__12865),
            .I(N__12857));
    Span4Mux_s1_h I__2108 (
            .O(N__12862),
            .I(N__12857));
    Span4Mux_h I__2107 (
            .O(N__12857),
            .I(N__12854));
    Odrv4 I__2106 (
            .O(N__12854),
            .I(\POWERLED.mult1_un96_sum ));
    InMux I__2105 (
            .O(N__12851),
            .I(\POWERLED.un1_dutycycle_1_cry_6 ));
    InMux I__2104 (
            .O(N__12848),
            .I(N__12844));
    InMux I__2103 (
            .O(N__12847),
            .I(N__12841));
    LocalMux I__2102 (
            .O(N__12844),
            .I(N__12838));
    LocalMux I__2101 (
            .O(N__12841),
            .I(N__12835));
    Span4Mux_v I__2100 (
            .O(N__12838),
            .I(N__12832));
    Span4Mux_h I__2099 (
            .O(N__12835),
            .I(N__12829));
    Span4Mux_h I__2098 (
            .O(N__12832),
            .I(N__12826));
    Odrv4 I__2097 (
            .O(N__12829),
            .I(\POWERLED.mult1_un89_sum ));
    Odrv4 I__2096 (
            .O(N__12826),
            .I(\POWERLED.mult1_un89_sum ));
    InMux I__2095 (
            .O(N__12821),
            .I(bfn_6_6_0_));
    InMux I__2094 (
            .O(N__12818),
            .I(N__12815));
    LocalMux I__2093 (
            .O(N__12815),
            .I(N__12812));
    Span4Mux_v I__2092 (
            .O(N__12812),
            .I(N__12808));
    InMux I__2091 (
            .O(N__12811),
            .I(N__12805));
    Span4Mux_h I__2090 (
            .O(N__12808),
            .I(N__12802));
    LocalMux I__2089 (
            .O(N__12805),
            .I(\POWERLED.mult1_un82_sum ));
    Odrv4 I__2088 (
            .O(N__12802),
            .I(\POWERLED.mult1_un82_sum ));
    InMux I__2087 (
            .O(N__12797),
            .I(\POWERLED.un1_dutycycle_1_cry_8 ));
    InMux I__2086 (
            .O(N__12794),
            .I(N__12790));
    InMux I__2085 (
            .O(N__12793),
            .I(N__12787));
    LocalMux I__2084 (
            .O(N__12790),
            .I(N__12784));
    LocalMux I__2083 (
            .O(N__12787),
            .I(\POWERLED.mult1_un75_sum ));
    Odrv12 I__2082 (
            .O(N__12784),
            .I(\POWERLED.mult1_un75_sum ));
    InMux I__2081 (
            .O(N__12779),
            .I(\POWERLED.un1_dutycycle_1_cry_9 ));
    InMux I__2080 (
            .O(N__12776),
            .I(\HDA_STRAP.un1_count_1_cry_11 ));
    InMux I__2079 (
            .O(N__12773),
            .I(\HDA_STRAP.un1_count_1_cry_12 ));
    InMux I__2078 (
            .O(N__12770),
            .I(\HDA_STRAP.un1_count_1_cry_13 ));
    InMux I__2077 (
            .O(N__12767),
            .I(\HDA_STRAP.un1_count_1_cry_14 ));
    InMux I__2076 (
            .O(N__12764),
            .I(bfn_6_3_0_));
    InMux I__2075 (
            .O(N__12761),
            .I(\HDA_STRAP.un1_count_1_cry_16 ));
    InMux I__2074 (
            .O(N__12758),
            .I(N__12754));
    InMux I__2073 (
            .O(N__12757),
            .I(N__12751));
    LocalMux I__2072 (
            .O(N__12754),
            .I(N__12746));
    LocalMux I__2071 (
            .O(N__12751),
            .I(N__12746));
    Span12Mux_s11_v I__2070 (
            .O(N__12746),
            .I(N__12743));
    Odrv12 I__2069 (
            .O(N__12743),
            .I(\POWERLED.un1_dutycycle_1_axb_0 ));
    CascadeMux I__2068 (
            .O(N__12740),
            .I(N__12737));
    InMux I__2067 (
            .O(N__12737),
            .I(N__12734));
    LocalMux I__2066 (
            .O(N__12734),
            .I(\POWERLED.un1_dutycycle_1_axb_1 ));
    InMux I__2065 (
            .O(N__12731),
            .I(N__12727));
    InMux I__2064 (
            .O(N__12730),
            .I(N__12724));
    LocalMux I__2063 (
            .O(N__12727),
            .I(N__12721));
    LocalMux I__2062 (
            .O(N__12724),
            .I(N__12718));
    Span4Mux_v I__2061 (
            .O(N__12721),
            .I(N__12715));
    Span12Mux_s11_v I__2060 (
            .O(N__12718),
            .I(N__12712));
    Odrv4 I__2059 (
            .O(N__12715),
            .I(\POWERLED.mult1_un138_sum ));
    Odrv12 I__2058 (
            .O(N__12712),
            .I(\POWERLED.mult1_un138_sum ));
    InMux I__2057 (
            .O(N__12707),
            .I(\POWERLED.un1_dutycycle_1_cry_0 ));
    InMux I__2056 (
            .O(N__12704),
            .I(N__12701));
    LocalMux I__2055 (
            .O(N__12701),
            .I(\POWERLED.dutycycle_RNI16B71Z0Z_5 ));
    CascadeMux I__2054 (
            .O(N__12698),
            .I(N__12694));
    InMux I__2053 (
            .O(N__12697),
            .I(N__12691));
    InMux I__2052 (
            .O(N__12694),
            .I(N__12688));
    LocalMux I__2051 (
            .O(N__12691),
            .I(\POWERLED.dutycycle_RNIFHLJZ0Z_0 ));
    LocalMux I__2050 (
            .O(N__12688),
            .I(\POWERLED.dutycycle_RNIFHLJZ0Z_0 ));
    InMux I__2049 (
            .O(N__12683),
            .I(N__12679));
    InMux I__2048 (
            .O(N__12682),
            .I(N__12676));
    LocalMux I__2047 (
            .O(N__12679),
            .I(N__12671));
    LocalMux I__2046 (
            .O(N__12676),
            .I(N__12671));
    Span4Mux_v I__2045 (
            .O(N__12671),
            .I(N__12668));
    Span4Mux_h I__2044 (
            .O(N__12668),
            .I(N__12665));
    Odrv4 I__2043 (
            .O(N__12665),
            .I(\POWERLED.mult1_un131_sum ));
    InMux I__2042 (
            .O(N__12662),
            .I(\POWERLED.un1_dutycycle_1_cry_1 ));
    InMux I__2041 (
            .O(N__12659),
            .I(\HDA_STRAP.un1_count_1_cry_2 ));
    InMux I__2040 (
            .O(N__12656),
            .I(\HDA_STRAP.un1_count_1_cry_3 ));
    InMux I__2039 (
            .O(N__12653),
            .I(\HDA_STRAP.un1_count_1_cry_4 ));
    InMux I__2038 (
            .O(N__12650),
            .I(\HDA_STRAP.un1_count_1_cry_5 ));
    InMux I__2037 (
            .O(N__12647),
            .I(\HDA_STRAP.un1_count_1_cry_6 ));
    InMux I__2036 (
            .O(N__12644),
            .I(bfn_6_2_0_));
    InMux I__2035 (
            .O(N__12641),
            .I(\HDA_STRAP.un1_count_1_cry_8 ));
    InMux I__2034 (
            .O(N__12638),
            .I(\HDA_STRAP.un1_count_1_cry_9 ));
    InMux I__2033 (
            .O(N__12635),
            .I(N__12632));
    LocalMux I__2032 (
            .O(N__12632),
            .I(\HDA_STRAP.count_RNO_0Z0Z_11 ));
    InMux I__2031 (
            .O(N__12629),
            .I(\HDA_STRAP.un1_count_1_cry_10 ));
    InMux I__2030 (
            .O(N__12626),
            .I(N__12623));
    LocalMux I__2029 (
            .O(N__12623),
            .I(N__12617));
    InMux I__2028 (
            .O(N__12622),
            .I(N__12614));
    InMux I__2027 (
            .O(N__12621),
            .I(N__12609));
    InMux I__2026 (
            .O(N__12620),
            .I(N__12609));
    Span4Mux_h I__2025 (
            .O(N__12617),
            .I(N__12606));
    LocalMux I__2024 (
            .O(N__12614),
            .I(\POWERLED.countZ0Z_13 ));
    LocalMux I__2023 (
            .O(N__12609),
            .I(\POWERLED.countZ0Z_13 ));
    Odrv4 I__2022 (
            .O(N__12606),
            .I(\POWERLED.countZ0Z_13 ));
    InMux I__2021 (
            .O(N__12599),
            .I(\POWERLED.un1_count_1_cry_12 ));
    InMux I__2020 (
            .O(N__12596),
            .I(N__12593));
    LocalMux I__2019 (
            .O(N__12593),
            .I(N__12587));
    InMux I__2018 (
            .O(N__12592),
            .I(N__12584));
    InMux I__2017 (
            .O(N__12591),
            .I(N__12581));
    InMux I__2016 (
            .O(N__12590),
            .I(N__12578));
    Span4Mux_h I__2015 (
            .O(N__12587),
            .I(N__12575));
    LocalMux I__2014 (
            .O(N__12584),
            .I(\POWERLED.countZ0Z_14 ));
    LocalMux I__2013 (
            .O(N__12581),
            .I(\POWERLED.countZ0Z_14 ));
    LocalMux I__2012 (
            .O(N__12578),
            .I(\POWERLED.countZ0Z_14 ));
    Odrv4 I__2011 (
            .O(N__12575),
            .I(\POWERLED.countZ0Z_14 ));
    InMux I__2010 (
            .O(N__12566),
            .I(\POWERLED.un1_count_1_cry_13 ));
    InMux I__2009 (
            .O(N__12563),
            .I(bfn_5_16_0_));
    InMux I__2008 (
            .O(N__12560),
            .I(N__12557));
    LocalMux I__2007 (
            .O(N__12557),
            .I(N__12553));
    InMux I__2006 (
            .O(N__12556),
            .I(N__12548));
    Span4Mux_h I__2005 (
            .O(N__12553),
            .I(N__12545));
    InMux I__2004 (
            .O(N__12552),
            .I(N__12540));
    InMux I__2003 (
            .O(N__12551),
            .I(N__12540));
    LocalMux I__2002 (
            .O(N__12548),
            .I(\POWERLED.countZ0Z_15 ));
    Odrv4 I__2001 (
            .O(N__12545),
            .I(\POWERLED.countZ0Z_15 ));
    LocalMux I__2000 (
            .O(N__12540),
            .I(\POWERLED.countZ0Z_15 ));
    CEMux I__1999 (
            .O(N__12533),
            .I(N__12530));
    LocalMux I__1998 (
            .O(N__12530),
            .I(N__12527));
    Odrv12 I__1997 (
            .O(N__12527),
            .I(\POWERLED.N_65_5 ));
    SRMux I__1996 (
            .O(N__12524),
            .I(N__12521));
    LocalMux I__1995 (
            .O(N__12521),
            .I(N__12516));
    SRMux I__1994 (
            .O(N__12520),
            .I(N__12511));
    SRMux I__1993 (
            .O(N__12519),
            .I(N__12508));
    Span4Mux_h I__1992 (
            .O(N__12516),
            .I(N__12505));
    SRMux I__1991 (
            .O(N__12515),
            .I(N__12502));
    InMux I__1990 (
            .O(N__12514),
            .I(N__12499));
    LocalMux I__1989 (
            .O(N__12511),
            .I(\POWERLED.curr_state_RNI75RB5Z0Z_0 ));
    LocalMux I__1988 (
            .O(N__12508),
            .I(\POWERLED.curr_state_RNI75RB5Z0Z_0 ));
    Odrv4 I__1987 (
            .O(N__12505),
            .I(\POWERLED.curr_state_RNI75RB5Z0Z_0 ));
    LocalMux I__1986 (
            .O(N__12502),
            .I(\POWERLED.curr_state_RNI75RB5Z0Z_0 ));
    LocalMux I__1985 (
            .O(N__12499),
            .I(\POWERLED.curr_state_RNI75RB5Z0Z_0 ));
    InMux I__1984 (
            .O(N__12488),
            .I(N__12485));
    LocalMux I__1983 (
            .O(N__12485),
            .I(\HDA_STRAP.count_RNO_0Z0Z_0 ));
    InMux I__1982 (
            .O(N__12482),
            .I(\HDA_STRAP.un1_count_1_cry_0 ));
    InMux I__1981 (
            .O(N__12479),
            .I(\HDA_STRAP.un1_count_1_cry_1 ));
    InMux I__1980 (
            .O(N__12476),
            .I(N__12473));
    LocalMux I__1979 (
            .O(N__12473),
            .I(N__12469));
    InMux I__1978 (
            .O(N__12472),
            .I(N__12464));
    Span4Mux_h I__1977 (
            .O(N__12469),
            .I(N__12461));
    InMux I__1976 (
            .O(N__12468),
            .I(N__12456));
    InMux I__1975 (
            .O(N__12467),
            .I(N__12456));
    LocalMux I__1974 (
            .O(N__12464),
            .I(\POWERLED.countZ0Z_4 ));
    Odrv4 I__1973 (
            .O(N__12461),
            .I(\POWERLED.countZ0Z_4 ));
    LocalMux I__1972 (
            .O(N__12456),
            .I(\POWERLED.countZ0Z_4 ));
    InMux I__1971 (
            .O(N__12449),
            .I(\POWERLED.un1_count_1_cry_3 ));
    InMux I__1970 (
            .O(N__12446),
            .I(N__12443));
    LocalMux I__1969 (
            .O(N__12443),
            .I(N__12437));
    InMux I__1968 (
            .O(N__12442),
            .I(N__12434));
    InMux I__1967 (
            .O(N__12441),
            .I(N__12429));
    InMux I__1966 (
            .O(N__12440),
            .I(N__12429));
    Span4Mux_v I__1965 (
            .O(N__12437),
            .I(N__12426));
    LocalMux I__1964 (
            .O(N__12434),
            .I(\POWERLED.countZ0Z_5 ));
    LocalMux I__1963 (
            .O(N__12429),
            .I(\POWERLED.countZ0Z_5 ));
    Odrv4 I__1962 (
            .O(N__12426),
            .I(\POWERLED.countZ0Z_5 ));
    InMux I__1961 (
            .O(N__12419),
            .I(\POWERLED.un1_count_1_cry_4 ));
    InMux I__1960 (
            .O(N__12416),
            .I(N__12413));
    LocalMux I__1959 (
            .O(N__12413),
            .I(N__12407));
    InMux I__1958 (
            .O(N__12412),
            .I(N__12404));
    InMux I__1957 (
            .O(N__12411),
            .I(N__12399));
    InMux I__1956 (
            .O(N__12410),
            .I(N__12399));
    Span4Mux_h I__1955 (
            .O(N__12407),
            .I(N__12396));
    LocalMux I__1954 (
            .O(N__12404),
            .I(\POWERLED.countZ0Z_6 ));
    LocalMux I__1953 (
            .O(N__12399),
            .I(\POWERLED.countZ0Z_6 ));
    Odrv4 I__1952 (
            .O(N__12396),
            .I(\POWERLED.countZ0Z_6 ));
    InMux I__1951 (
            .O(N__12389),
            .I(\POWERLED.un1_count_1_cry_5 ));
    CascadeMux I__1950 (
            .O(N__12386),
            .I(N__12381));
    InMux I__1949 (
            .O(N__12385),
            .I(N__12378));
    InMux I__1948 (
            .O(N__12384),
            .I(N__12372));
    InMux I__1947 (
            .O(N__12381),
            .I(N__12372));
    LocalMux I__1946 (
            .O(N__12378),
            .I(N__12369));
    InMux I__1945 (
            .O(N__12377),
            .I(N__12366));
    LocalMux I__1944 (
            .O(N__12372),
            .I(N__12361));
    Span4Mux_v I__1943 (
            .O(N__12369),
            .I(N__12361));
    LocalMux I__1942 (
            .O(N__12366),
            .I(\POWERLED.countZ0Z_7 ));
    Odrv4 I__1941 (
            .O(N__12361),
            .I(\POWERLED.countZ0Z_7 ));
    InMux I__1940 (
            .O(N__12356),
            .I(\POWERLED.un1_count_1_cry_6 ));
    InMux I__1939 (
            .O(N__12353),
            .I(N__12349));
    InMux I__1938 (
            .O(N__12352),
            .I(N__12344));
    LocalMux I__1937 (
            .O(N__12349),
            .I(N__12341));
    InMux I__1936 (
            .O(N__12348),
            .I(N__12336));
    InMux I__1935 (
            .O(N__12347),
            .I(N__12336));
    LocalMux I__1934 (
            .O(N__12344),
            .I(\POWERLED.countZ0Z_8 ));
    Odrv4 I__1933 (
            .O(N__12341),
            .I(\POWERLED.countZ0Z_8 ));
    LocalMux I__1932 (
            .O(N__12336),
            .I(\POWERLED.countZ0Z_8 ));
    InMux I__1931 (
            .O(N__12329),
            .I(\POWERLED.un1_count_1_cry_7 ));
    InMux I__1930 (
            .O(N__12326),
            .I(N__12322));
    CascadeMux I__1929 (
            .O(N__12325),
            .I(N__12317));
    LocalMux I__1928 (
            .O(N__12322),
            .I(N__12314));
    InMux I__1927 (
            .O(N__12321),
            .I(N__12311));
    InMux I__1926 (
            .O(N__12320),
            .I(N__12308));
    InMux I__1925 (
            .O(N__12317),
            .I(N__12305));
    Span4Mux_v I__1924 (
            .O(N__12314),
            .I(N__12302));
    LocalMux I__1923 (
            .O(N__12311),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__1922 (
            .O(N__12308),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__1921 (
            .O(N__12305),
            .I(\POWERLED.countZ0Z_9 ));
    Odrv4 I__1920 (
            .O(N__12302),
            .I(\POWERLED.countZ0Z_9 ));
    InMux I__1919 (
            .O(N__12293),
            .I(bfn_5_15_0_));
    InMux I__1918 (
            .O(N__12290),
            .I(N__12287));
    LocalMux I__1917 (
            .O(N__12287),
            .I(N__12283));
    InMux I__1916 (
            .O(N__12286),
            .I(N__12278));
    Span4Mux_v I__1915 (
            .O(N__12283),
            .I(N__12275));
    InMux I__1914 (
            .O(N__12282),
            .I(N__12270));
    InMux I__1913 (
            .O(N__12281),
            .I(N__12270));
    LocalMux I__1912 (
            .O(N__12278),
            .I(\POWERLED.countZ0Z_10 ));
    Odrv4 I__1911 (
            .O(N__12275),
            .I(\POWERLED.countZ0Z_10 ));
    LocalMux I__1910 (
            .O(N__12270),
            .I(\POWERLED.countZ0Z_10 ));
    InMux I__1909 (
            .O(N__12263),
            .I(\POWERLED.un1_count_1_cry_9 ));
    InMux I__1908 (
            .O(N__12260),
            .I(N__12257));
    LocalMux I__1907 (
            .O(N__12257),
            .I(N__12251));
    InMux I__1906 (
            .O(N__12256),
            .I(N__12248));
    InMux I__1905 (
            .O(N__12255),
            .I(N__12245));
    InMux I__1904 (
            .O(N__12254),
            .I(N__12242));
    Span4Mux_h I__1903 (
            .O(N__12251),
            .I(N__12239));
    LocalMux I__1902 (
            .O(N__12248),
            .I(\POWERLED.countZ0Z_11 ));
    LocalMux I__1901 (
            .O(N__12245),
            .I(\POWERLED.countZ0Z_11 ));
    LocalMux I__1900 (
            .O(N__12242),
            .I(\POWERLED.countZ0Z_11 ));
    Odrv4 I__1899 (
            .O(N__12239),
            .I(\POWERLED.countZ0Z_11 ));
    InMux I__1898 (
            .O(N__12230),
            .I(\POWERLED.un1_count_1_cry_10 ));
    InMux I__1897 (
            .O(N__12227),
            .I(N__12224));
    LocalMux I__1896 (
            .O(N__12224),
            .I(N__12218));
    InMux I__1895 (
            .O(N__12223),
            .I(N__12215));
    InMux I__1894 (
            .O(N__12222),
            .I(N__12212));
    InMux I__1893 (
            .O(N__12221),
            .I(N__12209));
    Span4Mux_h I__1892 (
            .O(N__12218),
            .I(N__12206));
    LocalMux I__1891 (
            .O(N__12215),
            .I(\POWERLED.countZ0Z_12 ));
    LocalMux I__1890 (
            .O(N__12212),
            .I(\POWERLED.countZ0Z_12 ));
    LocalMux I__1889 (
            .O(N__12209),
            .I(\POWERLED.countZ0Z_12 ));
    Odrv4 I__1888 (
            .O(N__12206),
            .I(\POWERLED.countZ0Z_12 ));
    InMux I__1887 (
            .O(N__12197),
            .I(\POWERLED.un1_count_1_cry_11 ));
    InMux I__1886 (
            .O(N__12194),
            .I(N__12190));
    InMux I__1885 (
            .O(N__12193),
            .I(N__12187));
    LocalMux I__1884 (
            .O(N__12190),
            .I(N__12184));
    LocalMux I__1883 (
            .O(N__12187),
            .I(\POWERLED.count_offZ0Z_8 ));
    Odrv4 I__1882 (
            .O(N__12184),
            .I(\POWERLED.count_offZ0Z_8 ));
    InMux I__1881 (
            .O(N__12179),
            .I(N__12175));
    InMux I__1880 (
            .O(N__12178),
            .I(N__12172));
    LocalMux I__1879 (
            .O(N__12175),
            .I(N__12169));
    LocalMux I__1878 (
            .O(N__12172),
            .I(\POWERLED.count_offZ0Z_6 ));
    Odrv4 I__1877 (
            .O(N__12169),
            .I(\POWERLED.count_offZ0Z_6 ));
    CascadeMux I__1876 (
            .O(N__12164),
            .I(N__12160));
    InMux I__1875 (
            .O(N__12163),
            .I(N__12157));
    InMux I__1874 (
            .O(N__12160),
            .I(N__12154));
    LocalMux I__1873 (
            .O(N__12157),
            .I(\POWERLED.count_offZ0Z_9 ));
    LocalMux I__1872 (
            .O(N__12154),
            .I(\POWERLED.count_offZ0Z_9 ));
    InMux I__1871 (
            .O(N__12149),
            .I(N__12145));
    InMux I__1870 (
            .O(N__12148),
            .I(N__12142));
    LocalMux I__1869 (
            .O(N__12145),
            .I(N__12139));
    LocalMux I__1868 (
            .O(N__12142),
            .I(\POWERLED.count_offZ0Z_5 ));
    Odrv4 I__1867 (
            .O(N__12139),
            .I(\POWERLED.count_offZ0Z_5 ));
    InMux I__1866 (
            .O(N__12134),
            .I(N__12131));
    LocalMux I__1865 (
            .O(N__12131),
            .I(\POWERLED.func_state_ns_0_a2_11_0 ));
    InMux I__1864 (
            .O(N__12128),
            .I(N__12125));
    LocalMux I__1863 (
            .O(N__12125),
            .I(\POWERLED.func_state_ns_0_a2_10_0 ));
    CascadeMux I__1862 (
            .O(N__12122),
            .I(\POWERLED.func_state_ns_0_a2_9_0_cascade_ ));
    InMux I__1861 (
            .O(N__12119),
            .I(N__12105));
    InMux I__1860 (
            .O(N__12118),
            .I(N__12098));
    InMux I__1859 (
            .O(N__12117),
            .I(N__12098));
    InMux I__1858 (
            .O(N__12116),
            .I(N__12098));
    InMux I__1857 (
            .O(N__12115),
            .I(N__12089));
    InMux I__1856 (
            .O(N__12114),
            .I(N__12089));
    InMux I__1855 (
            .O(N__12113),
            .I(N__12089));
    InMux I__1854 (
            .O(N__12112),
            .I(N__12089));
    InMux I__1853 (
            .O(N__12111),
            .I(N__12080));
    InMux I__1852 (
            .O(N__12110),
            .I(N__12080));
    InMux I__1851 (
            .O(N__12109),
            .I(N__12080));
    InMux I__1850 (
            .O(N__12108),
            .I(N__12080));
    LocalMux I__1849 (
            .O(N__12105),
            .I(N__12075));
    LocalMux I__1848 (
            .O(N__12098),
            .I(N__12075));
    LocalMux I__1847 (
            .O(N__12089),
            .I(\POWERLED.count_off_0_sqmuxa ));
    LocalMux I__1846 (
            .O(N__12080),
            .I(\POWERLED.count_off_0_sqmuxa ));
    Odrv12 I__1845 (
            .O(N__12075),
            .I(\POWERLED.count_off_0_sqmuxa ));
    CascadeMux I__1844 (
            .O(N__12068),
            .I(\POWERLED.count_off_0_sqmuxa_cascade_ ));
    InMux I__1843 (
            .O(N__12065),
            .I(N__12059));
    InMux I__1842 (
            .O(N__12064),
            .I(N__12052));
    InMux I__1841 (
            .O(N__12063),
            .I(N__12052));
    InMux I__1840 (
            .O(N__12062),
            .I(N__12052));
    LocalMux I__1839 (
            .O(N__12059),
            .I(N__12049));
    LocalMux I__1838 (
            .O(N__12052),
            .I(N__12046));
    Odrv4 I__1837 (
            .O(N__12049),
            .I(\POWERLED.N_85_1 ));
    Odrv12 I__1836 (
            .O(N__12046),
            .I(\POWERLED.N_85_1 ));
    InMux I__1835 (
            .O(N__12041),
            .I(N__12035));
    InMux I__1834 (
            .O(N__12040),
            .I(N__12030));
    InMux I__1833 (
            .O(N__12039),
            .I(N__12030));
    InMux I__1832 (
            .O(N__12038),
            .I(N__12027));
    LocalMux I__1831 (
            .O(N__12035),
            .I(N__12024));
    LocalMux I__1830 (
            .O(N__12030),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__1829 (
            .O(N__12027),
            .I(\POWERLED.countZ0Z_0 ));
    Odrv4 I__1828 (
            .O(N__12024),
            .I(\POWERLED.countZ0Z_0 ));
    InMux I__1827 (
            .O(N__12017),
            .I(N__12012));
    CascadeMux I__1826 (
            .O(N__12016),
            .I(N__12009));
    InMux I__1825 (
            .O(N__12015),
            .I(N__12006));
    LocalMux I__1824 (
            .O(N__12012),
            .I(N__12003));
    InMux I__1823 (
            .O(N__12009),
            .I(N__12000));
    LocalMux I__1822 (
            .O(N__12006),
            .I(N__11995));
    Span4Mux_s2_h I__1821 (
            .O(N__12003),
            .I(N__11995));
    LocalMux I__1820 (
            .O(N__12000),
            .I(\POWERLED.countZ0Z_1 ));
    Odrv4 I__1819 (
            .O(N__11995),
            .I(\POWERLED.countZ0Z_1 ));
    InMux I__1818 (
            .O(N__11990),
            .I(N__11987));
    LocalMux I__1817 (
            .O(N__11987),
            .I(N__11983));
    InMux I__1816 (
            .O(N__11986),
            .I(N__11978));
    Span4Mux_v I__1815 (
            .O(N__11983),
            .I(N__11975));
    InMux I__1814 (
            .O(N__11982),
            .I(N__11970));
    InMux I__1813 (
            .O(N__11981),
            .I(N__11970));
    LocalMux I__1812 (
            .O(N__11978),
            .I(\POWERLED.countZ0Z_2 ));
    Odrv4 I__1811 (
            .O(N__11975),
            .I(\POWERLED.countZ0Z_2 ));
    LocalMux I__1810 (
            .O(N__11970),
            .I(\POWERLED.countZ0Z_2 ));
    InMux I__1809 (
            .O(N__11963),
            .I(\POWERLED.un1_count_1_cry_1 ));
    InMux I__1808 (
            .O(N__11960),
            .I(N__11957));
    LocalMux I__1807 (
            .O(N__11957),
            .I(N__11953));
    InMux I__1806 (
            .O(N__11956),
            .I(N__11948));
    Span4Mux_h I__1805 (
            .O(N__11953),
            .I(N__11945));
    InMux I__1804 (
            .O(N__11952),
            .I(N__11940));
    InMux I__1803 (
            .O(N__11951),
            .I(N__11940));
    LocalMux I__1802 (
            .O(N__11948),
            .I(\POWERLED.countZ0Z_3 ));
    Odrv4 I__1801 (
            .O(N__11945),
            .I(\POWERLED.countZ0Z_3 ));
    LocalMux I__1800 (
            .O(N__11940),
            .I(\POWERLED.countZ0Z_3 ));
    InMux I__1799 (
            .O(N__11933),
            .I(\POWERLED.un1_count_1_cry_2 ));
    InMux I__1798 (
            .O(N__11930),
            .I(\POWERLED.un1_count_off_1_cry_8 ));
    InMux I__1797 (
            .O(N__11927),
            .I(\POWERLED.un1_count_off_1_cry_9 ));
    InMux I__1796 (
            .O(N__11924),
            .I(\POWERLED.un1_count_off_1_cry_10 ));
    InMux I__1795 (
            .O(N__11921),
            .I(\POWERLED.un1_count_off_1_cry_11 ));
    InMux I__1794 (
            .O(N__11918),
            .I(\POWERLED.un1_count_off_1_cry_12 ));
    InMux I__1793 (
            .O(N__11915),
            .I(\POWERLED.un1_count_off_1_cry_13 ));
    InMux I__1792 (
            .O(N__11912),
            .I(\POWERLED.un1_count_off_1_cry_14 ));
    InMux I__1791 (
            .O(N__11909),
            .I(N__11905));
    InMux I__1790 (
            .O(N__11908),
            .I(N__11902));
    LocalMux I__1789 (
            .O(N__11905),
            .I(\POWERLED.count_offZ0Z_12 ));
    LocalMux I__1788 (
            .O(N__11902),
            .I(\POWERLED.count_offZ0Z_12 ));
    InMux I__1787 (
            .O(N__11897),
            .I(N__11893));
    InMux I__1786 (
            .O(N__11896),
            .I(N__11890));
    LocalMux I__1785 (
            .O(N__11893),
            .I(\POWERLED.count_offZ0Z_13 ));
    LocalMux I__1784 (
            .O(N__11890),
            .I(\POWERLED.count_offZ0Z_13 ));
    CascadeMux I__1783 (
            .O(N__11885),
            .I(N__11881));
    InMux I__1782 (
            .O(N__11884),
            .I(N__11878));
    InMux I__1781 (
            .O(N__11881),
            .I(N__11875));
    LocalMux I__1780 (
            .O(N__11878),
            .I(\POWERLED.count_offZ0Z_15 ));
    LocalMux I__1779 (
            .O(N__11875),
            .I(\POWERLED.count_offZ0Z_15 ));
    InMux I__1778 (
            .O(N__11870),
            .I(N__11866));
    InMux I__1777 (
            .O(N__11869),
            .I(N__11863));
    LocalMux I__1776 (
            .O(N__11866),
            .I(N__11860));
    LocalMux I__1775 (
            .O(N__11863),
            .I(\POWERLED.count_offZ0Z_1 ));
    Odrv4 I__1774 (
            .O(N__11860),
            .I(\POWERLED.count_offZ0Z_1 ));
    InMux I__1773 (
            .O(N__11855),
            .I(N__11851));
    InMux I__1772 (
            .O(N__11854),
            .I(N__11848));
    LocalMux I__1771 (
            .O(N__11851),
            .I(\POWERLED.count_offZ0Z_11 ));
    LocalMux I__1770 (
            .O(N__11848),
            .I(\POWERLED.count_offZ0Z_11 ));
    InMux I__1769 (
            .O(N__11843),
            .I(N__11839));
    InMux I__1768 (
            .O(N__11842),
            .I(N__11836));
    LocalMux I__1767 (
            .O(N__11839),
            .I(N__11833));
    LocalMux I__1766 (
            .O(N__11836),
            .I(\POWERLED.count_offZ0Z_0 ));
    Odrv4 I__1765 (
            .O(N__11833),
            .I(\POWERLED.count_offZ0Z_0 ));
    CascadeMux I__1764 (
            .O(N__11828),
            .I(N__11824));
    InMux I__1763 (
            .O(N__11827),
            .I(N__11821));
    InMux I__1762 (
            .O(N__11824),
            .I(N__11818));
    LocalMux I__1761 (
            .O(N__11821),
            .I(\POWERLED.count_offZ0Z_14 ));
    LocalMux I__1760 (
            .O(N__11818),
            .I(\POWERLED.count_offZ0Z_14 ));
    InMux I__1759 (
            .O(N__11813),
            .I(N__11809));
    InMux I__1758 (
            .O(N__11812),
            .I(N__11806));
    LocalMux I__1757 (
            .O(N__11809),
            .I(\POWERLED.count_offZ0Z_10 ));
    LocalMux I__1756 (
            .O(N__11806),
            .I(\POWERLED.count_offZ0Z_10 ));
    InMux I__1755 (
            .O(N__11801),
            .I(\POWERLED.un1_count_off_1_cry_0 ));
    InMux I__1754 (
            .O(N__11798),
            .I(\POWERLED.un1_count_off_1_cry_1 ));
    InMux I__1753 (
            .O(N__11795),
            .I(\POWERLED.un1_count_off_1_cry_2 ));
    InMux I__1752 (
            .O(N__11792),
            .I(\POWERLED.un1_count_off_1_cry_3 ));
    InMux I__1751 (
            .O(N__11789),
            .I(\POWERLED.un1_count_off_1_cry_4 ));
    InMux I__1750 (
            .O(N__11786),
            .I(\POWERLED.un1_count_off_1_cry_5 ));
    InMux I__1749 (
            .O(N__11783),
            .I(\POWERLED.un1_count_off_1_cry_6 ));
    InMux I__1748 (
            .O(N__11780),
            .I(bfn_5_10_0_));
    CascadeMux I__1747 (
            .O(N__11777),
            .I(N__11774));
    InMux I__1746 (
            .O(N__11774),
            .I(N__11771));
    LocalMux I__1745 (
            .O(N__11771),
            .I(\POWERLED.un1_dutycycle_1_i_29 ));
    InMux I__1744 (
            .O(N__11768),
            .I(N__11765));
    LocalMux I__1743 (
            .O(N__11765),
            .I(N__11762));
    Odrv4 I__1742 (
            .O(N__11762),
            .I(\POWERLED.mult1_un61_sum_i ));
    InMux I__1741 (
            .O(N__11759),
            .I(N__11756));
    LocalMux I__1740 (
            .O(N__11756),
            .I(\POWERLED.mult1_un54_sum_i ));
    InMux I__1739 (
            .O(N__11753),
            .I(N__11750));
    LocalMux I__1738 (
            .O(N__11750),
            .I(N__11747));
    Odrv12 I__1737 (
            .O(N__11747),
            .I(\POWERLED.mult1_un75_sum_i ));
    InMux I__1736 (
            .O(N__11744),
            .I(N__11738));
    InMux I__1735 (
            .O(N__11743),
            .I(N__11738));
    LocalMux I__1734 (
            .O(N__11738),
            .I(N__11735));
    Span4Mux_h I__1733 (
            .O(N__11735),
            .I(N__11732));
    Odrv4 I__1732 (
            .O(N__11732),
            .I(\POWERLED.N_53 ));
    CascadeMux I__1731 (
            .O(N__11729),
            .I(N__11726));
    InMux I__1730 (
            .O(N__11726),
            .I(N__11723));
    LocalMux I__1729 (
            .O(N__11723),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_4 ));
    CascadeMux I__1728 (
            .O(N__11720),
            .I(N__11717));
    InMux I__1727 (
            .O(N__11717),
            .I(N__11714));
    LocalMux I__1726 (
            .O(N__11714),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_5 ));
    CascadeMux I__1725 (
            .O(N__11711),
            .I(N__11708));
    InMux I__1724 (
            .O(N__11708),
            .I(N__11705));
    LocalMux I__1723 (
            .O(N__11705),
            .I(\POWERLED.mult1_un47_sum_axb_4 ));
    InMux I__1722 (
            .O(N__11702),
            .I(N__11698));
    InMux I__1721 (
            .O(N__11701),
            .I(N__11695));
    LocalMux I__1720 (
            .O(N__11698),
            .I(\HDA_STRAP.N_5_0 ));
    LocalMux I__1719 (
            .O(N__11695),
            .I(\HDA_STRAP.N_5_0 ));
    InMux I__1718 (
            .O(N__11690),
            .I(N__11684));
    InMux I__1717 (
            .O(N__11689),
            .I(N__11684));
    LocalMux I__1716 (
            .O(N__11684),
            .I(\HDA_STRAP.curr_stateZ0Z_2 ));
    IoInMux I__1715 (
            .O(N__11681),
            .I(N__11678));
    LocalMux I__1714 (
            .O(N__11678),
            .I(N__11675));
    IoSpan4Mux I__1713 (
            .O(N__11675),
            .I(N__11672));
    Span4Mux_s0_h I__1712 (
            .O(N__11672),
            .I(N__11669));
    Span4Mux_h I__1711 (
            .O(N__11669),
            .I(N__11666));
    Odrv4 I__1710 (
            .O(N__11666),
            .I(hda_sdo_atp));
    InMux I__1709 (
            .O(N__11663),
            .I(N__11660));
    LocalMux I__1708 (
            .O(N__11660),
            .I(N__11657));
    Odrv12 I__1707 (
            .O(N__11657),
            .I(\POWERLED.mult1_un82_sum_i ));
    CascadeMux I__1706 (
            .O(N__11654),
            .I(N__11651));
    InMux I__1705 (
            .O(N__11651),
            .I(N__11648));
    LocalMux I__1704 (
            .O(N__11648),
            .I(\POWERLED.un1_dutycycle_1_i_28 ));
    CascadeMux I__1703 (
            .O(N__11645),
            .I(\POWERLED.un1_dutycycle_1_19_0_cascade_ ));
    CascadeMux I__1702 (
            .O(N__11642),
            .I(\POWERLED.un1_countlto15_5_cascade_ ));
    InMux I__1701 (
            .O(N__11639),
            .I(N__11636));
    LocalMux I__1700 (
            .O(N__11636),
            .I(\POWERLED.g0_0_4 ));
    InMux I__1699 (
            .O(N__11633),
            .I(N__11630));
    LocalMux I__1698 (
            .O(N__11630),
            .I(\POWERLED.un1_countlt6 ));
    InMux I__1697 (
            .O(N__11627),
            .I(N__11624));
    LocalMux I__1696 (
            .O(N__11624),
            .I(\POWERLED.g0_0_5 ));
    CascadeMux I__1695 (
            .O(N__11621),
            .I(\POWERLED.un1_countlto15_4_cascade_ ));
    InMux I__1694 (
            .O(N__11618),
            .I(N__11615));
    LocalMux I__1693 (
            .O(N__11615),
            .I(\POWERLED.un1_countlto15_7 ));
    InMux I__1692 (
            .O(N__11612),
            .I(N__11609));
    LocalMux I__1691 (
            .O(N__11609),
            .I(N__11606));
    Odrv4 I__1690 (
            .O(N__11606),
            .I(\POWERLED.count_RNIOVT24Z0Z_11 ));
    InMux I__1689 (
            .O(N__11603),
            .I(N__11597));
    InMux I__1688 (
            .O(N__11602),
            .I(N__11594));
    InMux I__1687 (
            .O(N__11601),
            .I(N__11591));
    InMux I__1686 (
            .O(N__11600),
            .I(N__11588));
    LocalMux I__1685 (
            .O(N__11597),
            .I(N__11585));
    LocalMux I__1684 (
            .O(N__11594),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    LocalMux I__1683 (
            .O(N__11591),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    LocalMux I__1682 (
            .O(N__11588),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    Odrv12 I__1681 (
            .O(N__11585),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    CascadeMux I__1680 (
            .O(N__11576),
            .I(\POWERLED.count_RNIOVT24Z0Z_11_cascade_ ));
    IoInMux I__1679 (
            .O(N__11573),
            .I(N__11570));
    LocalMux I__1678 (
            .O(N__11570),
            .I(N__11566));
    IoInMux I__1677 (
            .O(N__11569),
            .I(N__11563));
    Span4Mux_s3_h I__1676 (
            .O(N__11566),
            .I(N__11560));
    LocalMux I__1675 (
            .O(N__11563),
            .I(N__11557));
    Odrv4 I__1674 (
            .O(N__11560),
            .I(v5s_enn));
    Odrv12 I__1673 (
            .O(N__11557),
            .I(v5s_enn));
    InMux I__1672 (
            .O(N__11552),
            .I(N__11549));
    LocalMux I__1671 (
            .O(N__11549),
            .I(N__11546));
    Span4Mux_v I__1670 (
            .O(N__11546),
            .I(N__11543));
    Odrv4 I__1669 (
            .O(N__11543),
            .I(\POWERLED.mult1_un159_sum_i ));
    InMux I__1668 (
            .O(N__11540),
            .I(N__11537));
    LocalMux I__1667 (
            .O(N__11537),
            .I(N__11534));
    Odrv4 I__1666 (
            .O(N__11534),
            .I(\POWERLED.mult1_un152_sum_i ));
    CascadeMux I__1665 (
            .O(N__11531),
            .I(\POWERLED.un1_countlt6_0_cascade_ ));
    CascadeMux I__1664 (
            .O(N__11528),
            .I(\POWERLED.g0_0_7_cascade_ ));
    InMux I__1663 (
            .O(N__11525),
            .I(N__11522));
    LocalMux I__1662 (
            .O(N__11522),
            .I(N__11519));
    Span4Mux_s3_h I__1661 (
            .O(N__11519),
            .I(N__11516));
    Odrv4 I__1660 (
            .O(N__11516),
            .I(\POWERLED.un1_count_0 ));
    InMux I__1659 (
            .O(N__11513),
            .I(N__11509));
    InMux I__1658 (
            .O(N__11512),
            .I(N__11506));
    LocalMux I__1657 (
            .O(N__11509),
            .I(\POWERLED.mult1_un47_sum_cry_6_s ));
    LocalMux I__1656 (
            .O(N__11506),
            .I(\POWERLED.mult1_un47_sum_cry_6_s ));
    CascadeMux I__1655 (
            .O(N__11501),
            .I(N__11496));
    InMux I__1654 (
            .O(N__11500),
            .I(N__11488));
    InMux I__1653 (
            .O(N__11499),
            .I(N__11488));
    InMux I__1652 (
            .O(N__11496),
            .I(N__11488));
    InMux I__1651 (
            .O(N__11495),
            .I(N__11485));
    LocalMux I__1650 (
            .O(N__11488),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    LocalMux I__1649 (
            .O(N__11485),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    CascadeMux I__1648 (
            .O(N__11480),
            .I(N__11477));
    InMux I__1647 (
            .O(N__11477),
            .I(N__11474));
    LocalMux I__1646 (
            .O(N__11474),
            .I(N__11471));
    Odrv4 I__1645 (
            .O(N__11471),
            .I(\POWERLED.mult1_un54_sum_cry_6_THRU_CO ));
    InMux I__1644 (
            .O(N__11468),
            .I(\POWERLED.mult1_un61_sum_cry_7 ));
    InMux I__1643 (
            .O(N__11465),
            .I(N__11461));
    CascadeMux I__1642 (
            .O(N__11464),
            .I(N__11457));
    LocalMux I__1641 (
            .O(N__11461),
            .I(N__11454));
    InMux I__1640 (
            .O(N__11460),
            .I(N__11449));
    InMux I__1639 (
            .O(N__11457),
            .I(N__11449));
    Span4Mux_v I__1638 (
            .O(N__11454),
            .I(N__11442));
    LocalMux I__1637 (
            .O(N__11449),
            .I(N__11442));
    InMux I__1636 (
            .O(N__11448),
            .I(N__11439));
    InMux I__1635 (
            .O(N__11447),
            .I(N__11436));
    Odrv4 I__1634 (
            .O(N__11442),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__1633 (
            .O(N__11439),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__1632 (
            .O(N__11436),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    CascadeMux I__1631 (
            .O(N__11429),
            .I(N__11425));
    CascadeMux I__1630 (
            .O(N__11428),
            .I(N__11421));
    InMux I__1629 (
            .O(N__11425),
            .I(N__11414));
    InMux I__1628 (
            .O(N__11424),
            .I(N__11414));
    InMux I__1627 (
            .O(N__11421),
            .I(N__11414));
    LocalMux I__1626 (
            .O(N__11414),
            .I(N__11411));
    Odrv4 I__1625 (
            .O(N__11411),
            .I(\POWERLED.mult1_un61_sum_i_0_8 ));
    InMux I__1624 (
            .O(N__11408),
            .I(N__11405));
    LocalMux I__1623 (
            .O(N__11405),
            .I(N__11402));
    Span4Mux_h I__1622 (
            .O(N__11402),
            .I(N__11399));
    Odrv4 I__1621 (
            .O(N__11399),
            .I(\POWERLED.mult1_un110_sum_i ));
    InMux I__1620 (
            .O(N__11396),
            .I(N__11393));
    LocalMux I__1619 (
            .O(N__11393),
            .I(N__11390));
    Span4Mux_s3_h I__1618 (
            .O(N__11390),
            .I(N__11387));
    Sp12to4 I__1617 (
            .O(N__11387),
            .I(N__11384));
    Odrv12 I__1616 (
            .O(N__11384),
            .I(\POWERLED.mult1_un138_sum_i ));
    InMux I__1615 (
            .O(N__11381),
            .I(N__11378));
    LocalMux I__1614 (
            .O(N__11378),
            .I(N__11375));
    Span4Mux_h I__1613 (
            .O(N__11375),
            .I(N__11372));
    Odrv4 I__1612 (
            .O(N__11372),
            .I(\POWERLED.mult1_un124_sum_i ));
    InMux I__1611 (
            .O(N__11369),
            .I(N__11366));
    LocalMux I__1610 (
            .O(N__11366),
            .I(N__11363));
    Odrv4 I__1609 (
            .O(N__11363),
            .I(\POWERLED.mult1_un117_sum_i ));
    InMux I__1608 (
            .O(N__11360),
            .I(N__11357));
    LocalMux I__1607 (
            .O(N__11357),
            .I(N__11353));
    InMux I__1606 (
            .O(N__11356),
            .I(N__11350));
    Odrv4 I__1605 (
            .O(N__11353),
            .I(\POWERLED.mult1_un138_sum_cry_6_s ));
    LocalMux I__1604 (
            .O(N__11350),
            .I(\POWERLED.mult1_un138_sum_cry_6_s ));
    CascadeMux I__1603 (
            .O(N__11345),
            .I(N__11342));
    InMux I__1602 (
            .O(N__11342),
            .I(N__11339));
    LocalMux I__1601 (
            .O(N__11339),
            .I(N__11336));
    Odrv4 I__1600 (
            .O(N__11336),
            .I(\POWERLED.mult1_un145_sum_axb_7_l_fx ));
    CascadeMux I__1599 (
            .O(N__11333),
            .I(N__11327));
    InMux I__1598 (
            .O(N__11332),
            .I(N__11320));
    InMux I__1597 (
            .O(N__11331),
            .I(N__11320));
    InMux I__1596 (
            .O(N__11330),
            .I(N__11315));
    InMux I__1595 (
            .O(N__11327),
            .I(N__11315));
    InMux I__1594 (
            .O(N__11326),
            .I(N__11312));
    InMux I__1593 (
            .O(N__11325),
            .I(N__11309));
    LocalMux I__1592 (
            .O(N__11320),
            .I(N__11306));
    LocalMux I__1591 (
            .O(N__11315),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__1590 (
            .O(N__11312),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__1589 (
            .O(N__11309),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    Odrv12 I__1588 (
            .O(N__11306),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    InMux I__1587 (
            .O(N__11297),
            .I(N__11294));
    LocalMux I__1586 (
            .O(N__11294),
            .I(N__11291));
    Span4Mux_s3_h I__1585 (
            .O(N__11291),
            .I(N__11288));
    Odrv4 I__1584 (
            .O(N__11288),
            .I(\POWERLED.un1_count_2_4 ));
    InMux I__1583 (
            .O(N__11285),
            .I(N__11282));
    LocalMux I__1582 (
            .O(N__11282),
            .I(N__11279));
    Odrv12 I__1581 (
            .O(N__11279),
            .I(\POWERLED.mult1_un68_sum_i ));
    CascadeMux I__1580 (
            .O(N__11276),
            .I(N__11273));
    InMux I__1579 (
            .O(N__11273),
            .I(N__11270));
    LocalMux I__1578 (
            .O(N__11270),
            .I(N__11267));
    Odrv4 I__1577 (
            .O(N__11267),
            .I(\POWERLED.mult1_un61_sum_cry_3_s ));
    InMux I__1576 (
            .O(N__11264),
            .I(\POWERLED.mult1_un61_sum_cry_2 ));
    CascadeMux I__1575 (
            .O(N__11261),
            .I(N__11258));
    InMux I__1574 (
            .O(N__11258),
            .I(N__11255));
    LocalMux I__1573 (
            .O(N__11255),
            .I(N__11252));
    Span4Mux_h I__1572 (
            .O(N__11252),
            .I(N__11249));
    Odrv4 I__1571 (
            .O(N__11249),
            .I(\POWERLED.mult1_un54_sum_cry_3_s ));
    InMux I__1570 (
            .O(N__11246),
            .I(N__11243));
    LocalMux I__1569 (
            .O(N__11243),
            .I(N__11240));
    Odrv4 I__1568 (
            .O(N__11240),
            .I(\POWERLED.mult1_un61_sum_cry_4_s ));
    InMux I__1567 (
            .O(N__11237),
            .I(\POWERLED.mult1_un61_sum_cry_3 ));
    InMux I__1566 (
            .O(N__11234),
            .I(N__11231));
    LocalMux I__1565 (
            .O(N__11231),
            .I(N__11228));
    Odrv12 I__1564 (
            .O(N__11228),
            .I(\POWERLED.mult1_un54_sum_cry_4_s ));
    CascadeMux I__1563 (
            .O(N__11225),
            .I(N__11222));
    InMux I__1562 (
            .O(N__11222),
            .I(N__11219));
    LocalMux I__1561 (
            .O(N__11219),
            .I(N__11216));
    Odrv4 I__1560 (
            .O(N__11216),
            .I(\POWERLED.mult1_un61_sum_cry_5_s ));
    InMux I__1559 (
            .O(N__11213),
            .I(\POWERLED.mult1_un61_sum_cry_4 ));
    CascadeMux I__1558 (
            .O(N__11210),
            .I(N__11207));
    InMux I__1557 (
            .O(N__11207),
            .I(N__11204));
    LocalMux I__1556 (
            .O(N__11204),
            .I(N__11201));
    Odrv4 I__1555 (
            .O(N__11201),
            .I(\POWERLED.mult1_un54_sum_cry_5_s ));
    InMux I__1554 (
            .O(N__11198),
            .I(N__11195));
    LocalMux I__1553 (
            .O(N__11195),
            .I(N__11192));
    Odrv4 I__1552 (
            .O(N__11192),
            .I(\POWERLED.mult1_un61_sum_cry_6_s ));
    InMux I__1551 (
            .O(N__11189),
            .I(\POWERLED.mult1_un61_sum_cry_5 ));
    InMux I__1550 (
            .O(N__11186),
            .I(N__11183));
    LocalMux I__1549 (
            .O(N__11183),
            .I(N__11180));
    Odrv4 I__1548 (
            .O(N__11180),
            .I(\POWERLED.mult1_un54_sum_cry_6_s ));
    CascadeMux I__1547 (
            .O(N__11177),
            .I(N__11173));
    CascadeMux I__1546 (
            .O(N__11176),
            .I(N__11169));
    InMux I__1545 (
            .O(N__11173),
            .I(N__11162));
    InMux I__1544 (
            .O(N__11172),
            .I(N__11162));
    InMux I__1543 (
            .O(N__11169),
            .I(N__11162));
    LocalMux I__1542 (
            .O(N__11162),
            .I(\POWERLED.mult1_un54_sum_i_8 ));
    InMux I__1541 (
            .O(N__11159),
            .I(N__11156));
    LocalMux I__1540 (
            .O(N__11156),
            .I(N__11153));
    Odrv4 I__1539 (
            .O(N__11153),
            .I(\POWERLED.mult1_un68_sum_axb_8 ));
    InMux I__1538 (
            .O(N__11150),
            .I(\POWERLED.mult1_un61_sum_cry_6 ));
    InMux I__1537 (
            .O(N__11147),
            .I(\POWERLED.mult1_un54_sum_cry_5 ));
    InMux I__1536 (
            .O(N__11144),
            .I(\POWERLED.mult1_un54_sum_cry_6 ));
    InMux I__1535 (
            .O(N__11141),
            .I(\POWERLED.mult1_un54_sum_cry_7 ));
    CascadeMux I__1534 (
            .O(N__11138),
            .I(N__11135));
    InMux I__1533 (
            .O(N__11135),
            .I(N__11132));
    LocalMux I__1532 (
            .O(N__11132),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    InMux I__1531 (
            .O(N__11129),
            .I(\POWERLED.mult1_un47_sum_cry_2 ));
    CascadeMux I__1530 (
            .O(N__11126),
            .I(N__11123));
    InMux I__1529 (
            .O(N__11123),
            .I(N__11120));
    LocalMux I__1528 (
            .O(N__11120),
            .I(\POWERLED.mult1_un47_sum_cry_4_s ));
    InMux I__1527 (
            .O(N__11117),
            .I(\POWERLED.mult1_un47_sum_cry_3 ));
    CascadeMux I__1526 (
            .O(N__11114),
            .I(N__11111));
    InMux I__1525 (
            .O(N__11111),
            .I(N__11108));
    LocalMux I__1524 (
            .O(N__11108),
            .I(\POWERLED.mult1_un47_sum_cry_5_s ));
    InMux I__1523 (
            .O(N__11105),
            .I(\POWERLED.mult1_un47_sum_cry_4 ));
    InMux I__1522 (
            .O(N__11102),
            .I(\POWERLED.mult1_un47_sum_cry_5 ));
    InMux I__1521 (
            .O(N__11099),
            .I(N__11096));
    LocalMux I__1520 (
            .O(N__11096),
            .I(\POWERLED.mult1_un54_sum_cry_7_THRU_CO ));
    InMux I__1519 (
            .O(N__11093),
            .I(\POWERLED.mult1_un47_sum_cry_6 ));
    CascadeMux I__1518 (
            .O(N__11090),
            .I(\POWERLED.un1_count_2_cry_15_THRU_CO_cascade_ ));
    CEMux I__1517 (
            .O(N__11087),
            .I(N__11084));
    LocalMux I__1516 (
            .O(N__11084),
            .I(N__11081));
    Span4Mux_v I__1515 (
            .O(N__11081),
            .I(N__11078));
    Odrv4 I__1514 (
            .O(N__11078),
            .I(\POWERLED.pwm_out_RNOZ0 ));
    InMux I__1513 (
            .O(N__11075),
            .I(N__11072));
    LocalMux I__1512 (
            .O(N__11072),
            .I(N__11069));
    Span4Mux_s3_v I__1511 (
            .O(N__11069),
            .I(N__11066));
    Odrv4 I__1510 (
            .O(N__11066),
            .I(vpp_ok));
    IoInMux I__1509 (
            .O(N__11063),
            .I(N__11060));
    LocalMux I__1508 (
            .O(N__11060),
            .I(N__11057));
    Span4Mux_s1_v I__1507 (
            .O(N__11057),
            .I(N__11054));
    Odrv4 I__1506 (
            .O(N__11054),
            .I(vddq_en));
    InMux I__1505 (
            .O(N__11051),
            .I(N__11048));
    LocalMux I__1504 (
            .O(N__11048),
            .I(N__11045));
    Span4Mux_v I__1503 (
            .O(N__11045),
            .I(N__11042));
    Span4Mux_h I__1502 (
            .O(N__11042),
            .I(N__11039));
    Odrv4 I__1501 (
            .O(N__11039),
            .I(gpio_fpga_soc_1));
    CascadeMux I__1500 (
            .O(N__11036),
            .I(\HDA_STRAP.N_5_0_cascade_ ));
    IoInMux I__1499 (
            .O(N__11033),
            .I(N__11030));
    LocalMux I__1498 (
            .O(N__11030),
            .I(N__11026));
    InMux I__1497 (
            .O(N__11029),
            .I(N__11022));
    Span4Mux_s0_h I__1496 (
            .O(N__11026),
            .I(N__11018));
    IoInMux I__1495 (
            .O(N__11025),
            .I(N__11015));
    LocalMux I__1494 (
            .O(N__11022),
            .I(N__11012));
    InMux I__1493 (
            .O(N__11021),
            .I(N__11009));
    Sp12to4 I__1492 (
            .O(N__11018),
            .I(N__11006));
    LocalMux I__1491 (
            .O(N__11015),
            .I(N__11003));
    Span4Mux_v I__1490 (
            .O(N__11012),
            .I(N__10998));
    LocalMux I__1489 (
            .O(N__11009),
            .I(N__10998));
    Span12Mux_v I__1488 (
            .O(N__11006),
            .I(N__10995));
    Span4Mux_s0_h I__1487 (
            .O(N__11003),
            .I(N__10990));
    Span4Mux_h I__1486 (
            .O(N__10998),
            .I(N__10990));
    Odrv12 I__1485 (
            .O(N__10995),
            .I(pch_pwrok));
    Odrv4 I__1484 (
            .O(N__10990),
            .I(pch_pwrok));
    CascadeMux I__1483 (
            .O(N__10985),
            .I(N__10982));
    InMux I__1482 (
            .O(N__10982),
            .I(N__10979));
    LocalMux I__1481 (
            .O(N__10979),
            .I(\HDA_STRAP.m14_ns_1 ));
    InMux I__1480 (
            .O(N__10976),
            .I(\POWERLED.mult1_un54_sum_cry_2 ));
    InMux I__1479 (
            .O(N__10973),
            .I(\POWERLED.mult1_un54_sum_cry_3 ));
    InMux I__1478 (
            .O(N__10970),
            .I(\POWERLED.mult1_un54_sum_cry_4 ));
    InMux I__1477 (
            .O(N__10967),
            .I(N__10964));
    LocalMux I__1476 (
            .O(N__10964),
            .I(N__10961));
    Odrv12 I__1475 (
            .O(N__10961),
            .I(\POWERLED.un1_count_2_9 ));
    CascadeMux I__1474 (
            .O(N__10958),
            .I(N__10955));
    InMux I__1473 (
            .O(N__10955),
            .I(N__10952));
    LocalMux I__1472 (
            .O(N__10952),
            .I(\POWERLED.count_i_9 ));
    InMux I__1471 (
            .O(N__10949),
            .I(N__10946));
    LocalMux I__1470 (
            .O(N__10946),
            .I(\POWERLED.un1_count_2_10 ));
    CascadeMux I__1469 (
            .O(N__10943),
            .I(N__10940));
    InMux I__1468 (
            .O(N__10940),
            .I(N__10937));
    LocalMux I__1467 (
            .O(N__10937),
            .I(\POWERLED.count_i_10 ));
    InMux I__1466 (
            .O(N__10934),
            .I(N__10931));
    LocalMux I__1465 (
            .O(N__10931),
            .I(N__10928));
    Odrv12 I__1464 (
            .O(N__10928),
            .I(\POWERLED.un1_count_2_11 ));
    CascadeMux I__1463 (
            .O(N__10925),
            .I(N__10922));
    InMux I__1462 (
            .O(N__10922),
            .I(N__10919));
    LocalMux I__1461 (
            .O(N__10919),
            .I(\POWERLED.count_i_11 ));
    InMux I__1460 (
            .O(N__10916),
            .I(N__10913));
    LocalMux I__1459 (
            .O(N__10913),
            .I(N__10910));
    Span4Mux_v I__1458 (
            .O(N__10910),
            .I(N__10907));
    Odrv4 I__1457 (
            .O(N__10907),
            .I(\POWERLED.un1_count_2_12 ));
    CascadeMux I__1456 (
            .O(N__10904),
            .I(N__10901));
    InMux I__1455 (
            .O(N__10901),
            .I(N__10898));
    LocalMux I__1454 (
            .O(N__10898),
            .I(N__10895));
    Odrv4 I__1453 (
            .O(N__10895),
            .I(\POWERLED.count_i_12 ));
    InMux I__1452 (
            .O(N__10892),
            .I(N__10889));
    LocalMux I__1451 (
            .O(N__10889),
            .I(N__10886));
    Span12Mux_s4_v I__1450 (
            .O(N__10886),
            .I(N__10883));
    Odrv12 I__1449 (
            .O(N__10883),
            .I(\POWERLED.un1_count_2_13 ));
    CascadeMux I__1448 (
            .O(N__10880),
            .I(N__10877));
    InMux I__1447 (
            .O(N__10877),
            .I(N__10874));
    LocalMux I__1446 (
            .O(N__10874),
            .I(\POWERLED.count_i_13 ));
    InMux I__1445 (
            .O(N__10871),
            .I(N__10868));
    LocalMux I__1444 (
            .O(N__10868),
            .I(N__10865));
    Span4Mux_v I__1443 (
            .O(N__10865),
            .I(N__10862));
    Odrv4 I__1442 (
            .O(N__10862),
            .I(\POWERLED.un1_count_2_14 ));
    CascadeMux I__1441 (
            .O(N__10859),
            .I(N__10856));
    InMux I__1440 (
            .O(N__10856),
            .I(N__10853));
    LocalMux I__1439 (
            .O(N__10853),
            .I(N__10850));
    Odrv4 I__1438 (
            .O(N__10850),
            .I(\POWERLED.count_i_14 ));
    InMux I__1437 (
            .O(N__10847),
            .I(N__10844));
    LocalMux I__1436 (
            .O(N__10844),
            .I(N__10841));
    Span4Mux_s3_v I__1435 (
            .O(N__10841),
            .I(N__10838));
    Odrv4 I__1434 (
            .O(N__10838),
            .I(\POWERLED.un1_count_2_15 ));
    CascadeMux I__1433 (
            .O(N__10835),
            .I(N__10832));
    InMux I__1432 (
            .O(N__10832),
            .I(N__10829));
    LocalMux I__1431 (
            .O(N__10829),
            .I(\POWERLED.count_i_15 ));
    InMux I__1430 (
            .O(N__10826),
            .I(bfn_2_15_0_));
    InMux I__1429 (
            .O(N__10823),
            .I(N__10820));
    LocalMux I__1428 (
            .O(N__10820),
            .I(\POWERLED.un1_count_2_cry_15_THRU_CO ));
    CascadeMux I__1427 (
            .O(N__10817),
            .I(N__10814));
    InMux I__1426 (
            .O(N__10814),
            .I(N__10811));
    LocalMux I__1425 (
            .O(N__10811),
            .I(\POWERLED.un1_count_2_1 ));
    InMux I__1424 (
            .O(N__10808),
            .I(N__10805));
    LocalMux I__1423 (
            .O(N__10805),
            .I(N__10802));
    Odrv4 I__1422 (
            .O(N__10802),
            .I(\POWERLED.count_i_1 ));
    InMux I__1421 (
            .O(N__10799),
            .I(N__10796));
    LocalMux I__1420 (
            .O(N__10796),
            .I(\POWERLED.un1_count_2_2 ));
    CascadeMux I__1419 (
            .O(N__10793),
            .I(N__10790));
    InMux I__1418 (
            .O(N__10790),
            .I(N__10787));
    LocalMux I__1417 (
            .O(N__10787),
            .I(\POWERLED.count_i_2 ));
    InMux I__1416 (
            .O(N__10784),
            .I(N__10781));
    LocalMux I__1415 (
            .O(N__10781),
            .I(N__10778));
    Odrv4 I__1414 (
            .O(N__10778),
            .I(\POWERLED.un1_count_2_3 ));
    CascadeMux I__1413 (
            .O(N__10775),
            .I(N__10772));
    InMux I__1412 (
            .O(N__10772),
            .I(N__10769));
    LocalMux I__1411 (
            .O(N__10769),
            .I(\POWERLED.count_i_3 ));
    CascadeMux I__1410 (
            .O(N__10766),
            .I(N__10763));
    InMux I__1409 (
            .O(N__10763),
            .I(N__10760));
    LocalMux I__1408 (
            .O(N__10760),
            .I(N__10757));
    Odrv4 I__1407 (
            .O(N__10757),
            .I(\POWERLED.count_i_4 ));
    InMux I__1406 (
            .O(N__10754),
            .I(N__10751));
    LocalMux I__1405 (
            .O(N__10751),
            .I(N__10748));
    Odrv12 I__1404 (
            .O(N__10748),
            .I(\POWERLED.un1_count_2_5 ));
    CascadeMux I__1403 (
            .O(N__10745),
            .I(N__10742));
    InMux I__1402 (
            .O(N__10742),
            .I(N__10739));
    LocalMux I__1401 (
            .O(N__10739),
            .I(\POWERLED.count_i_5 ));
    InMux I__1400 (
            .O(N__10736),
            .I(N__10733));
    LocalMux I__1399 (
            .O(N__10733),
            .I(N__10730));
    Odrv12 I__1398 (
            .O(N__10730),
            .I(\POWERLED.un1_count_2_6 ));
    CascadeMux I__1397 (
            .O(N__10727),
            .I(N__10724));
    InMux I__1396 (
            .O(N__10724),
            .I(N__10721));
    LocalMux I__1395 (
            .O(N__10721),
            .I(N__10718));
    Odrv4 I__1394 (
            .O(N__10718),
            .I(\POWERLED.count_i_6 ));
    InMux I__1393 (
            .O(N__10715),
            .I(N__10712));
    LocalMux I__1392 (
            .O(N__10712),
            .I(N__10709));
    Odrv4 I__1391 (
            .O(N__10709),
            .I(\POWERLED.un1_count_2_7 ));
    CascadeMux I__1390 (
            .O(N__10706),
            .I(N__10703));
    InMux I__1389 (
            .O(N__10703),
            .I(N__10700));
    LocalMux I__1388 (
            .O(N__10700),
            .I(N__10697));
    Odrv4 I__1387 (
            .O(N__10697),
            .I(\POWERLED.count_i_7 ));
    InMux I__1386 (
            .O(N__10694),
            .I(N__10691));
    LocalMux I__1385 (
            .O(N__10691),
            .I(N__10688));
    Odrv12 I__1384 (
            .O(N__10688),
            .I(\POWERLED.un1_count_2_8 ));
    CascadeMux I__1383 (
            .O(N__10685),
            .I(N__10682));
    InMux I__1382 (
            .O(N__10682),
            .I(N__10679));
    LocalMux I__1381 (
            .O(N__10679),
            .I(\POWERLED.count_i_8 ));
    CascadeMux I__1380 (
            .O(N__10676),
            .I(N__10673));
    InMux I__1379 (
            .O(N__10673),
            .I(N__10670));
    LocalMux I__1378 (
            .O(N__10670),
            .I(\POWERLED.mult1_un152_sum_cry_3_s ));
    InMux I__1377 (
            .O(N__10667),
            .I(\POWERLED.mult1_un152_sum_cry_2 ));
    CascadeMux I__1376 (
            .O(N__10664),
            .I(N__10661));
    InMux I__1375 (
            .O(N__10661),
            .I(N__10658));
    LocalMux I__1374 (
            .O(N__10658),
            .I(\POWERLED.mult1_un145_sum_cry_3_s ));
    InMux I__1373 (
            .O(N__10655),
            .I(N__10652));
    LocalMux I__1372 (
            .O(N__10652),
            .I(\POWERLED.mult1_un152_sum_cry_4_s ));
    InMux I__1371 (
            .O(N__10649),
            .I(\POWERLED.mult1_un152_sum_cry_3 ));
    InMux I__1370 (
            .O(N__10646),
            .I(N__10643));
    LocalMux I__1369 (
            .O(N__10643),
            .I(\POWERLED.mult1_un145_sum_cry_4_s ));
    CascadeMux I__1368 (
            .O(N__10640),
            .I(N__10637));
    InMux I__1367 (
            .O(N__10637),
            .I(N__10634));
    LocalMux I__1366 (
            .O(N__10634),
            .I(\POWERLED.mult1_un152_sum_cry_5_s ));
    InMux I__1365 (
            .O(N__10631),
            .I(\POWERLED.mult1_un152_sum_cry_4 ));
    CascadeMux I__1364 (
            .O(N__10628),
            .I(N__10623));
    InMux I__1363 (
            .O(N__10627),
            .I(N__10619));
    InMux I__1362 (
            .O(N__10626),
            .I(N__10614));
    InMux I__1361 (
            .O(N__10623),
            .I(N__10614));
    InMux I__1360 (
            .O(N__10622),
            .I(N__10611));
    LocalMux I__1359 (
            .O(N__10619),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__1358 (
            .O(N__10614),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__1357 (
            .O(N__10611),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    CascadeMux I__1356 (
            .O(N__10604),
            .I(N__10601));
    InMux I__1355 (
            .O(N__10601),
            .I(N__10598));
    LocalMux I__1354 (
            .O(N__10598),
            .I(\POWERLED.mult1_un145_sum_cry_5_s ));
    InMux I__1353 (
            .O(N__10595),
            .I(N__10592));
    LocalMux I__1352 (
            .O(N__10592),
            .I(\POWERLED.mult1_un152_sum_cry_6_s ));
    InMux I__1351 (
            .O(N__10589),
            .I(\POWERLED.mult1_un152_sum_cry_5 ));
    InMux I__1350 (
            .O(N__10586),
            .I(N__10583));
    LocalMux I__1349 (
            .O(N__10583),
            .I(\POWERLED.mult1_un145_sum_cry_6_s ));
    CascadeMux I__1348 (
            .O(N__10580),
            .I(N__10576));
    CascadeMux I__1347 (
            .O(N__10579),
            .I(N__10572));
    InMux I__1346 (
            .O(N__10576),
            .I(N__10565));
    InMux I__1345 (
            .O(N__10575),
            .I(N__10565));
    InMux I__1344 (
            .O(N__10572),
            .I(N__10565));
    LocalMux I__1343 (
            .O(N__10565),
            .I(\POWERLED.mult1_un145_sum_i_0_8 ));
    InMux I__1342 (
            .O(N__10562),
            .I(N__10559));
    LocalMux I__1341 (
            .O(N__10559),
            .I(\POWERLED.mult1_un159_sum_axb_7 ));
    InMux I__1340 (
            .O(N__10556),
            .I(\POWERLED.mult1_un152_sum_cry_6 ));
    InMux I__1339 (
            .O(N__10553),
            .I(N__10550));
    LocalMux I__1338 (
            .O(N__10550),
            .I(\POWERLED.mult1_un152_sum_axb_8 ));
    InMux I__1337 (
            .O(N__10547),
            .I(\POWERLED.mult1_un152_sum_cry_7 ));
    CascadeMux I__1336 (
            .O(N__10544),
            .I(N__10539));
    InMux I__1335 (
            .O(N__10543),
            .I(N__10535));
    InMux I__1334 (
            .O(N__10542),
            .I(N__10530));
    InMux I__1333 (
            .O(N__10539),
            .I(N__10530));
    InMux I__1332 (
            .O(N__10538),
            .I(N__10527));
    LocalMux I__1331 (
            .O(N__10535),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__1330 (
            .O(N__10530),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__1329 (
            .O(N__10527),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    CascadeMux I__1328 (
            .O(N__10520),
            .I(\POWERLED.mult1_un152_sum_s_8_cascade_ ));
    CascadeMux I__1327 (
            .O(N__10517),
            .I(N__10513));
    CascadeMux I__1326 (
            .O(N__10516),
            .I(N__10509));
    InMux I__1325 (
            .O(N__10513),
            .I(N__10502));
    InMux I__1324 (
            .O(N__10512),
            .I(N__10502));
    InMux I__1323 (
            .O(N__10509),
            .I(N__10502));
    LocalMux I__1322 (
            .O(N__10502),
            .I(\POWERLED.mult1_un152_sum_i_0_8 ));
    CascadeMux I__1321 (
            .O(N__10499),
            .I(N__10496));
    InMux I__1320 (
            .O(N__10496),
            .I(N__10493));
    LocalMux I__1319 (
            .O(N__10493),
            .I(\POWERLED.un1_count_2_0 ));
    InMux I__1318 (
            .O(N__10490),
            .I(N__10487));
    LocalMux I__1317 (
            .O(N__10487),
            .I(\POWERLED.count_i_0_0 ));
    CascadeMux I__1316 (
            .O(N__10484),
            .I(N__10481));
    InMux I__1315 (
            .O(N__10481),
            .I(N__10478));
    LocalMux I__1314 (
            .O(N__10478),
            .I(\POWERLED.mult1_un138_sum_i_0_8 ));
    InMux I__1313 (
            .O(N__10475),
            .I(\POWERLED.mult1_un145_sum_cry_2 ));
    InMux I__1312 (
            .O(N__10472),
            .I(N__10468));
    InMux I__1311 (
            .O(N__10471),
            .I(N__10465));
    LocalMux I__1310 (
            .O(N__10468),
            .I(\POWERLED.mult1_un138_sum_cry_3_s ));
    LocalMux I__1309 (
            .O(N__10465),
            .I(\POWERLED.mult1_un138_sum_cry_3_s ));
    CascadeMux I__1308 (
            .O(N__10460),
            .I(N__10457));
    InMux I__1307 (
            .O(N__10457),
            .I(N__10454));
    LocalMux I__1306 (
            .O(N__10454),
            .I(\POWERLED.mult1_un145_sum_axb_4_l_fx ));
    InMux I__1305 (
            .O(N__10451),
            .I(\POWERLED.mult1_un145_sum_cry_3 ));
    InMux I__1304 (
            .O(N__10448),
            .I(N__10445));
    LocalMux I__1303 (
            .O(N__10445),
            .I(N__10442));
    Odrv4 I__1302 (
            .O(N__10442),
            .I(\POWERLED.mult1_un138_sum_cry_4_s ));
    InMux I__1301 (
            .O(N__10439),
            .I(\POWERLED.mult1_un145_sum_cry_4 ));
    CascadeMux I__1300 (
            .O(N__10436),
            .I(N__10433));
    InMux I__1299 (
            .O(N__10433),
            .I(N__10430));
    LocalMux I__1298 (
            .O(N__10430),
            .I(\POWERLED.mult1_un138_sum_cry_5_s ));
    InMux I__1297 (
            .O(N__10427),
            .I(\POWERLED.mult1_un145_sum_cry_5 ));
    InMux I__1296 (
            .O(N__10424),
            .I(\POWERLED.mult1_un145_sum_cry_6 ));
    InMux I__1295 (
            .O(N__10421),
            .I(N__10418));
    LocalMux I__1294 (
            .O(N__10418),
            .I(\POWERLED.mult1_un145_sum_axb_8 ));
    InMux I__1293 (
            .O(N__10415),
            .I(\POWERLED.mult1_un145_sum_cry_7 ));
    CascadeMux I__1292 (
            .O(N__10412),
            .I(\POWERLED.mult1_un145_sum_s_8_cascade_ ));
    InMux I__1291 (
            .O(N__10409),
            .I(N__10406));
    LocalMux I__1290 (
            .O(N__10406),
            .I(N__10403));
    Odrv4 I__1289 (
            .O(N__10403),
            .I(\POWERLED.mult1_un145_sum_i ));
    CascadeMux I__1288 (
            .O(N__10400),
            .I(\POWERLED.mult1_un117_sum_s_8_cascade_ ));
    CascadeMux I__1287 (
            .O(N__10397),
            .I(N__10393));
    CascadeMux I__1286 (
            .O(N__10396),
            .I(N__10389));
    InMux I__1285 (
            .O(N__10393),
            .I(N__10382));
    InMux I__1284 (
            .O(N__10392),
            .I(N__10382));
    InMux I__1283 (
            .O(N__10389),
            .I(N__10382));
    LocalMux I__1282 (
            .O(N__10382),
            .I(\POWERLED.mult1_un117_sum_i_0_8 ));
    CascadeMux I__1281 (
            .O(N__10379),
            .I(N__10374));
    InMux I__1280 (
            .O(N__10378),
            .I(N__10370));
    InMux I__1279 (
            .O(N__10377),
            .I(N__10365));
    InMux I__1278 (
            .O(N__10374),
            .I(N__10365));
    InMux I__1277 (
            .O(N__10373),
            .I(N__10362));
    LocalMux I__1276 (
            .O(N__10370),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__1275 (
            .O(N__10365),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__1274 (
            .O(N__10362),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    CascadeMux I__1273 (
            .O(N__10355),
            .I(N__10350));
    InMux I__1272 (
            .O(N__10354),
            .I(N__10346));
    InMux I__1271 (
            .O(N__10353),
            .I(N__10341));
    InMux I__1270 (
            .O(N__10350),
            .I(N__10341));
    InMux I__1269 (
            .O(N__10349),
            .I(N__10338));
    LocalMux I__1268 (
            .O(N__10346),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__1267 (
            .O(N__10341),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__1266 (
            .O(N__10338),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    InMux I__1265 (
            .O(N__10331),
            .I(N__10328));
    LocalMux I__1264 (
            .O(N__10328),
            .I(N__10325));
    Odrv4 I__1263 (
            .O(N__10325),
            .I(\POWERLED.mult1_un131_sum_i ));
    InMux I__1262 (
            .O(N__10322),
            .I(N__10318));
    CascadeMux I__1261 (
            .O(N__10321),
            .I(N__10314));
    LocalMux I__1260 (
            .O(N__10318),
            .I(N__10310));
    InMux I__1259 (
            .O(N__10317),
            .I(N__10305));
    InMux I__1258 (
            .O(N__10314),
            .I(N__10305));
    InMux I__1257 (
            .O(N__10313),
            .I(N__10302));
    Odrv4 I__1256 (
            .O(N__10310),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__1255 (
            .O(N__10305),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__1254 (
            .O(N__10302),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    InMux I__1253 (
            .O(N__10295),
            .I(N__10292));
    LocalMux I__1252 (
            .O(N__10292),
            .I(N__10289));
    Span4Mux_s1_h I__1251 (
            .O(N__10289),
            .I(N__10286));
    Odrv4 I__1250 (
            .O(N__10286),
            .I(\POWERLED.mult1_un89_sum_i ));
    CascadeMux I__1249 (
            .O(N__10283),
            .I(N__10280));
    InMux I__1248 (
            .O(N__10280),
            .I(N__10277));
    LocalMux I__1247 (
            .O(N__10277),
            .I(\POWERLED.mult1_un117_sum_cry_3_s ));
    InMux I__1246 (
            .O(N__10274),
            .I(\POWERLED.mult1_un117_sum_cry_2 ));
    CascadeMux I__1245 (
            .O(N__10271),
            .I(N__10268));
    InMux I__1244 (
            .O(N__10268),
            .I(N__10265));
    LocalMux I__1243 (
            .O(N__10265),
            .I(\POWERLED.mult1_un110_sum_cry_3_s ));
    InMux I__1242 (
            .O(N__10262),
            .I(N__10259));
    LocalMux I__1241 (
            .O(N__10259),
            .I(\POWERLED.mult1_un117_sum_cry_4_s ));
    InMux I__1240 (
            .O(N__10256),
            .I(\POWERLED.mult1_un117_sum_cry_3 ));
    InMux I__1239 (
            .O(N__10253),
            .I(N__10250));
    LocalMux I__1238 (
            .O(N__10250),
            .I(\POWERLED.mult1_un110_sum_cry_4_s ));
    CascadeMux I__1237 (
            .O(N__10247),
            .I(N__10244));
    InMux I__1236 (
            .O(N__10244),
            .I(N__10241));
    LocalMux I__1235 (
            .O(N__10241),
            .I(\POWERLED.mult1_un117_sum_cry_5_s ));
    InMux I__1234 (
            .O(N__10238),
            .I(\POWERLED.mult1_un117_sum_cry_4 ));
    CascadeMux I__1233 (
            .O(N__10235),
            .I(N__10230));
    InMux I__1232 (
            .O(N__10234),
            .I(N__10226));
    InMux I__1231 (
            .O(N__10233),
            .I(N__10221));
    InMux I__1230 (
            .O(N__10230),
            .I(N__10221));
    InMux I__1229 (
            .O(N__10229),
            .I(N__10218));
    LocalMux I__1228 (
            .O(N__10226),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__1227 (
            .O(N__10221),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__1226 (
            .O(N__10218),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    CascadeMux I__1225 (
            .O(N__10211),
            .I(N__10208));
    InMux I__1224 (
            .O(N__10208),
            .I(N__10205));
    LocalMux I__1223 (
            .O(N__10205),
            .I(\POWERLED.mult1_un110_sum_cry_5_s ));
    InMux I__1222 (
            .O(N__10202),
            .I(N__10199));
    LocalMux I__1221 (
            .O(N__10199),
            .I(\POWERLED.mult1_un117_sum_cry_6_s ));
    InMux I__1220 (
            .O(N__10196),
            .I(\POWERLED.mult1_un117_sum_cry_5 ));
    InMux I__1219 (
            .O(N__10193),
            .I(N__10190));
    LocalMux I__1218 (
            .O(N__10190),
            .I(\POWERLED.mult1_un110_sum_cry_6_s ));
    CascadeMux I__1217 (
            .O(N__10187),
            .I(N__10183));
    CascadeMux I__1216 (
            .O(N__10186),
            .I(N__10179));
    InMux I__1215 (
            .O(N__10183),
            .I(N__10172));
    InMux I__1214 (
            .O(N__10182),
            .I(N__10172));
    InMux I__1213 (
            .O(N__10179),
            .I(N__10172));
    LocalMux I__1212 (
            .O(N__10172),
            .I(\POWERLED.mult1_un110_sum_i_0_8 ));
    InMux I__1211 (
            .O(N__10169),
            .I(N__10166));
    LocalMux I__1210 (
            .O(N__10166),
            .I(\POWERLED.mult1_un124_sum_axb_8 ));
    InMux I__1209 (
            .O(N__10163),
            .I(\POWERLED.mult1_un117_sum_cry_6 ));
    InMux I__1208 (
            .O(N__10160),
            .I(N__10157));
    LocalMux I__1207 (
            .O(N__10157),
            .I(\POWERLED.mult1_un117_sum_axb_8 ));
    InMux I__1206 (
            .O(N__10154),
            .I(\POWERLED.mult1_un117_sum_cry_7 ));
    InMux I__1205 (
            .O(N__10151),
            .I(\POWERLED.mult1_un68_sum_cry_7 ));
    CascadeMux I__1204 (
            .O(N__10148),
            .I(N__10144));
    CascadeMux I__1203 (
            .O(N__10147),
            .I(N__10140));
    InMux I__1202 (
            .O(N__10144),
            .I(N__10133));
    InMux I__1201 (
            .O(N__10143),
            .I(N__10133));
    InMux I__1200 (
            .O(N__10140),
            .I(N__10133));
    LocalMux I__1199 (
            .O(N__10133),
            .I(\POWERLED.mult1_un68_sum_i_0_8 ));
    InMux I__1198 (
            .O(N__10130),
            .I(N__10126));
    CascadeMux I__1197 (
            .O(N__10129),
            .I(N__10122));
    LocalMux I__1196 (
            .O(N__10126),
            .I(N__10118));
    InMux I__1195 (
            .O(N__10125),
            .I(N__10113));
    InMux I__1194 (
            .O(N__10122),
            .I(N__10113));
    InMux I__1193 (
            .O(N__10121),
            .I(N__10110));
    Odrv4 I__1192 (
            .O(N__10118),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__1191 (
            .O(N__10113),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__1190 (
            .O(N__10110),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    InMux I__1189 (
            .O(N__10103),
            .I(N__10099));
    CascadeMux I__1188 (
            .O(N__10102),
            .I(N__10095));
    LocalMux I__1187 (
            .O(N__10099),
            .I(N__10091));
    InMux I__1186 (
            .O(N__10098),
            .I(N__10086));
    InMux I__1185 (
            .O(N__10095),
            .I(N__10086));
    InMux I__1184 (
            .O(N__10094),
            .I(N__10083));
    Odrv4 I__1183 (
            .O(N__10091),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__1182 (
            .O(N__10086),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__1181 (
            .O(N__10083),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    CascadeMux I__1180 (
            .O(N__10076),
            .I(N__10071));
    InMux I__1179 (
            .O(N__10075),
            .I(N__10066));
    InMux I__1178 (
            .O(N__10074),
            .I(N__10061));
    InMux I__1177 (
            .O(N__10071),
            .I(N__10061));
    InMux I__1176 (
            .O(N__10070),
            .I(N__10058));
    InMux I__1175 (
            .O(N__10069),
            .I(N__10055));
    LocalMux I__1174 (
            .O(N__10066),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__1173 (
            .O(N__10061),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__1172 (
            .O(N__10058),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__1171 (
            .O(N__10055),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    InMux I__1170 (
            .O(N__10046),
            .I(N__10042));
    CascadeMux I__1169 (
            .O(N__10045),
            .I(N__10038));
    LocalMux I__1168 (
            .O(N__10042),
            .I(N__10034));
    InMux I__1167 (
            .O(N__10041),
            .I(N__10029));
    InMux I__1166 (
            .O(N__10038),
            .I(N__10029));
    InMux I__1165 (
            .O(N__10037),
            .I(N__10026));
    Odrv4 I__1164 (
            .O(N__10034),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__1163 (
            .O(N__10029),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__1162 (
            .O(N__10026),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    InMux I__1161 (
            .O(N__10019),
            .I(N__10016));
    LocalMux I__1160 (
            .O(N__10016),
            .I(\POWERLED.mult1_un103_sum_i ));
    CascadeMux I__1159 (
            .O(N__10013),
            .I(N__10008));
    InMux I__1158 (
            .O(N__10012),
            .I(N__10004));
    InMux I__1157 (
            .O(N__10011),
            .I(N__9999));
    InMux I__1156 (
            .O(N__10008),
            .I(N__9999));
    InMux I__1155 (
            .O(N__10007),
            .I(N__9996));
    LocalMux I__1154 (
            .O(N__10004),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__1153 (
            .O(N__9999),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__1152 (
            .O(N__9996),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    InMux I__1151 (
            .O(N__9989),
            .I(N__9986));
    LocalMux I__1150 (
            .O(N__9986),
            .I(\POWERLED.mult1_un82_sum_axb_8 ));
    InMux I__1149 (
            .O(N__9983),
            .I(\POWERLED.mult1_un75_sum_cry_6 ));
    InMux I__1148 (
            .O(N__9980),
            .I(\POWERLED.mult1_un75_sum_cry_7 ));
    CascadeMux I__1147 (
            .O(N__9977),
            .I(\POWERLED.mult1_un75_sum_s_8_cascade_ ));
    CascadeMux I__1146 (
            .O(N__9974),
            .I(N__9970));
    CascadeMux I__1145 (
            .O(N__9973),
            .I(N__9966));
    InMux I__1144 (
            .O(N__9970),
            .I(N__9959));
    InMux I__1143 (
            .O(N__9969),
            .I(N__9959));
    InMux I__1142 (
            .O(N__9966),
            .I(N__9959));
    LocalMux I__1141 (
            .O(N__9959),
            .I(\POWERLED.mult1_un75_sum_i_0_8 ));
    CascadeMux I__1140 (
            .O(N__9956),
            .I(N__9953));
    InMux I__1139 (
            .O(N__9953),
            .I(N__9950));
    LocalMux I__1138 (
            .O(N__9950),
            .I(\POWERLED.mult1_un68_sum_cry_3_s ));
    InMux I__1137 (
            .O(N__9947),
            .I(\POWERLED.mult1_un68_sum_cry_2 ));
    InMux I__1136 (
            .O(N__9944),
            .I(N__9941));
    LocalMux I__1135 (
            .O(N__9941),
            .I(\POWERLED.mult1_un68_sum_cry_4_s ));
    InMux I__1134 (
            .O(N__9938),
            .I(\POWERLED.mult1_un68_sum_cry_3 ));
    CascadeMux I__1133 (
            .O(N__9935),
            .I(N__9932));
    InMux I__1132 (
            .O(N__9932),
            .I(N__9929));
    LocalMux I__1131 (
            .O(N__9929),
            .I(\POWERLED.mult1_un68_sum_cry_5_s ));
    InMux I__1130 (
            .O(N__9926),
            .I(\POWERLED.mult1_un68_sum_cry_4 ));
    InMux I__1129 (
            .O(N__9923),
            .I(N__9920));
    LocalMux I__1128 (
            .O(N__9920),
            .I(\POWERLED.mult1_un68_sum_cry_6_s ));
    InMux I__1127 (
            .O(N__9917),
            .I(\POWERLED.mult1_un68_sum_cry_5 ));
    InMux I__1126 (
            .O(N__9914),
            .I(N__9911));
    LocalMux I__1125 (
            .O(N__9911),
            .I(\POWERLED.mult1_un75_sum_axb_8 ));
    InMux I__1124 (
            .O(N__9908),
            .I(\POWERLED.mult1_un68_sum_cry_6 ));
    InMux I__1123 (
            .O(N__9905),
            .I(N__9902));
    LocalMux I__1122 (
            .O(N__9902),
            .I(\POWERLED.mult1_un89_sum_axb_8 ));
    InMux I__1121 (
            .O(N__9899),
            .I(\POWERLED.mult1_un82_sum_cry_6 ));
    InMux I__1120 (
            .O(N__9896),
            .I(\POWERLED.mult1_un82_sum_cry_7 ));
    CascadeMux I__1119 (
            .O(N__9893),
            .I(\POWERLED.mult1_un82_sum_s_8_cascade_ ));
    CascadeMux I__1118 (
            .O(N__9890),
            .I(N__9886));
    CascadeMux I__1117 (
            .O(N__9889),
            .I(N__9882));
    InMux I__1116 (
            .O(N__9886),
            .I(N__9875));
    InMux I__1115 (
            .O(N__9885),
            .I(N__9875));
    InMux I__1114 (
            .O(N__9882),
            .I(N__9875));
    LocalMux I__1113 (
            .O(N__9875),
            .I(\POWERLED.mult1_un82_sum_i_0_8 ));
    CascadeMux I__1112 (
            .O(N__9872),
            .I(N__9869));
    InMux I__1111 (
            .O(N__9869),
            .I(N__9866));
    LocalMux I__1110 (
            .O(N__9866),
            .I(\POWERLED.mult1_un75_sum_cry_3_s ));
    InMux I__1109 (
            .O(N__9863),
            .I(\POWERLED.mult1_un75_sum_cry_2 ));
    InMux I__1108 (
            .O(N__9860),
            .I(N__9857));
    LocalMux I__1107 (
            .O(N__9857),
            .I(\POWERLED.mult1_un75_sum_cry_4_s ));
    InMux I__1106 (
            .O(N__9854),
            .I(\POWERLED.mult1_un75_sum_cry_3 ));
    CascadeMux I__1105 (
            .O(N__9851),
            .I(N__9848));
    InMux I__1104 (
            .O(N__9848),
            .I(N__9845));
    LocalMux I__1103 (
            .O(N__9845),
            .I(\POWERLED.mult1_un75_sum_cry_5_s ));
    InMux I__1102 (
            .O(N__9842),
            .I(\POWERLED.mult1_un75_sum_cry_4 ));
    InMux I__1101 (
            .O(N__9839),
            .I(N__9836));
    LocalMux I__1100 (
            .O(N__9836),
            .I(\POWERLED.mult1_un75_sum_cry_6_s ));
    InMux I__1099 (
            .O(N__9833),
            .I(\POWERLED.mult1_un75_sum_cry_5 ));
    InMux I__1098 (
            .O(N__9830),
            .I(N__9826));
    InMux I__1097 (
            .O(N__9829),
            .I(N__9823));
    LocalMux I__1096 (
            .O(N__9826),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    LocalMux I__1095 (
            .O(N__9823),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    InMux I__1094 (
            .O(N__9818),
            .I(\PCH_PWRGD.un1_count_1_cry_12 ));
    InMux I__1093 (
            .O(N__9815),
            .I(N__9811));
    InMux I__1092 (
            .O(N__9814),
            .I(N__9808));
    LocalMux I__1091 (
            .O(N__9811),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    LocalMux I__1090 (
            .O(N__9808),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    InMux I__1089 (
            .O(N__9803),
            .I(\PCH_PWRGD.un1_count_1_cry_13 ));
    InMux I__1088 (
            .O(N__9800),
            .I(bfn_2_4_0_));
    CascadeMux I__1087 (
            .O(N__9797),
            .I(N__9793));
    InMux I__1086 (
            .O(N__9796),
            .I(N__9790));
    InMux I__1085 (
            .O(N__9793),
            .I(N__9787));
    LocalMux I__1084 (
            .O(N__9790),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    LocalMux I__1083 (
            .O(N__9787),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    CEMux I__1082 (
            .O(N__9782),
            .I(N__9779));
    LocalMux I__1081 (
            .O(N__9779),
            .I(N__9776));
    Span4Mux_v I__1080 (
            .O(N__9776),
            .I(N__9773));
    Odrv4 I__1079 (
            .O(N__9773),
            .I(\PCH_PWRGD.N_65_3 ));
    SRMux I__1078 (
            .O(N__9770),
            .I(N__9765));
    SRMux I__1077 (
            .O(N__9769),
            .I(N__9762));
    SRMux I__1076 (
            .O(N__9768),
            .I(N__9759));
    LocalMux I__1075 (
            .O(N__9765),
            .I(\PCH_PWRGD.curr_state_RNI7N705Z0Z_0 ));
    LocalMux I__1074 (
            .O(N__9762),
            .I(\PCH_PWRGD.curr_state_RNI7N705Z0Z_0 ));
    LocalMux I__1073 (
            .O(N__9759),
            .I(\PCH_PWRGD.curr_state_RNI7N705Z0Z_0 ));
    CascadeMux I__1072 (
            .O(N__9752),
            .I(N__9749));
    InMux I__1071 (
            .O(N__9749),
            .I(N__9746));
    LocalMux I__1070 (
            .O(N__9746),
            .I(\POWERLED.mult1_un82_sum_cry_3_s ));
    InMux I__1069 (
            .O(N__9743),
            .I(\POWERLED.mult1_un82_sum_cry_2 ));
    InMux I__1068 (
            .O(N__9740),
            .I(N__9737));
    LocalMux I__1067 (
            .O(N__9737),
            .I(\POWERLED.mult1_un82_sum_cry_4_s ));
    InMux I__1066 (
            .O(N__9734),
            .I(\POWERLED.mult1_un82_sum_cry_3 ));
    CascadeMux I__1065 (
            .O(N__9731),
            .I(N__9728));
    InMux I__1064 (
            .O(N__9728),
            .I(N__9725));
    LocalMux I__1063 (
            .O(N__9725),
            .I(\POWERLED.mult1_un82_sum_cry_5_s ));
    InMux I__1062 (
            .O(N__9722),
            .I(\POWERLED.mult1_un82_sum_cry_4 ));
    InMux I__1061 (
            .O(N__9719),
            .I(N__9716));
    LocalMux I__1060 (
            .O(N__9716),
            .I(\POWERLED.mult1_un82_sum_cry_6_s ));
    InMux I__1059 (
            .O(N__9713),
            .I(\POWERLED.mult1_un82_sum_cry_5 ));
    InMux I__1058 (
            .O(N__9710),
            .I(N__9706));
    InMux I__1057 (
            .O(N__9709),
            .I(N__9703));
    LocalMux I__1056 (
            .O(N__9706),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    LocalMux I__1055 (
            .O(N__9703),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    InMux I__1054 (
            .O(N__9698),
            .I(\PCH_PWRGD.un1_count_1_cry_4 ));
    InMux I__1053 (
            .O(N__9695),
            .I(N__9691));
    InMux I__1052 (
            .O(N__9694),
            .I(N__9688));
    LocalMux I__1051 (
            .O(N__9691),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    LocalMux I__1050 (
            .O(N__9688),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    InMux I__1049 (
            .O(N__9683),
            .I(\PCH_PWRGD.un1_count_1_cry_5 ));
    CascadeMux I__1048 (
            .O(N__9680),
            .I(N__9676));
    InMux I__1047 (
            .O(N__9679),
            .I(N__9673));
    InMux I__1046 (
            .O(N__9676),
            .I(N__9670));
    LocalMux I__1045 (
            .O(N__9673),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    LocalMux I__1044 (
            .O(N__9670),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    InMux I__1043 (
            .O(N__9665),
            .I(\PCH_PWRGD.un1_count_1_cry_6 ));
    InMux I__1042 (
            .O(N__9662),
            .I(N__9658));
    InMux I__1041 (
            .O(N__9661),
            .I(N__9655));
    LocalMux I__1040 (
            .O(N__9658),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    LocalMux I__1039 (
            .O(N__9655),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    InMux I__1038 (
            .O(N__9650),
            .I(bfn_2_3_0_));
    InMux I__1037 (
            .O(N__9647),
            .I(N__9643));
    InMux I__1036 (
            .O(N__9646),
            .I(N__9640));
    LocalMux I__1035 (
            .O(N__9643),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    LocalMux I__1034 (
            .O(N__9640),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    InMux I__1033 (
            .O(N__9635),
            .I(\PCH_PWRGD.un1_count_1_cry_8 ));
    CascadeMux I__1032 (
            .O(N__9632),
            .I(N__9628));
    InMux I__1031 (
            .O(N__9631),
            .I(N__9625));
    InMux I__1030 (
            .O(N__9628),
            .I(N__9622));
    LocalMux I__1029 (
            .O(N__9625),
            .I(\PCH_PWRGD.countZ0Z_10 ));
    LocalMux I__1028 (
            .O(N__9622),
            .I(\PCH_PWRGD.countZ0Z_10 ));
    InMux I__1027 (
            .O(N__9617),
            .I(\PCH_PWRGD.un1_count_1_cry_9 ));
    CascadeMux I__1026 (
            .O(N__9614),
            .I(N__9610));
    InMux I__1025 (
            .O(N__9613),
            .I(N__9607));
    InMux I__1024 (
            .O(N__9610),
            .I(N__9604));
    LocalMux I__1023 (
            .O(N__9607),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    LocalMux I__1022 (
            .O(N__9604),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    InMux I__1021 (
            .O(N__9599),
            .I(\PCH_PWRGD.un1_count_1_cry_10 ));
    InMux I__1020 (
            .O(N__9596),
            .I(N__9592));
    InMux I__1019 (
            .O(N__9595),
            .I(N__9589));
    LocalMux I__1018 (
            .O(N__9592),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    LocalMux I__1017 (
            .O(N__9589),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    InMux I__1016 (
            .O(N__9584),
            .I(\PCH_PWRGD.un1_count_1_cry_11 ));
    InMux I__1015 (
            .O(N__9581),
            .I(N__9578));
    LocalMux I__1014 (
            .O(N__9578),
            .I(N__9575));
    Odrv12 I__1013 (
            .O(N__9575),
            .I(\POWERLED.mult1_un96_sum_i ));
    InMux I__1012 (
            .O(N__9572),
            .I(N__9569));
    LocalMux I__1011 (
            .O(N__9569),
            .I(N__9565));
    CascadeMux I__1010 (
            .O(N__9568),
            .I(N__9561));
    Span12Mux_s4_v I__1009 (
            .O(N__9565),
            .I(N__9557));
    InMux I__1008 (
            .O(N__9564),
            .I(N__9552));
    InMux I__1007 (
            .O(N__9561),
            .I(N__9552));
    InMux I__1006 (
            .O(N__9560),
            .I(N__9549));
    Odrv12 I__1005 (
            .O(N__9557),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__1004 (
            .O(N__9552),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__1003 (
            .O(N__9549),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    IoInMux I__1002 (
            .O(N__9542),
            .I(N__9539));
    LocalMux I__1001 (
            .O(N__9539),
            .I(N__9536));
    Odrv4 I__1000 (
            .O(N__9536),
            .I(pwrbtn_led));
    CascadeMux I__999 (
            .O(N__9533),
            .I(N__9529));
    InMux I__998 (
            .O(N__9532),
            .I(N__9526));
    InMux I__997 (
            .O(N__9529),
            .I(N__9523));
    LocalMux I__996 (
            .O(N__9526),
            .I(N__9518));
    LocalMux I__995 (
            .O(N__9523),
            .I(N__9518));
    Odrv4 I__994 (
            .O(N__9518),
            .I(\PCH_PWRGD.un1_curr_state10_0 ));
    InMux I__993 (
            .O(N__9515),
            .I(N__9511));
    InMux I__992 (
            .O(N__9514),
            .I(N__9508));
    LocalMux I__991 (
            .O(N__9511),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    LocalMux I__990 (
            .O(N__9508),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    InMux I__989 (
            .O(N__9503),
            .I(N__9499));
    InMux I__988 (
            .O(N__9502),
            .I(N__9496));
    LocalMux I__987 (
            .O(N__9499),
            .I(\PCH_PWRGD.countZ0Z_1 ));
    LocalMux I__986 (
            .O(N__9496),
            .I(\PCH_PWRGD.countZ0Z_1 ));
    InMux I__985 (
            .O(N__9491),
            .I(\PCH_PWRGD.un1_count_1_cry_0 ));
    InMux I__984 (
            .O(N__9488),
            .I(N__9484));
    InMux I__983 (
            .O(N__9487),
            .I(N__9481));
    LocalMux I__982 (
            .O(N__9484),
            .I(\PCH_PWRGD.countZ0Z_2 ));
    LocalMux I__981 (
            .O(N__9481),
            .I(\PCH_PWRGD.countZ0Z_2 ));
    InMux I__980 (
            .O(N__9476),
            .I(\PCH_PWRGD.un1_count_1_cry_1 ));
    InMux I__979 (
            .O(N__9473),
            .I(N__9469));
    InMux I__978 (
            .O(N__9472),
            .I(N__9466));
    LocalMux I__977 (
            .O(N__9469),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    LocalMux I__976 (
            .O(N__9466),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    InMux I__975 (
            .O(N__9461),
            .I(\PCH_PWRGD.un1_count_1_cry_2 ));
    InMux I__974 (
            .O(N__9458),
            .I(N__9454));
    InMux I__973 (
            .O(N__9457),
            .I(N__9451));
    LocalMux I__972 (
            .O(N__9454),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    LocalMux I__971 (
            .O(N__9451),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    InMux I__970 (
            .O(N__9446),
            .I(\PCH_PWRGD.un1_count_1_cry_3 ));
    CascadeMux I__969 (
            .O(N__9443),
            .I(N__9440));
    InMux I__968 (
            .O(N__9440),
            .I(N__9437));
    LocalMux I__967 (
            .O(N__9437),
            .I(\POWERLED.mult1_un159_sum_cry_2_s ));
    CascadeMux I__966 (
            .O(N__9434),
            .I(N__9431));
    InMux I__965 (
            .O(N__9431),
            .I(N__9428));
    LocalMux I__964 (
            .O(N__9428),
            .I(\POWERLED.mult1_un159_sum_cry_3_s ));
    InMux I__963 (
            .O(N__9425),
            .I(N__9422));
    LocalMux I__962 (
            .O(N__9422),
            .I(\POWERLED.mult1_un159_sum_cry_4_s ));
    CascadeMux I__961 (
            .O(N__9419),
            .I(N__9415));
    InMux I__960 (
            .O(N__9418),
            .I(N__9410));
    InMux I__959 (
            .O(N__9415),
            .I(N__9403));
    InMux I__958 (
            .O(N__9414),
            .I(N__9403));
    InMux I__957 (
            .O(N__9413),
            .I(N__9403));
    LocalMux I__956 (
            .O(N__9410),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__955 (
            .O(N__9403),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    InMux I__954 (
            .O(N__9398),
            .I(N__9395));
    LocalMux I__953 (
            .O(N__9395),
            .I(\POWERLED.mult1_un159_sum_cry_5_s ));
    CascadeMux I__952 (
            .O(N__9392),
            .I(N__9388));
    CascadeMux I__951 (
            .O(N__9391),
            .I(N__9384));
    InMux I__950 (
            .O(N__9388),
            .I(N__9377));
    InMux I__949 (
            .O(N__9387),
            .I(N__9377));
    InMux I__948 (
            .O(N__9384),
            .I(N__9377));
    LocalMux I__947 (
            .O(N__9377),
            .I(G_407));
    InMux I__946 (
            .O(N__9374),
            .I(N__9371));
    LocalMux I__945 (
            .O(N__9371),
            .I(\POWERLED.mult1_un166_sum_axb_6 ));
    InMux I__944 (
            .O(N__9368),
            .I(\POWERLED.mult1_un166_sum_cry_5 ));
    InMux I__943 (
            .O(N__9365),
            .I(\POWERLED.mult1_un138_sum_cry_7 ));
    CascadeMux I__942 (
            .O(N__9362),
            .I(\POWERLED.mult1_un138_sum_s_8_cascade_ ));
    InMux I__941 (
            .O(N__9359),
            .I(\POWERLED.mult1_un159_sum_cry_1 ));
    InMux I__940 (
            .O(N__9356),
            .I(\POWERLED.mult1_un159_sum_cry_2 ));
    InMux I__939 (
            .O(N__9353),
            .I(\POWERLED.mult1_un159_sum_cry_3 ));
    InMux I__938 (
            .O(N__9350),
            .I(\POWERLED.mult1_un159_sum_cry_4 ));
    InMux I__937 (
            .O(N__9347),
            .I(\POWERLED.mult1_un159_sum_cry_5 ));
    InMux I__936 (
            .O(N__9344),
            .I(\POWERLED.mult1_un159_sum_cry_6 ));
    CascadeMux I__935 (
            .O(N__9341),
            .I(\POWERLED.mult1_un159_sum_s_7_cascade_ ));
    InMux I__934 (
            .O(N__9338),
            .I(N__9335));
    LocalMux I__933 (
            .O(N__9335),
            .I(\POWERLED.mult1_un131_sum_axb_8 ));
    InMux I__932 (
            .O(N__9332),
            .I(\POWERLED.mult1_un131_sum_cry_7 ));
    CascadeMux I__931 (
            .O(N__9329),
            .I(\POWERLED.mult1_un131_sum_s_8_cascade_ ));
    InMux I__930 (
            .O(N__9326),
            .I(\POWERLED.mult1_un138_sum_cry_2 ));
    CascadeMux I__929 (
            .O(N__9323),
            .I(N__9320));
    InMux I__928 (
            .O(N__9320),
            .I(N__9317));
    LocalMux I__927 (
            .O(N__9317),
            .I(\POWERLED.mult1_un131_sum_cry_3_s ));
    InMux I__926 (
            .O(N__9314),
            .I(\POWERLED.mult1_un138_sum_cry_3 ));
    InMux I__925 (
            .O(N__9311),
            .I(N__9308));
    LocalMux I__924 (
            .O(N__9308),
            .I(\POWERLED.mult1_un131_sum_cry_4_s ));
    InMux I__923 (
            .O(N__9305),
            .I(\POWERLED.mult1_un138_sum_cry_4 ));
    CascadeMux I__922 (
            .O(N__9302),
            .I(N__9299));
    InMux I__921 (
            .O(N__9299),
            .I(N__9296));
    LocalMux I__920 (
            .O(N__9296),
            .I(\POWERLED.mult1_un131_sum_cry_5_s ));
    InMux I__919 (
            .O(N__9293),
            .I(\POWERLED.mult1_un138_sum_cry_5 ));
    InMux I__918 (
            .O(N__9290),
            .I(N__9287));
    LocalMux I__917 (
            .O(N__9287),
            .I(\POWERLED.mult1_un131_sum_cry_6_s ));
    CascadeMux I__916 (
            .O(N__9284),
            .I(N__9280));
    CascadeMux I__915 (
            .O(N__9283),
            .I(N__9276));
    InMux I__914 (
            .O(N__9280),
            .I(N__9269));
    InMux I__913 (
            .O(N__9279),
            .I(N__9269));
    InMux I__912 (
            .O(N__9276),
            .I(N__9269));
    LocalMux I__911 (
            .O(N__9269),
            .I(\POWERLED.mult1_un131_sum_i_0_8 ));
    InMux I__910 (
            .O(N__9266),
            .I(\POWERLED.mult1_un138_sum_cry_6 ));
    InMux I__909 (
            .O(N__9263),
            .I(N__9260));
    LocalMux I__908 (
            .O(N__9260),
            .I(\POWERLED.mult1_un138_sum_axb_8 ));
    InMux I__907 (
            .O(N__9257),
            .I(\POWERLED.mult1_un124_sum_cry_6 ));
    InMux I__906 (
            .O(N__9254),
            .I(\POWERLED.mult1_un124_sum_cry_7 ));
    CascadeMux I__905 (
            .O(N__9251),
            .I(\POWERLED.mult1_un124_sum_s_8_cascade_ ));
    InMux I__904 (
            .O(N__9248),
            .I(\POWERLED.mult1_un131_sum_cry_2 ));
    CascadeMux I__903 (
            .O(N__9245),
            .I(N__9242));
    InMux I__902 (
            .O(N__9242),
            .I(N__9239));
    LocalMux I__901 (
            .O(N__9239),
            .I(\POWERLED.mult1_un124_sum_cry_3_s ));
    InMux I__900 (
            .O(N__9236),
            .I(\POWERLED.mult1_un131_sum_cry_3 ));
    InMux I__899 (
            .O(N__9233),
            .I(N__9230));
    LocalMux I__898 (
            .O(N__9230),
            .I(\POWERLED.mult1_un124_sum_cry_4_s ));
    InMux I__897 (
            .O(N__9227),
            .I(\POWERLED.mult1_un131_sum_cry_4 ));
    CascadeMux I__896 (
            .O(N__9224),
            .I(N__9221));
    InMux I__895 (
            .O(N__9221),
            .I(N__9218));
    LocalMux I__894 (
            .O(N__9218),
            .I(\POWERLED.mult1_un124_sum_cry_5_s ));
    InMux I__893 (
            .O(N__9215),
            .I(\POWERLED.mult1_un131_sum_cry_5 ));
    InMux I__892 (
            .O(N__9212),
            .I(N__9209));
    LocalMux I__891 (
            .O(N__9209),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    CascadeMux I__890 (
            .O(N__9206),
            .I(N__9202));
    CascadeMux I__889 (
            .O(N__9205),
            .I(N__9198));
    InMux I__888 (
            .O(N__9202),
            .I(N__9191));
    InMux I__887 (
            .O(N__9201),
            .I(N__9191));
    InMux I__886 (
            .O(N__9198),
            .I(N__9191));
    LocalMux I__885 (
            .O(N__9191),
            .I(\POWERLED.mult1_un124_sum_i_0_8 ));
    InMux I__884 (
            .O(N__9188),
            .I(\POWERLED.mult1_un131_sum_cry_6 ));
    CascadeMux I__883 (
            .O(N__9185),
            .I(N__9182));
    InMux I__882 (
            .O(N__9182),
            .I(N__9179));
    LocalMux I__881 (
            .O(N__9179),
            .I(\POWERLED.mult1_un103_sum_cry_5_s ));
    InMux I__880 (
            .O(N__9176),
            .I(\POWERLED.mult1_un110_sum_cry_5 ));
    InMux I__879 (
            .O(N__9173),
            .I(N__9170));
    LocalMux I__878 (
            .O(N__9170),
            .I(\POWERLED.mult1_un103_sum_cry_6_s ));
    CascadeMux I__877 (
            .O(N__9167),
            .I(N__9163));
    CascadeMux I__876 (
            .O(N__9166),
            .I(N__9159));
    InMux I__875 (
            .O(N__9163),
            .I(N__9152));
    InMux I__874 (
            .O(N__9162),
            .I(N__9152));
    InMux I__873 (
            .O(N__9159),
            .I(N__9152));
    LocalMux I__872 (
            .O(N__9152),
            .I(\POWERLED.mult1_un103_sum_i_0_8 ));
    InMux I__871 (
            .O(N__9149),
            .I(\POWERLED.mult1_un110_sum_cry_6 ));
    InMux I__870 (
            .O(N__9146),
            .I(N__9143));
    LocalMux I__869 (
            .O(N__9143),
            .I(\POWERLED.mult1_un110_sum_axb_8 ));
    InMux I__868 (
            .O(N__9140),
            .I(\POWERLED.mult1_un110_sum_cry_7 ));
    CascadeMux I__867 (
            .O(N__9137),
            .I(\POWERLED.mult1_un110_sum_s_8_cascade_ ));
    InMux I__866 (
            .O(N__9134),
            .I(\POWERLED.mult1_un124_sum_cry_2 ));
    InMux I__865 (
            .O(N__9131),
            .I(\POWERLED.mult1_un124_sum_cry_3 ));
    InMux I__864 (
            .O(N__9128),
            .I(\POWERLED.mult1_un124_sum_cry_4 ));
    InMux I__863 (
            .O(N__9125),
            .I(\POWERLED.mult1_un124_sum_cry_5 ));
    CascadeMux I__862 (
            .O(N__9122),
            .I(N__9119));
    InMux I__861 (
            .O(N__9119),
            .I(N__9116));
    LocalMux I__860 (
            .O(N__9116),
            .I(\POWERLED.mult1_un96_sum_cry_5_s ));
    InMux I__859 (
            .O(N__9113),
            .I(\POWERLED.mult1_un103_sum_cry_5 ));
    InMux I__858 (
            .O(N__9110),
            .I(N__9107));
    LocalMux I__857 (
            .O(N__9107),
            .I(\POWERLED.mult1_un96_sum_cry_6_s ));
    CascadeMux I__856 (
            .O(N__9104),
            .I(N__9100));
    CascadeMux I__855 (
            .O(N__9103),
            .I(N__9096));
    InMux I__854 (
            .O(N__9100),
            .I(N__9089));
    InMux I__853 (
            .O(N__9099),
            .I(N__9089));
    InMux I__852 (
            .O(N__9096),
            .I(N__9089));
    LocalMux I__851 (
            .O(N__9089),
            .I(\POWERLED.mult1_un96_sum_i_0_8 ));
    InMux I__850 (
            .O(N__9086),
            .I(\POWERLED.mult1_un103_sum_cry_6 ));
    InMux I__849 (
            .O(N__9083),
            .I(N__9080));
    LocalMux I__848 (
            .O(N__9080),
            .I(\POWERLED.mult1_un103_sum_axb_8 ));
    InMux I__847 (
            .O(N__9077),
            .I(\POWERLED.mult1_un103_sum_cry_7 ));
    CascadeMux I__846 (
            .O(N__9074),
            .I(\POWERLED.mult1_un103_sum_s_8_cascade_ ));
    InMux I__845 (
            .O(N__9071),
            .I(\POWERLED.mult1_un110_sum_cry_2 ));
    CascadeMux I__844 (
            .O(N__9068),
            .I(N__9065));
    InMux I__843 (
            .O(N__9065),
            .I(N__9062));
    LocalMux I__842 (
            .O(N__9062),
            .I(\POWERLED.mult1_un103_sum_cry_3_s ));
    InMux I__841 (
            .O(N__9059),
            .I(\POWERLED.mult1_un110_sum_cry_3 ));
    InMux I__840 (
            .O(N__9056),
            .I(N__9053));
    LocalMux I__839 (
            .O(N__9053),
            .I(\POWERLED.mult1_un103_sum_cry_4_s ));
    InMux I__838 (
            .O(N__9050),
            .I(\POWERLED.mult1_un110_sum_cry_4 ));
    InMux I__837 (
            .O(N__9047),
            .I(N__9044));
    LocalMux I__836 (
            .O(N__9044),
            .I(\POWERLED.mult1_un89_sum_cry_4_s ));
    InMux I__835 (
            .O(N__9041),
            .I(\POWERLED.mult1_un96_sum_cry_4 ));
    CascadeMux I__834 (
            .O(N__9038),
            .I(N__9035));
    InMux I__833 (
            .O(N__9035),
            .I(N__9032));
    LocalMux I__832 (
            .O(N__9032),
            .I(\POWERLED.mult1_un89_sum_cry_5_s ));
    InMux I__831 (
            .O(N__9029),
            .I(\POWERLED.mult1_un96_sum_cry_5 ));
    InMux I__830 (
            .O(N__9026),
            .I(N__9023));
    LocalMux I__829 (
            .O(N__9023),
            .I(\POWERLED.mult1_un89_sum_cry_6_s ));
    CascadeMux I__828 (
            .O(N__9020),
            .I(N__9016));
    CascadeMux I__827 (
            .O(N__9019),
            .I(N__9012));
    InMux I__826 (
            .O(N__9016),
            .I(N__9005));
    InMux I__825 (
            .O(N__9015),
            .I(N__9005));
    InMux I__824 (
            .O(N__9012),
            .I(N__9005));
    LocalMux I__823 (
            .O(N__9005),
            .I(\POWERLED.mult1_un89_sum_i_0_8 ));
    InMux I__822 (
            .O(N__9002),
            .I(\POWERLED.mult1_un96_sum_cry_6 ));
    InMux I__821 (
            .O(N__8999),
            .I(N__8996));
    LocalMux I__820 (
            .O(N__8996),
            .I(\POWERLED.mult1_un96_sum_axb_8 ));
    InMux I__819 (
            .O(N__8993),
            .I(\POWERLED.mult1_un96_sum_cry_7 ));
    CascadeMux I__818 (
            .O(N__8990),
            .I(\POWERLED.mult1_un96_sum_s_8_cascade_ ));
    InMux I__817 (
            .O(N__8987),
            .I(\POWERLED.mult1_un103_sum_cry_2 ));
    CascadeMux I__816 (
            .O(N__8984),
            .I(N__8981));
    InMux I__815 (
            .O(N__8981),
            .I(N__8978));
    LocalMux I__814 (
            .O(N__8978),
            .I(\POWERLED.mult1_un96_sum_cry_3_s ));
    InMux I__813 (
            .O(N__8975),
            .I(\POWERLED.mult1_un103_sum_cry_3 ));
    InMux I__812 (
            .O(N__8972),
            .I(N__8969));
    LocalMux I__811 (
            .O(N__8969),
            .I(\POWERLED.mult1_un96_sum_cry_4_s ));
    InMux I__810 (
            .O(N__8966),
            .I(\POWERLED.mult1_un103_sum_cry_4 ));
    InMux I__809 (
            .O(N__8963),
            .I(\POWERLED.mult1_un89_sum_cry_3 ));
    InMux I__808 (
            .O(N__8960),
            .I(\POWERLED.mult1_un89_sum_cry_4 ));
    InMux I__807 (
            .O(N__8957),
            .I(\POWERLED.mult1_un89_sum_cry_5 ));
    InMux I__806 (
            .O(N__8954),
            .I(\POWERLED.mult1_un89_sum_cry_6 ));
    InMux I__805 (
            .O(N__8951),
            .I(\POWERLED.mult1_un89_sum_cry_7 ));
    CascadeMux I__804 (
            .O(N__8948),
            .I(\POWERLED.mult1_un89_sum_s_8_cascade_ ));
    InMux I__803 (
            .O(N__8945),
            .I(\POWERLED.mult1_un96_sum_cry_2 ));
    CascadeMux I__802 (
            .O(N__8942),
            .I(N__8939));
    InMux I__801 (
            .O(N__8939),
            .I(N__8936));
    LocalMux I__800 (
            .O(N__8936),
            .I(\POWERLED.mult1_un89_sum_cry_3_s ));
    InMux I__799 (
            .O(N__8933),
            .I(\POWERLED.mult1_un96_sum_cry_3 ));
    CascadeMux I__798 (
            .O(N__8930),
            .I(\PCH_PWRGD.curr_state_RNI7N705Z0Z_0_cascade_ ));
    InMux I__797 (
            .O(N__8927),
            .I(N__8924));
    LocalMux I__796 (
            .O(N__8924),
            .I(\PCH_PWRGD.un4_count_8 ));
    CascadeMux I__795 (
            .O(N__8921),
            .I(\PCH_PWRGD.N_3_i_cascade_ ));
    InMux I__794 (
            .O(N__8918),
            .I(N__8912));
    InMux I__793 (
            .O(N__8917),
            .I(N__8912));
    LocalMux I__792 (
            .O(N__8912),
            .I(N__8909));
    Span4Mux_v I__791 (
            .O(N__8909),
            .I(N__8906));
    Span4Mux_v I__790 (
            .O(N__8906),
            .I(N__8903));
    Odrv4 I__789 (
            .O(N__8903),
            .I(vr_ready_vccin));
    InMux I__788 (
            .O(N__8900),
            .I(N__8887));
    InMux I__787 (
            .O(N__8899),
            .I(N__8887));
    InMux I__786 (
            .O(N__8898),
            .I(N__8887));
    InMux I__785 (
            .O(N__8897),
            .I(N__8887));
    InMux I__784 (
            .O(N__8896),
            .I(N__8884));
    LocalMux I__783 (
            .O(N__8887),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__782 (
            .O(N__8884),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    InMux I__781 (
            .O(N__8879),
            .I(N__8873));
    InMux I__780 (
            .O(N__8878),
            .I(N__8873));
    LocalMux I__779 (
            .O(N__8873),
            .I(\PCH_PWRGD.N_1_i ));
    CascadeMux I__778 (
            .O(N__8870),
            .I(N__8866));
    InMux I__777 (
            .O(N__8869),
            .I(N__8862));
    InMux I__776 (
            .O(N__8866),
            .I(N__8859));
    InMux I__775 (
            .O(N__8865),
            .I(N__8856));
    LocalMux I__774 (
            .O(N__8862),
            .I(N__8853));
    LocalMux I__773 (
            .O(N__8859),
            .I(\PCH_PWRGD.N_3_i ));
    LocalMux I__772 (
            .O(N__8856),
            .I(\PCH_PWRGD.N_3_i ));
    Odrv4 I__771 (
            .O(N__8853),
            .I(\PCH_PWRGD.N_3_i ));
    InMux I__770 (
            .O(N__8846),
            .I(N__8839));
    InMux I__769 (
            .O(N__8845),
            .I(N__8830));
    InMux I__768 (
            .O(N__8844),
            .I(N__8830));
    InMux I__767 (
            .O(N__8843),
            .I(N__8830));
    InMux I__766 (
            .O(N__8842),
            .I(N__8830));
    LocalMux I__765 (
            .O(N__8839),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__764 (
            .O(N__8830),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    InMux I__763 (
            .O(N__8825),
            .I(\POWERLED.mult1_un89_sum_cry_2 ));
    InMux I__762 (
            .O(N__8822),
            .I(N__8819));
    LocalMux I__761 (
            .O(N__8819),
            .I(\PCH_PWRGD.un4_count_11 ));
    InMux I__760 (
            .O(N__8816),
            .I(N__8813));
    LocalMux I__759 (
            .O(N__8813),
            .I(\PCH_PWRGD.un4_count_9 ));
    CascadeMux I__758 (
            .O(N__8810),
            .I(\PCH_PWRGD.un4_count_10_cascade_ ));
    CascadeMux I__757 (
            .O(N__8807),
            .I(\PCH_PWRGD.N_1_i_cascade_ ));
    CascadeMux I__756 (
            .O(N__8804),
            .I(\PCH_PWRGD.un1_curr_state_0_sqmuxa_0_cascade_ ));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(\POWERLED.dutycycle_cry_6 ),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(\POWERLED.dutycycle_cry_14 ),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_5_0_));
    defparam IN_MUX_bfv_2_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_5_0_));
    defparam IN_MUX_bfv_2_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_6_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_4_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_7_0_));
    defparam IN_MUX_bfv_4_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_5_0_));
    defparam IN_MUX_bfv_4_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_6_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_8_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(\POWERLED.un1_count_1_cry_8 ),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_5_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_16_0_ (
            .carryinitin(\POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO ),
            .carryinitout(bfn_5_16_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(\COUNTER.un4_counter_7 ),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_9_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_1_0_));
    defparam IN_MUX_bfv_9_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_2_0_ (
            .carryinitin(\COUNTER.counter_1_cry_8 ),
            .carryinitout(bfn_9_2_0_));
    defparam IN_MUX_bfv_9_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_3_0_ (
            .carryinitin(\COUNTER.counter_1_cry_16 ),
            .carryinitout(bfn_9_3_0_));
    defparam IN_MUX_bfv_9_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_4_0_ (
            .carryinitin(\COUNTER.counter_1_cry_24 ),
            .carryinitout(bfn_9_4_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_7 ),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(\POWERLED.un1_count_2_cry_7 ),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(\POWERLED.un1_count_2_cry_15 ),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_1_cry_7 ),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_1_cry_15 ),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(\POWERLED.un1_count_off_1_cry_7 ),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\POWERLED.un1_count_clk_1_cry_7 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(\POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_2_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_2_0_));
    defparam IN_MUX_bfv_2_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_3_0_ (
            .carryinitin(\PCH_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_2_3_0_));
    defparam IN_MUX_bfv_2_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_4_0_ (
            .carryinitin(\PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_2_4_0_));
    defparam IN_MUX_bfv_6_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_1_0_));
    defparam IN_MUX_bfv_6_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_2_0_ (
            .carryinitin(\HDA_STRAP.un1_count_1_cry_7 ),
            .carryinitout(bfn_6_2_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(\HDA_STRAP.un1_count_1_cry_15 ),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(\ALL_SYS_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(\ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_8_7_0_));
    ICE_GB \COUNTER.tmp_RNIRH3P_0  (
            .USERSIGNALTOGLOBALBUFFER(N__17737),
            .GLOBALBUFFEROUTPUT(N_65_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIESHJ_1_LC_1_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIESHJ_1_LC_1_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIESHJ_1_LC_1_2_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \PCH_PWRGD.count_RNIESHJ_1_LC_1_2_0  (
            .in0(N__9694),
            .in1(N__9487),
            .in2(N__9632),
            .in3(N__9502),
            .lcout(\PCH_PWRGD.un4_count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI7J2B_3_LC_1_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI7J2B_3_LC_1_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI7J2B_3_LC_1_2_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNI7J2B_3_LC_1_2_2  (
            .in0(N__9709),
            .in1(N__9457),
            .in2(N__9680),
            .in3(N__9472),
            .lcout(\PCH_PWRGD.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIN5IJ_0_LC_1_3_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIN5IJ_0_LC_1_3_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIN5IJ_0_LC_1_3_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PCH_PWRGD.count_RNIN5IJ_0_LC_1_3_1  (
            .in0(N__9646),
            .in1(N__9514),
            .in2(N__9614),
            .in3(N__9661),
            .lcout(),
            .ltout(\PCH_PWRGD.un4_count_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_1_3_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_1_3_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_1_3_2  (
            .in0(N__8822),
            .in1(N__8816),
            .in2(N__8810),
            .in3(N__8927),
            .lcout(\PCH_PWRGD.N_1_i ),
            .ltout(\PCH_PWRGD.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIC5474_0_LC_1_3_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIC5474_0_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIC5474_0_LC_1_3_3 .LUT_INIT=16'b1100111011011111;
    LogicCell40 \PCH_PWRGD.curr_state_RNIC5474_0_LC_1_3_3  (
            .in0(N__8846),
            .in1(N__8896),
            .in2(N__8807),
            .in3(N__8869),
            .lcout(),
            .ltout(\PCH_PWRGD.un1_curr_state_0_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI7N705_0_LC_1_3_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI7N705_0_LC_1_3_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI7N705_0_LC_1_3_4 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI7N705_0_LC_1_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8804),
            .in3(N__20059),
            .lcout(\PCH_PWRGD.curr_state_RNI7N705Z0Z_0 ),
            .ltout(\PCH_PWRGD.curr_state_RNI7N705Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_esr_RNO_0_15_LC_1_3_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_esr_RNO_0_15_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_esr_RNO_0_15_LC_1_3_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \PCH_PWRGD.count_esr_RNO_0_15_LC_1_3_5  (
            .in0(N__20060),
            .in1(_gnd_net_),
            .in2(N__8930),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.N_65_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_esr_RNIFR521_15_LC_1_3_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_esr_RNIFR521_15_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_esr_RNIFR521_15_LC_1_3_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \PCH_PWRGD.count_esr_RNIFR521_15_LC_1_3_7  (
            .in0(N__9814),
            .in1(N__9829),
            .in2(N__9797),
            .in3(N__9595),
            .lcout(\PCH_PWRGD.un4_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_sys_pwrok_LC_1_4_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_sys_pwrok_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_sys_pwrok_LC_1_4_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \PCH_PWRGD.un2_sys_pwrok_LC_1_4_0  (
            .in0(N__19283),
            .in1(N__8918),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.N_3_i ),
            .ltout(\PCH_PWRGD.N_3_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_0_LC_1_4_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_0_LC_1_4_1 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_0_LC_1_4_1 .LUT_INIT=16'b0100010010100000;
    LogicCell40 \PCH_PWRGD.curr_state_0_LC_1_4_1  (
            .in0(N__8898),
            .in1(N__8878),
            .in2(N__8921),
            .in3(N__8845),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20560),
            .ce(N__19787),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.pch_pwrok_LC_1_4_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.pch_pwrok_LC_1_4_5 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.pch_pwrok_LC_1_4_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \PCH_PWRGD.pch_pwrok_LC_1_4_5  (
            .in0(N__8900),
            .in1(N__8844),
            .in2(_gnd_net_),
            .in3(N__8865),
            .lcout(pch_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20560),
            .ce(N__19787),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIHKNI1_0_LC_1_4_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIHKNI1_0_LC_1_4_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIHKNI1_0_LC_1_4_6 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \PCH_PWRGD.curr_state_RNIHKNI1_0_LC_1_4_6  (
            .in0(N__8842),
            .in1(N__8897),
            .in2(N__19286),
            .in3(N__8917),
            .lcout(\PCH_PWRGD.un1_curr_state10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_1_LC_1_4_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_1_LC_1_4_7 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_1_LC_1_4_7 .LUT_INIT=16'b0001000101010000;
    LogicCell40 \PCH_PWRGD.curr_state_1_LC_1_4_7  (
            .in0(N__8899),
            .in1(N__8879),
            .in2(N__8870),
            .in3(N__8843),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20560),
            .ce(N__19787),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_1_5_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_1_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(N__12848),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_5_0_),
            .carryout(\POWERLED.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_1_5_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_1_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_1_5_1  (
            .in0(_gnd_net_),
            .in1(N__11663),
            .in2(N__9889),
            .in3(N__8825),
            .lcout(\POWERLED.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_1_5_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_1_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_1_5_2  (
            .in0(_gnd_net_),
            .in1(N__9885),
            .in2(N__9752),
            .in3(N__8963),
            .lcout(\POWERLED.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_1_5_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_1_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_1_5_3  (
            .in0(_gnd_net_),
            .in1(N__9740),
            .in2(N__10102),
            .in3(N__8960),
            .lcout(\POWERLED.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_1_5_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_1_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_1_5_4  (
            .in0(_gnd_net_),
            .in1(N__10098),
            .in2(N__9731),
            .in3(N__8957),
            .lcout(\POWERLED.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_1_5_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_1_5_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_1_5_5  (
            .in0(N__10121),
            .in1(N__9719),
            .in2(N__9890),
            .in3(N__8954),
            .lcout(\POWERLED.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_1_5_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_1_5_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_1_5_6  (
            .in0(_gnd_net_),
            .in1(N__9905),
            .in2(_gnd_net_),
            .in3(N__8951),
            .lcout(\POWERLED.mult1_un89_sum_s_8 ),
            .ltout(\POWERLED.mult1_un89_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_5_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_5_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8948),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_1_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_1_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__12874),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(\POWERLED.mult1_un96_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_1_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_1_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__10295),
            .in2(N__9019),
            .in3(N__8945),
            .lcout(\POWERLED.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_1_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_1_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(N__9015),
            .in2(N__8942),
            .in3(N__8933),
            .lcout(\POWERLED.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_1_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_1_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(N__9047),
            .in2(N__10129),
            .in3(N__9041),
            .lcout(\POWERLED.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_1_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_1_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(N__10125),
            .in2(N__9038),
            .in3(N__9029),
            .lcout(\POWERLED.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_1_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_1_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_1_6_5  (
            .in0(N__9560),
            .in1(N__9026),
            .in2(N__9020),
            .in3(N__9002),
            .lcout(\POWERLED.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_1_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_1_6_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(N__8999),
            .in2(_gnd_net_),
            .in3(N__8993),
            .lcout(\POWERLED.mult1_un96_sum_s_8 ),
            .ltout(\POWERLED.mult1_un96_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_6_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_6_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8990),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__12916),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(\POWERLED.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(N__9581),
            .in2(N__9103),
            .in3(N__8987),
            .lcout(\POWERLED.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_7_2  (
            .in0(_gnd_net_),
            .in1(N__9099),
            .in2(N__8984),
            .in3(N__8975),
            .lcout(\POWERLED.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_7_3  (
            .in0(_gnd_net_),
            .in1(N__8972),
            .in2(N__9568),
            .in3(N__8966),
            .lcout(\POWERLED.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_7_4  (
            .in0(_gnd_net_),
            .in1(N__9564),
            .in2(N__9122),
            .in3(N__9113),
            .lcout(\POWERLED.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_7_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_7_5  (
            .in0(N__10007),
            .in1(N__9110),
            .in2(N__9104),
            .in3(N__9086),
            .lcout(\POWERLED.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_7_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_7_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_7_6  (
            .in0(_gnd_net_),
            .in1(N__9083),
            .in2(_gnd_net_),
            .in3(N__9077),
            .lcout(\POWERLED.mult1_un103_sum_s_8 ),
            .ltout(\POWERLED.mult1_un103_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_7_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9074),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(N__12950),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_8_0_),
            .carryout(\POWERLED.mult1_un110_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_8_1  (
            .in0(_gnd_net_),
            .in1(N__10019),
            .in2(N__9166),
            .in3(N__9071),
            .lcout(\POWERLED.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(N__9162),
            .in2(N__9068),
            .in3(N__9059),
            .lcout(\POWERLED.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_8_3  (
            .in0(_gnd_net_),
            .in1(N__9056),
            .in2(N__10013),
            .in3(N__9050),
            .lcout(\POWERLED.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(N__10011),
            .in2(N__9185),
            .in3(N__9176),
            .lcout(\POWERLED.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_8_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_8_5  (
            .in0(N__10229),
            .in1(N__9173),
            .in2(N__9167),
            .in3(N__9149),
            .lcout(\POWERLED.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_8_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_8_6  (
            .in0(_gnd_net_),
            .in1(N__9146),
            .in2(_gnd_net_),
            .in3(N__9140),
            .lcout(\POWERLED.mult1_un110_sum_s_8 ),
            .ltout(\POWERLED.mult1_un110_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_1_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_1_8_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_1_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9137),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_1_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_1_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(N__13007),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\POWERLED.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_1_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_1_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(N__11369),
            .in2(N__10396),
            .in3(N__9134),
            .lcout(\POWERLED.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_1_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_1_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__10392),
            .in2(N__10283),
            .in3(N__9131),
            .lcout(\POWERLED.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_1_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_1_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(N__10262),
            .in2(N__10321),
            .in3(N__9128),
            .lcout(\POWERLED.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_1_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_1_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(N__10317),
            .in2(N__10247),
            .in3(N__9125),
            .lcout(\POWERLED.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_1_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_1_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_1_9_5  (
            .in0(N__10373),
            .in1(N__10202),
            .in2(N__10397),
            .in3(N__9257),
            .lcout(\POWERLED.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_1_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_1_9_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_1_9_6  (
            .in0(_gnd_net_),
            .in1(N__10169),
            .in2(_gnd_net_),
            .in3(N__9254),
            .lcout(\POWERLED.mult1_un124_sum_s_8 ),
            .ltout(\POWERLED.mult1_un124_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_9_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9251),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__12682),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\POWERLED.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__11381),
            .in2(N__9205),
            .in3(N__9248),
            .lcout(\POWERLED.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__9201),
            .in2(N__9245),
            .in3(N__9236),
            .lcout(\POWERLED.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__9233),
            .in2(N__10379),
            .in3(N__9227),
            .lcout(\POWERLED.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__10377),
            .in2(N__9224),
            .in3(N__9215),
            .lcout(\POWERLED.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_10_5  (
            .in0(N__10349),
            .in1(N__9212),
            .in2(N__9206),
            .in3(N__9188),
            .lcout(\POWERLED.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_10_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(N__9338),
            .in2(_gnd_net_),
            .in3(N__9332),
            .lcout(\POWERLED.mult1_un131_sum_s_8 ),
            .ltout(\POWERLED.mult1_un131_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_10_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9329),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__12730),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\POWERLED.mult1_un138_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__10331),
            .in2(N__9283),
            .in3(N__9326),
            .lcout(\POWERLED.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__9279),
            .in2(N__9323),
            .in3(N__9314),
            .lcout(\POWERLED.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__9311),
            .in2(N__10355),
            .in3(N__9305),
            .lcout(\POWERLED.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__10353),
            .in2(N__9302),
            .in3(N__9293),
            .lcout(\POWERLED.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_11_5  (
            .in0(N__11326),
            .in1(N__9290),
            .in2(N__9284),
            .in3(N__9266),
            .lcout(\POWERLED.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__9263),
            .in2(_gnd_net_),
            .in3(N__9365),
            .lcout(\POWERLED.mult1_un138_sum_s_8 ),
            .ltout(\POWERLED.mult1_un138_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9362),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_1_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_1_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__14129),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\POWERLED.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_1_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_1_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__11540),
            .in2(N__10516),
            .in3(N__9359),
            .lcout(\POWERLED.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_1_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_1_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__10512),
            .in2(N__10676),
            .in3(N__9356),
            .lcout(\POWERLED.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_1_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_1_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__10655),
            .in2(N__10544),
            .in3(N__9353),
            .lcout(\POWERLED.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_1_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_1_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(N__10542),
            .in2(N__10640),
            .in3(N__9350),
            .lcout(\POWERLED.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_1_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_1_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_1_12_5  (
            .in0(N__9418),
            .in1(N__10595),
            .in2(N__10517),
            .in3(N__9347),
            .lcout(\POWERLED.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_1_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_1_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__10562),
            .in2(_gnd_net_),
            .in3(N__9344),
            .lcout(\POWERLED.mult1_un159_sum_s_7 ),
            .ltout(\POWERLED.mult1_un159_sum_s_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_1_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_1_12_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9341),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_1_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_1_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__14209),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\POWERLED.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_1_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_1_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__11552),
            .in2(N__9391),
            .in3(N__9413),
            .lcout(G_407),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_0 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_1_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_1_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__9387),
            .in2(N__9443),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_1_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_1_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__9414),
            .in2(N__9434),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_1_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_1_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__9425),
            .in2(N__9419),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_1_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_1_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__9398),
            .in2(N__9392),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_1_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_1_13_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__9374),
            .in2(_gnd_net_),
            .in3(N__9368),
            .lcout(\POWERLED.un1_count_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_1_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_1_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_1_13_7  (
            .in0(N__10543),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_1_14_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_1_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12878),
            .lcout(\POWERLED.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_1_14_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_1_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9572),
            .lcout(\POWERLED.un1_count_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_LC_1_14_6 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_LC_1_14_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.pwm_out_LC_1_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.pwm_out_LC_1_14_6  (
            .in0(N__11602),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwrbtn_led),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20628),
            .ce(N__11087),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_0_LC_1_15_6 .C_ON=1'b0;
    defparam \POWERLED.curr_state_0_LC_1_15_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.curr_state_0_LC_1_15_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \POWERLED.curr_state_0_LC_1_15_6  (
            .in0(N__11601),
            .in1(N__11612),
            .in2(_gnd_net_),
            .in3(N__10823),
            .lcout(\POWERLED.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20629),
            .ce(N__19812),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_0_LC_2_2_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_0_LC_2_2_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_0_LC_2_2_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_0_LC_2_2_0  (
            .in0(N__20074),
            .in1(N__9515),
            .in2(N__9533),
            .in3(N__9532),
            .lcout(\PCH_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_2_2_0_),
            .carryout(\PCH_PWRGD.un1_count_1_cry_0 ),
            .clk(N__20466),
            .ce(),
            .sr(N__9769));
    defparam \PCH_PWRGD.count_1_LC_2_2_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_1_LC_2_2_1 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_1_LC_2_2_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_1_LC_2_2_1  (
            .in0(N__20067),
            .in1(N__9503),
            .in2(_gnd_net_),
            .in3(N__9491),
            .lcout(\PCH_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_0 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_1 ),
            .clk(N__20466),
            .ce(),
            .sr(N__9769));
    defparam \PCH_PWRGD.count_2_LC_2_2_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_2_LC_2_2_2 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_2_LC_2_2_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_2_LC_2_2_2  (
            .in0(N__20075),
            .in1(N__9488),
            .in2(_gnd_net_),
            .in3(N__9476),
            .lcout(\PCH_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_1 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_2 ),
            .clk(N__20466),
            .ce(),
            .sr(N__9769));
    defparam \PCH_PWRGD.count_3_LC_2_2_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_3_LC_2_2_3 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_3_LC_2_2_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_3_LC_2_2_3  (
            .in0(N__20068),
            .in1(N__9473),
            .in2(_gnd_net_),
            .in3(N__9461),
            .lcout(\PCH_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_2 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_3 ),
            .clk(N__20466),
            .ce(),
            .sr(N__9769));
    defparam \PCH_PWRGD.count_4_LC_2_2_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_4_LC_2_2_4 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_4_LC_2_2_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_4_LC_2_2_4  (
            .in0(N__20076),
            .in1(N__9458),
            .in2(_gnd_net_),
            .in3(N__9446),
            .lcout(\PCH_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_3 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_4 ),
            .clk(N__20466),
            .ce(),
            .sr(N__9769));
    defparam \PCH_PWRGD.count_5_LC_2_2_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_5_LC_2_2_5 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_5_LC_2_2_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_5_LC_2_2_5  (
            .in0(N__20069),
            .in1(N__9710),
            .in2(_gnd_net_),
            .in3(N__9698),
            .lcout(\PCH_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_4 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_5 ),
            .clk(N__20466),
            .ce(),
            .sr(N__9769));
    defparam \PCH_PWRGD.count_6_LC_2_2_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_6_LC_2_2_6 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_6_LC_2_2_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_6_LC_2_2_6  (
            .in0(N__20077),
            .in1(N__9695),
            .in2(_gnd_net_),
            .in3(N__9683),
            .lcout(\PCH_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_5 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_6 ),
            .clk(N__20466),
            .ce(),
            .sr(N__9769));
    defparam \PCH_PWRGD.count_7_LC_2_2_7 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_7_LC_2_2_7 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_7_LC_2_2_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_7_LC_2_2_7  (
            .in0(N__20070),
            .in1(N__9679),
            .in2(_gnd_net_),
            .in3(N__9665),
            .lcout(\PCH_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_6 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_7 ),
            .clk(N__20466),
            .ce(),
            .sr(N__9769));
    defparam \PCH_PWRGD.count_8_LC_2_3_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_8_LC_2_3_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_8_LC_2_3_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_8_LC_2_3_0  (
            .in0(N__20117),
            .in1(N__9662),
            .in2(_gnd_net_),
            .in3(N__9650),
            .lcout(\PCH_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_2_3_0_),
            .carryout(\PCH_PWRGD.un1_count_1_cry_8 ),
            .clk(N__20532),
            .ce(),
            .sr(N__9768));
    defparam \PCH_PWRGD.count_9_LC_2_3_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_9_LC_2_3_1 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_9_LC_2_3_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_9_LC_2_3_1  (
            .in0(N__20102),
            .in1(N__9647),
            .in2(_gnd_net_),
            .in3(N__9635),
            .lcout(\PCH_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_8 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_9 ),
            .clk(N__20532),
            .ce(),
            .sr(N__9768));
    defparam \PCH_PWRGD.count_10_LC_2_3_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_10_LC_2_3_2 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_10_LC_2_3_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_10_LC_2_3_2  (
            .in0(N__20114),
            .in1(N__9631),
            .in2(_gnd_net_),
            .in3(N__9617),
            .lcout(\PCH_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_9 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_10 ),
            .clk(N__20532),
            .ce(),
            .sr(N__9768));
    defparam \PCH_PWRGD.count_11_LC_2_3_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_11_LC_2_3_3 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_11_LC_2_3_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_11_LC_2_3_3  (
            .in0(N__20100),
            .in1(N__9613),
            .in2(_gnd_net_),
            .in3(N__9599),
            .lcout(\PCH_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_10 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_11 ),
            .clk(N__20532),
            .ce(),
            .sr(N__9768));
    defparam \PCH_PWRGD.count_12_LC_2_3_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_12_LC_2_3_4 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_12_LC_2_3_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_12_LC_2_3_4  (
            .in0(N__20115),
            .in1(N__9596),
            .in2(_gnd_net_),
            .in3(N__9584),
            .lcout(\PCH_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_11 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_12 ),
            .clk(N__20532),
            .ce(),
            .sr(N__9768));
    defparam \PCH_PWRGD.count_13_LC_2_3_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_13_LC_2_3_5 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_13_LC_2_3_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_13_LC_2_3_5  (
            .in0(N__20101),
            .in1(N__9830),
            .in2(_gnd_net_),
            .in3(N__9818),
            .lcout(\PCH_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_12 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_13 ),
            .clk(N__20532),
            .ce(),
            .sr(N__9768));
    defparam \PCH_PWRGD.count_14_LC_2_3_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_14_LC_2_3_6 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_14_LC_2_3_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_14_LC_2_3_6  (
            .in0(N__20116),
            .in1(N__9815),
            .in2(_gnd_net_),
            .in3(N__9803),
            .lcout(\PCH_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_13 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_14 ),
            .clk(N__20532),
            .ce(),
            .sr(N__9768));
    defparam \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_3_7 .C_ON=1'b1;
    defparam \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_3_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_3_7  (
            .in0(_gnd_net_),
            .in1(N__18395),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_14 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_esr_15_LC_2_4_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_esr_15_LC_2_4_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_esr_15_LC_2_4_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \PCH_PWRGD.count_esr_15_LC_2_4_0  (
            .in0(_gnd_net_),
            .in1(N__9796),
            .in2(_gnd_net_),
            .in3(N__9800),
            .lcout(\PCH_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20542),
            .ce(N__9782),
            .sr(N__9770));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_2_5_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_2_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_2_5_0  (
            .in0(_gnd_net_),
            .in1(N__12818),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_5_0_),
            .carryout(\POWERLED.mult1_un82_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_2_5_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_2_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_2_5_1  (
            .in0(_gnd_net_),
            .in1(N__11753),
            .in2(N__9973),
            .in3(N__9743),
            .lcout(\POWERLED.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_2_5_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_2_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_2_5_2  (
            .in0(_gnd_net_),
            .in1(N__9969),
            .in2(N__9872),
            .in3(N__9734),
            .lcout(\POWERLED.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_2_5_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_2_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_2_5_3  (
            .in0(_gnd_net_),
            .in1(N__9860),
            .in2(N__10045),
            .in3(N__9722),
            .lcout(\POWERLED.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_2_5_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_2_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_2_5_4  (
            .in0(_gnd_net_),
            .in1(N__10041),
            .in2(N__9851),
            .in3(N__9713),
            .lcout(\POWERLED.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_2_5_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_2_5_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_2_5_5  (
            .in0(N__10094),
            .in1(N__9839),
            .in2(N__9974),
            .in3(N__9899),
            .lcout(\POWERLED.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_2_5_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_2_5_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_2_5_6  (
            .in0(_gnd_net_),
            .in1(N__9989),
            .in2(_gnd_net_),
            .in3(N__9896),
            .lcout(\POWERLED.mult1_un82_sum_s_8 ),
            .ltout(\POWERLED.mult1_un82_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_2_5_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_2_5_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_2_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9893),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(N__12794),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_6_0_),
            .carryout(\POWERLED.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_2_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_2_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(N__11285),
            .in2(N__10147),
            .in3(N__9863),
            .lcout(\POWERLED.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_2_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_2_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_2_6_2  (
            .in0(_gnd_net_),
            .in1(N__10143),
            .in2(N__9956),
            .in3(N__9854),
            .lcout(\POWERLED.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_2_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_2_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_2_6_3  (
            .in0(_gnd_net_),
            .in1(N__9944),
            .in2(N__10076),
            .in3(N__9842),
            .lcout(\POWERLED.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_2_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_2_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_2_6_4  (
            .in0(_gnd_net_),
            .in1(N__10074),
            .in2(N__9935),
            .in3(N__9833),
            .lcout(\POWERLED.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_2_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_2_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_2_6_5  (
            .in0(N__10037),
            .in1(N__9923),
            .in2(N__10148),
            .in3(N__9983),
            .lcout(\POWERLED.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_2_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_2_6_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_2_6_6  (
            .in0(_gnd_net_),
            .in1(N__9914),
            .in2(_gnd_net_),
            .in3(N__9980),
            .lcout(\POWERLED.mult1_un75_sum_s_8 ),
            .ltout(\POWERLED.mult1_un75_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_2_6_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_2_6_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_2_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9977),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_2_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_2_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_2_7_0  (
            .in0(_gnd_net_),
            .in1(N__13184),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_7_0_),
            .carryout(\POWERLED.mult1_un68_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_2_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_2_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(N__11768),
            .in2(N__11428),
            .in3(N__9947),
            .lcout(\POWERLED.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_2_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_2_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(N__11424),
            .in2(N__11276),
            .in3(N__9938),
            .lcout(\POWERLED.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_2_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_2_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_2_7_3  (
            .in0(_gnd_net_),
            .in1(N__11246),
            .in2(N__11464),
            .in3(N__9926),
            .lcout(\POWERLED.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_2_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_2_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_2_7_4  (
            .in0(_gnd_net_),
            .in1(N__11460),
            .in2(N__11225),
            .in3(N__9917),
            .lcout(\POWERLED.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_2_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_2_7_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_2_7_5  (
            .in0(N__10070),
            .in1(N__11198),
            .in2(N__11429),
            .in3(N__9908),
            .lcout(\POWERLED.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_2_7_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_2_7_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_2_7_6  (
            .in0(_gnd_net_),
            .in1(N__11159),
            .in2(_gnd_net_),
            .in3(N__10151),
            .lcout(\POWERLED.mult1_un68_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_2_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_2_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_2_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10069),
            .lcout(\POWERLED.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_2_8_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_2_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10234),
            .lcout(\POWERLED.un1_count_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_8_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_8_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_8_1  (
            .in0(_gnd_net_),
            .in1(N__10130),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_8_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_8_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(N__10103),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_2_8_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_2_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_2_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10075),
            .lcout(\POWERLED.un1_count_2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_8_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10046),
            .lcout(\POWERLED.un1_count_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_2_8_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_2_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12917),
            .lcout(\POWERLED.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_2_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_2_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10012),
            .lcout(\POWERLED.un1_count_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12847),
            .lcout(\POWERLED.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(N__12979),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(\POWERLED.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(N__11408),
            .in2(N__10186),
            .in3(N__10274),
            .lcout(\POWERLED.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(N__10182),
            .in2(N__10271),
            .in3(N__10256),
            .lcout(\POWERLED.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__10253),
            .in2(N__10235),
            .in3(N__10238),
            .lcout(\POWERLED.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__10233),
            .in2(N__10211),
            .in3(N__10196),
            .lcout(\POWERLED.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_9_5  (
            .in0(N__10313),
            .in1(N__10193),
            .in2(N__10187),
            .in3(N__10163),
            .lcout(\POWERLED.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_9_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__10160),
            .in2(_gnd_net_),
            .in3(N__10154),
            .lcout(\POWERLED.mult1_un117_sum_s_8 ),
            .ltout(\POWERLED.mult1_un117_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_2_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_2_9_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10400),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_2_10_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_2_10_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_2_10_0  (
            .in0(N__10378),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_10_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_10_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_10_1  (
            .in0(N__10354),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_4_l_fx_LC_2_10_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_4_l_fx_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_4_l_fx_LC_2_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_4_l_fx_LC_2_10_2  (
            .in0(N__10472),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11325),
            .lcout(\POWERLED.mult1_un145_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_2_10_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_2_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10627),
            .lcout(\POWERLED.un1_count_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_10_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12683),
            .lcout(\POWERLED.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_2_10_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_2_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_2_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12758),
            .lcout(\POWERLED.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10322),
            .lcout(\POWERLED.un1_count_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_2_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_2_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11465),
            .lcout(\POWERLED.un1_count_2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_2_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_2_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__12757),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\POWERLED.mult1_un145_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_2_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_2_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__11396),
            .in2(N__10484),
            .in3(N__10475),
            .lcout(\POWERLED.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_2_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_2_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__10471),
            .in2(N__10460),
            .in3(N__10451),
            .lcout(\POWERLED.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_2_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_2_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__10448),
            .in2(N__11333),
            .in3(N__10439),
            .lcout(\POWERLED.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_2_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_2_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__11330),
            .in2(N__10436),
            .in3(N__10427),
            .lcout(\POWERLED.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_2_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_2_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_2_11_5  (
            .in0(N__10622),
            .in1(N__11356),
            .in2(N__11345),
            .in3(N__10424),
            .lcout(\POWERLED.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_2_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_2_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__10421),
            .in2(_gnd_net_),
            .in3(N__10415),
            .lcout(\POWERLED.mult1_un145_sum_s_8 ),
            .ltout(\POWERLED.mult1_un145_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_2_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_2_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10412),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_2_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_2_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__14752),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\POWERLED.mult1_un152_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_2_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_2_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__10409),
            .in2(N__10579),
            .in3(N__10667),
            .lcout(\POWERLED.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_2_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_2_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__10575),
            .in2(N__10664),
            .in3(N__10649),
            .lcout(\POWERLED.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_2_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_2_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__10646),
            .in2(N__10628),
            .in3(N__10631),
            .lcout(\POWERLED.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_2_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_2_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__10626),
            .in2(N__10604),
            .in3(N__10589),
            .lcout(\POWERLED.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_2_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_2_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_2_12_5  (
            .in0(N__10538),
            .in1(N__10586),
            .in2(N__10580),
            .in3(N__10556),
            .lcout(\POWERLED.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_2_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_2_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(N__10553),
            .in2(_gnd_net_),
            .in3(N__10547),
            .lcout(\POWERLED.mult1_un152_sum_s_8 ),
            .ltout(\POWERLED.mult1_un152_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_2_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_2_12_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10520),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_0_c_inv_LC_2_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_0_c_inv_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_0_c_inv_LC_2_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_0_c_inv_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__10490),
            .in2(N__10499),
            .in3(N__12041),
            .lcout(\POWERLED.count_i_0_0 ),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\POWERLED.un1_count_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_1_c_inv_LC_2_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_1_c_inv_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_1_c_inv_LC_2_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_1_c_inv_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__10808),
            .in2(N__10817),
            .in3(N__12017),
            .lcout(\POWERLED.count_i_1 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_0 ),
            .carryout(\POWERLED.un1_count_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_2_c_inv_LC_2_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_2_c_inv_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_2_c_inv_LC_2_13_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_count_2_cry_2_c_inv_LC_2_13_2  (
            .in0(N__11990),
            .in1(N__10799),
            .in2(N__10793),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_i_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_1 ),
            .carryout(\POWERLED.un1_count_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_3_c_inv_LC_2_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_3_c_inv_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_3_c_inv_LC_2_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_3_c_inv_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__10784),
            .in2(N__10775),
            .in3(N__11960),
            .lcout(\POWERLED.count_i_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_2 ),
            .carryout(\POWERLED.un1_count_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_4_c_inv_LC_2_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_4_c_inv_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_4_c_inv_LC_2_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_4_c_inv_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__11297),
            .in2(N__10766),
            .in3(N__12476),
            .lcout(\POWERLED.count_i_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_3 ),
            .carryout(\POWERLED.un1_count_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_5_c_inv_LC_2_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_5_c_inv_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_5_c_inv_LC_2_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_5_c_inv_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__10754),
            .in2(N__10745),
            .in3(N__12446),
            .lcout(\POWERLED.count_i_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_4 ),
            .carryout(\POWERLED.un1_count_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_6_c_inv_LC_2_13_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_6_c_inv_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_6_c_inv_LC_2_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_6_c_inv_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(N__10736),
            .in2(N__10727),
            .in3(N__12416),
            .lcout(\POWERLED.count_i_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_5 ),
            .carryout(\POWERLED.un1_count_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_7_c_inv_LC_2_13_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_7_c_inv_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_7_c_inv_LC_2_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_7_c_inv_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__10715),
            .in2(N__10706),
            .in3(N__12385),
            .lcout(\POWERLED.count_i_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_6 ),
            .carryout(\POWERLED.un1_count_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_8_c_inv_LC_2_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_8_c_inv_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_8_c_inv_LC_2_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_8_c_inv_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__10694),
            .in2(N__10685),
            .in3(N__12353),
            .lcout(\POWERLED.count_i_8 ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\POWERLED.un1_count_2_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_9_c_inv_LC_2_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_9_c_inv_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_9_c_inv_LC_2_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_9_c_inv_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__10967),
            .in2(N__10958),
            .in3(N__12326),
            .lcout(\POWERLED.count_i_9 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_8 ),
            .carryout(\POWERLED.un1_count_2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_10_c_inv_LC_2_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_10_c_inv_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_10_c_inv_LC_2_14_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_count_2_cry_10_c_inv_LC_2_14_2  (
            .in0(N__12290),
            .in1(N__10949),
            .in2(N__10943),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_i_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_9 ),
            .carryout(\POWERLED.un1_count_2_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_11_c_inv_LC_2_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_11_c_inv_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_11_c_inv_LC_2_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_11_c_inv_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__10934),
            .in2(N__10925),
            .in3(N__12260),
            .lcout(\POWERLED.count_i_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_10 ),
            .carryout(\POWERLED.un1_count_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_12_c_inv_LC_2_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_12_c_inv_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_12_c_inv_LC_2_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_12_c_inv_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__10916),
            .in2(N__10904),
            .in3(N__12227),
            .lcout(\POWERLED.count_i_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_11 ),
            .carryout(\POWERLED.un1_count_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_13_c_inv_LC_2_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_13_c_inv_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_13_c_inv_LC_2_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_13_c_inv_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__10892),
            .in2(N__10880),
            .in3(N__12626),
            .lcout(\POWERLED.count_i_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_12 ),
            .carryout(\POWERLED.un1_count_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_14_c_inv_LC_2_14_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_14_c_inv_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_14_c_inv_LC_2_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_14_c_inv_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__10871),
            .in2(N__10859),
            .in3(N__12596),
            .lcout(\POWERLED.count_i_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_13 ),
            .carryout(\POWERLED.un1_count_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_15_c_inv_LC_2_14_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_15_c_inv_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_15_c_inv_LC_2_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_15_c_inv_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__10847),
            .in2(N__10835),
            .in3(N__12560),
            .lcout(\POWERLED.count_i_15 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_14 ),
            .carryout(\POWERLED.un1_count_2_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_2_15_0 .C_ON=1'b0;
    defparam \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_2_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10826),
            .lcout(\POWERLED.un1_count_2_cry_15_THRU_CO ),
            .ltout(\POWERLED.un1_count_2_cry_15_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_LC_2_15_1 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_LC_2_15_1 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \POWERLED.pwm_out_RNO_LC_2_15_1  (
            .in0(N__11600),
            .in1(N__11525),
            .in2(N__11090),
            .in3(N__17738),
            .lcout(\POWERLED.pwm_out_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_vddq_en_LC_2_15_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_vddq_en_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_vddq_en_LC_2_15_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \VPP_VDDQ.un1_vddq_en_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(N__11075),
            .in2(_gnd_net_),
            .in3(N__15659),
            .lcout(vddq_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNI1S0J_0_LC_4_2_4 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNI1S0J_0_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNI1S0J_0_LC_4_2_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \HDA_STRAP.curr_state_RNI1S0J_0_LC_4_2_4  (
            .in0(_gnd_net_),
            .in1(N__11021),
            .in2(_gnd_net_),
            .in3(N__15777),
            .lcout(\HDA_STRAP.N_5_0 ),
            .ltout(\HDA_STRAP.N_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_4_2_5 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_4_2_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_4_2_5 .LUT_INIT=16'b0000101101010101;
    LogicCell40 \HDA_STRAP.curr_state_RNO_0_0_LC_4_2_5  (
            .in0(N__15778),
            .in1(N__11051),
            .in2(N__11036),
            .in3(N__15867),
            .lcout(\HDA_STRAP.m14_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_0_LC_4_3_7 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_0_LC_4_3_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_0_LC_4_3_7 .LUT_INIT=16'b1111000010100011;
    LogicCell40 \HDA_STRAP.curr_state_0_LC_4_3_7  (
            .in0(N__11029),
            .in1(N__15735),
            .in2(N__10985),
            .in3(N__15914),
            .lcout(\HDA_STRAP.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20428),
            .ce(N__19740),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_5_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_5_0  (
            .in0(_gnd_net_),
            .in1(N__13139),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_5_0_),
            .carryout(\POWERLED.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_5_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_5_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11654),
            .in3(N__10976),
            .lcout(\POWERLED.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_5_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_5_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11138),
            .in3(N__10973),
            .lcout(\POWERLED.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_5_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(N__18387),
            .in2(N__11126),
            .in3(N__10970),
            .lcout(\POWERLED.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_5_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(N__18388),
            .in2(N__11114),
            .in3(N__11147),
            .lcout(\POWERLED.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_4_5_5 .C_ON=1'b1;
    defparam \POWERLED.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_4_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_4_5_5  (
            .in0(_gnd_net_),
            .in1(N__11512),
            .in2(_gnd_net_),
            .in3(N__11144),
            .lcout(\POWERLED.mult1_un54_sum_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_4_5_6 .C_ON=1'b0;
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_4_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_4_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11141),
            .lcout(\POWERLED.mult1_un54_sum_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13118),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_6_0_),
            .carryout(\POWERLED.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_6_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11777),
            .in3(N__11129),
            .lcout(\POWERLED.mult1_un47_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_6_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11711),
            .in3(N__11117),
            .lcout(\POWERLED.mult1_un47_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_6_3  (
            .in0(_gnd_net_),
            .in1(N__18376),
            .in2(N__11729),
            .in3(N__11105),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_4_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_4_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_4_6_4  (
            .in0(_gnd_net_),
            .in1(N__18377),
            .in2(N__11720),
            .in3(N__11102),
            .lcout(\POWERLED.mult1_un47_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_6_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_6_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_6_5  (
            .in0(_gnd_net_),
            .in1(N__11099),
            .in2(_gnd_net_),
            .in3(N__11093),
            .lcout(\POWERLED.mult1_un54_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_4_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_4_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_4_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13183),
            .lcout(\POWERLED.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_6_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11495),
            .lcout(\POWERLED.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(N__13160),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_7_0_),
            .carryout(\POWERLED.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(N__11759),
            .in2(N__11176),
            .in3(N__11264),
            .lcout(\POWERLED.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_4_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_4_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_4_7_2  (
            .in0(_gnd_net_),
            .in1(N__11172),
            .in2(N__11261),
            .in3(N__11237),
            .lcout(\POWERLED.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_4_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_4_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_4_7_3  (
            .in0(_gnd_net_),
            .in1(N__11234),
            .in2(N__11501),
            .in3(N__11213),
            .lcout(\POWERLED.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_4_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_4_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(N__11499),
            .in2(N__11210),
            .in3(N__11189),
            .lcout(\POWERLED.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_4_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_4_7_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_4_7_5  (
            .in0(N__11448),
            .in1(N__11186),
            .in2(N__11177),
            .in3(N__11150),
            .lcout(\POWERLED.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_4_7_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_4_7_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_4_7_6  (
            .in0(N__11513),
            .in1(N__11500),
            .in2(N__11480),
            .in3(N__11468),
            .lcout(\POWERLED.mult1_un61_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_4_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_4_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_4_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11447),
            .lcout(\POWERLED.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_8_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12949),
            .lcout(\POWERLED.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_4_9_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_4_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12731),
            .lcout(\POWERLED.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_4_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_4_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13006),
            .lcout(\POWERLED.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12983),
            .lcout(\POWERLED.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIV4PD6_1_LC_4_10_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIV4PD6_1_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIV4PD6_1_LC_4_10_1 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \POWERLED.func_state_RNIV4PD6_1_LC_4_10_1  (
            .in0(N__13706),
            .in1(N__15302),
            .in2(_gnd_net_),
            .in3(N__13529),
            .lcout(\POWERLED.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_7_l_fx_LC_4_11_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_7_l_fx_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_7_l_fx_LC_4_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_7_l_fx_LC_4_11_5  (
            .in0(N__11360),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11331),
            .lcout(\POWERLED.mult1_un145_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_4_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_4_11_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_4_11_6  (
            .in0(N__11332),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_EN_i_i_i_LC_4_12_3 .C_ON=1'b0;
    defparam \POWERLED.VCCST_EN_i_i_i_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_EN_i_i_i_LC_4_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.VCCST_EN_i_i_i_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15019),
            .lcout(v5s_enn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_12_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14127),
            .lcout(\POWERLED.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_4_12_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_4_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14753),
            .lcout(\POWERLED.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_1_LC_4_13_2 .C_ON=1'b0;
    defparam \POWERLED.count_1_LC_4_13_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_1_LC_4_13_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \POWERLED.count_1_LC_4_13_2  (
            .in0(N__12015),
            .in1(N__12040),
            .in2(_gnd_net_),
            .in3(N__20123),
            .lcout(\POWERLED.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20615),
            .ce(),
            .sr(N__12524));
    defparam \POWERLED.count_0_LC_4_13_6 .C_ON=1'b0;
    defparam \POWERLED.count_0_LC_4_13_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_0_LC_4_13_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.count_0_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__12039),
            .in2(_gnd_net_),
            .in3(N__20122),
            .lcout(\POWERLED.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20615),
            .ce(),
            .sr(N__12524));
    defparam \POWERLED.pwm_out_RNO_4_LC_4_14_0 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_4_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_4_LC_4_14_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.pwm_out_RNO_4_LC_4_14_0  (
            .in0(N__12468),
            .in1(N__11952),
            .in2(_gnd_net_),
            .in3(N__11982),
            .lcout(),
            .ltout(\POWERLED.un1_countlt6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_2_LC_4_14_1 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_2_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_2_LC_4_14_1 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \POWERLED.pwm_out_RNO_2_LC_4_14_1  (
            .in0(N__12441),
            .in1(N__11627),
            .in2(N__11531),
            .in3(N__12411),
            .lcout(),
            .ltout(\POWERLED.g0_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_0_LC_4_14_2 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_0_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_0_LC_4_14_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.pwm_out_RNO_0_LC_4_14_2  (
            .in0(N__12282),
            .in1(N__12384),
            .in2(N__11528),
            .in3(N__11639),
            .lcout(\POWERLED.un1_count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNID4E61_7_LC_4_14_3 .C_ON=1'b0;
    defparam \POWERLED.count_RNID4E61_7_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNID4E61_7_LC_4_14_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_RNID4E61_7_LC_4_14_3  (
            .in0(N__12320),
            .in1(N__12347),
            .in2(N__12386),
            .in3(N__12281),
            .lcout(),
            .ltout(\POWERLED.un1_countlto15_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI6IPJ2_5_LC_4_14_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI6IPJ2_5_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI6IPJ2_5_LC_4_14_4 .LUT_INIT=16'b1111000001110000;
    LogicCell40 \POWERLED.count_RNI6IPJ2_5_LC_4_14_4  (
            .in0(N__12410),
            .in1(N__12440),
            .in2(N__11642),
            .in3(N__11633),
            .lcout(\POWERLED.un1_countlto15_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_1_LC_4_14_5 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_1_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_1_LC_4_14_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.pwm_out_RNO_1_LC_4_14_5  (
            .in0(N__12222),
            .in1(N__12254),
            .in2(_gnd_net_),
            .in3(N__12348),
            .lcout(\POWERLED.g0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNICO6R_2_LC_4_14_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNICO6R_2_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNICO6R_2_LC_4_14_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.count_RNICO6R_2_LC_4_14_6  (
            .in0(N__12467),
            .in1(N__11951),
            .in2(_gnd_net_),
            .in3(N__11981),
            .lcout(\POWERLED.un1_countlt6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_3_LC_4_15_2 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_3_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_3_LC_4_15_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.pwm_out_RNO_3_LC_4_15_2  (
            .in0(N__12621),
            .in1(N__12591),
            .in2(N__12325),
            .in3(N__12551),
            .lcout(\POWERLED.g0_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_esr_RNIBHMO_15_LC_4_15_3 .C_ON=1'b0;
    defparam \POWERLED.count_esr_RNIBHMO_15_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_esr_RNIBHMO_15_LC_4_15_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.count_esr_RNIBHMO_15_LC_4_15_3  (
            .in0(N__12552),
            .in1(N__12590),
            .in2(_gnd_net_),
            .in3(N__12620),
            .lcout(),
            .ltout(\POWERLED.un1_countlto15_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIOVT24_11_LC_4_15_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNIOVT24_11_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIOVT24_11_LC_4_15_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.count_RNIOVT24_11_LC_4_15_4  (
            .in0(N__12221),
            .in1(N__12255),
            .in2(N__11621),
            .in3(N__11618),
            .lcout(\POWERLED.count_RNIOVT24Z0Z_11 ),
            .ltout(\POWERLED.count_RNIOVT24Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNI75RB5_0_LC_4_15_5 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI75RB5_0_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI75RB5_0_LC_4_15_5 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \POWERLED.curr_state_RNI75RB5_0_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__11603),
            .in2(N__11576),
            .in3(N__20063),
            .lcout(\POWERLED.curr_state_RNI75RB5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_esr_RNO_0_15_LC_4_16_0 .C_ON=1'b0;
    defparam \POWERLED.count_esr_RNO_0_15_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_esr_RNO_0_15_LC_4_16_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \POWERLED.count_esr_RNO_0_15_LC_4_16_0  (
            .in0(N__12514),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20066),
            .lcout(\POWERLED.N_65_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_0_LC_5_1_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_0_LC_5_1_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_0_LC_5_1_2 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \HDA_STRAP.count_0_LC_5_1_2  (
            .in0(N__15807),
            .in1(N__15737),
            .in2(N__15901),
            .in3(N__12488),
            .lcout(\HDA_STRAP.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20443),
            .ce(N__19784),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_1_LC_5_1_7 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_1_LC_5_1_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_1_LC_5_1_7 .LUT_INIT=16'b0000100011111000;
    LogicCell40 \HDA_STRAP.curr_state_1_LC_5_1_7  (
            .in0(N__15736),
            .in1(N__15808),
            .in2(N__15900),
            .in3(N__11702),
            .lcout(\HDA_STRAP.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20443),
            .ce(N__19784),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_11_LC_5_2_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_11_LC_5_2_0 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_11_LC_5_2_0 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \HDA_STRAP.count_11_LC_5_2_0  (
            .in0(N__15787),
            .in1(N__15734),
            .in2(N__15899),
            .in3(N__12635),
            .lcout(\HDA_STRAP.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20467),
            .ce(N__19763),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_2_LC_5_2_1 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_2_LC_5_2_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_2_LC_5_2_1 .LUT_INIT=16'b0010111000001100;
    LogicCell40 \HDA_STRAP.curr_state_2_LC_5_2_1  (
            .in0(N__11701),
            .in1(N__11689),
            .in2(N__14036),
            .in3(N__15872),
            .lcout(\HDA_STRAP.curr_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20467),
            .ce(N__19763),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.HDA_SDO_FPGA_LC_5_2_7 .C_ON=1'b0;
    defparam \HDA_STRAP.HDA_SDO_FPGA_LC_5_2_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.HDA_SDO_FPGA_LC_5_2_7 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \HDA_STRAP.HDA_SDO_FPGA_LC_5_2_7  (
            .in0(N__15788),
            .in1(N__15868),
            .in2(_gnd_net_),
            .in3(N__11690),
            .lcout(hda_sdo_atp),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20467),
            .ce(N__19763),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIFHLJ_0_0_LC_5_5_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIFHLJ_0_0_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIFHLJ_0_0_LC_5_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNIFHLJ_0_0_LC_5_5_0  (
            .in0(_gnd_net_),
            .in1(N__14604),
            .in2(N__14110),
            .in3(N__14177),
            .lcout(\POWERLED.un1_dutycycle_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI16B71_5_LC_5_5_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI16B71_5_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI16B71_5_LC_5_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI16B71_5_LC_5_5_1  (
            .in0(N__12697),
            .in1(N__14530),
            .in2(N__14751),
            .in3(N__14088),
            .lcout(\POWERLED.dutycycle_RNI16B71Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_5_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_5_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12811),
            .lcout(\POWERLED.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_5_5_3 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_5_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13114),
            .lcout(\POWERLED.un1_dutycycle_1_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNIMOAE_5_LC_5_5_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNIMOAE_5_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNIMOAE_5_LC_5_5_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_fast_RNIMOAE_5_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(N__16081),
            .in2(_gnd_net_),
            .in3(N__13041),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_1_19_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIEJ021_4_LC_5_5_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIEJ021_4_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIEJ021_4_LC_5_5_5 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \POWERLED.dutycycle_RNIEJ021_4_LC_5_5_5  (
            .in0(N__14605),
            .in1(N__14398),
            .in2(N__11645),
            .in3(N__14666),
            .lcout(\POWERLED.dutycycle_RNIEJ021Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_5_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_5_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_5_6  (
            .in0(N__12793),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIFHLJ_0_LC_5_6_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIFHLJ_0_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIFHLJ_0_LC_5_6_0 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_RNIFHLJ_0_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(N__14606),
            .in2(N__14111),
            .in3(N__14178),
            .lcout(\POWERLED.dutycycle_RNIFHLJZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_LC_5_6_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_1_LC_5_6_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \POWERLED.dutycycle_1_LC_5_6_2  (
            .in0(N__16769),
            .in1(N__11744),
            .in2(_gnd_net_),
            .in3(N__14051),
            .lcout(\POWERLED.dutycycleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20471),
            .ce(N__19773),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_0_LC_5_6_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_0_LC_5_6_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_0_LC_5_6_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \POWERLED.dutycycle_0_LC_5_6_5  (
            .in0(N__11743),
            .in1(N__16770),
            .in2(_gnd_net_),
            .in3(N__14144),
            .lcout(\POWERLED.dutycycleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20471),
            .ce(N__19773),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNIVCSK_5_LC_5_6_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNIVCSK_5_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNIVCSK_5_LC_5_6_6 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_fast_RNIVCSK_5_LC_5_6_6  (
            .in0(_gnd_net_),
            .in1(N__14736),
            .in2(N__14112),
            .in3(N__13042),
            .lcout(\POWERLED.dutycycle_fast_RNIVCSKZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_5_LC_5_6_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_5_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_fast_5_LC_5_6_7 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \POWERLED.dutycycle_fast_5_LC_5_6_7  (
            .in0(N__13430),
            .in1(N__16771),
            .in2(N__13593),
            .in3(N__14486),
            .lcout(\POWERLED.dutycycle_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20471),
            .ce(N__19773),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_7_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_7_0 .LUT_INIT=16'b1111110000000011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(N__13069),
            .in2(N__13097),
            .in3(N__13051),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_5_7_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_5_7_1 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_5_7_1  (
            .in0(N__13052),
            .in1(_gnd_net_),
            .in2(N__13073),
            .in3(N__13095),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_7_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_7_2 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13096),
            .in3(N__13068),
            .lcout(\POWERLED.mult1_un47_sum_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_5_7_3 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_5_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13088),
            .lcout(\POWERLED.un1_dutycycle_1_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_5_7_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_5_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_5_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13156),
            .lcout(\POWERLED.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_5_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_5_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_5_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13135),
            .lcout(\POWERLED.mult1_un54_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI4I7Q_0_5_LC_5_8_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI4I7Q_0_5_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI4I7Q_0_5_LC_5_8_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI4I7Q_0_5_LC_5_8_0  (
            .in0(N__14123),
            .in1(N__14196),
            .in2(N__14532),
            .in3(N__14444),
            .lcout(\POWERLED.N_234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_5_LC_5_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_5_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_5_LC_5_8_1 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \POWERLED.dutycycle_5_LC_5_8_1  (
            .in0(N__16773),
            .in1(N__13421),
            .in2(N__13594),
            .in3(N__14485),
            .lcout(\POWERLED.dutycycleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20564),
            .ce(N__19798),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6NI81_5_LC_5_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6NI81_5_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6NI81_5_LC_5_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI6NI81_5_LC_5_8_2  (
            .in0(N__13021),
            .in1(N__16242),
            .in2(N__14531),
            .in3(N__14443),
            .lcout(\POWERLED.dutycycle_RNI6NI81Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_6_LC_5_8_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_6_LC_5_8_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_6_LC_5_8_3 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \POWERLED.dutycycle_6_LC_5_8_3  (
            .in0(N__16774),
            .in1(N__13422),
            .in2(N__13595),
            .in3(N__14416),
            .lcout(\POWERLED.dutycycleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20564),
            .ce(N__19798),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_6_LC_5_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_6_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_fast_6_LC_5_8_4 .LUT_INIT=16'b1111110010101010;
    LogicCell40 \POWERLED.dutycycle_fast_6_LC_5_8_4  (
            .in0(N__14417),
            .in1(N__13586),
            .in2(N__13429),
            .in3(N__16775),
            .lcout(\POWERLED.dutycycle_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20564),
            .ce(N__19798),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJNBA1_6_LC_5_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJNBA1_6_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJNBA1_6_LC_5_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNIJNBA1_6_LC_5_8_6  (
            .in0(N__13198),
            .in1(N__14442),
            .in2(N__16292),
            .in3(N__14385),
            .lcout(\POWERLED.dutycycle_RNIJNBA1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNILMLM_6_LC_5_8_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNILMLM_6_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNILMLM_6_LC_5_8_7 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_fast_RNILMLM_6_LC_5_8_7  (
            .in0(_gnd_net_),
            .in1(N__16288),
            .in2(N__14397),
            .in3(N__13218),
            .lcout(\POWERLED.dutycycle_fast_RNILMLMZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_0_LC_5_9_0 .C_ON=1'b1;
    defparam \POWERLED.count_off_0_LC_5_9_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_0_LC_5_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_0_LC_5_9_0  (
            .in0(N__12062),
            .in1(N__11842),
            .in2(N__13457),
            .in3(N__13456),
            .lcout(\POWERLED.count_offZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\POWERLED.un1_count_off_1_cry_0 ),
            .clk(N__20585),
            .ce(N__19797),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_1_LC_5_9_1 .C_ON=1'b1;
    defparam \POWERLED.count_off_1_LC_5_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_1_LC_5_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_1_LC_5_9_1  (
            .in0(N__12116),
            .in1(N__11869),
            .in2(_gnd_net_),
            .in3(N__11801),
            .lcout(\POWERLED.count_offZ0Z_1 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_0 ),
            .carryout(\POWERLED.un1_count_off_1_cry_1 ),
            .clk(N__20585),
            .ce(N__19797),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_2_LC_5_9_2 .C_ON=1'b1;
    defparam \POWERLED.count_off_2_LC_5_9_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_2_LC_5_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_2_LC_5_9_2  (
            .in0(N__12063),
            .in1(N__13325),
            .in2(_gnd_net_),
            .in3(N__11798),
            .lcout(\POWERLED.count_offZ0Z_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_1 ),
            .carryout(\POWERLED.un1_count_off_1_cry_2 ),
            .clk(N__20585),
            .ce(N__19797),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_3_LC_5_9_3 .C_ON=1'b1;
    defparam \POWERLED.count_off_3_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_3_LC_5_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_3_LC_5_9_3  (
            .in0(N__12117),
            .in1(N__13367),
            .in2(_gnd_net_),
            .in3(N__11795),
            .lcout(\POWERLED.count_offZ0Z_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_2 ),
            .carryout(\POWERLED.un1_count_off_1_cry_3 ),
            .clk(N__20585),
            .ce(N__19797),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_4_LC_5_9_4 .C_ON=1'b1;
    defparam \POWERLED.count_off_4_LC_5_9_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_4_LC_5_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_4_LC_5_9_4  (
            .in0(N__12119),
            .in1(N__13339),
            .in2(_gnd_net_),
            .in3(N__11792),
            .lcout(\POWERLED.count_offZ0Z_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_3 ),
            .carryout(\POWERLED.un1_count_off_1_cry_4 ),
            .clk(N__20585),
            .ce(N__19797),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_5_LC_5_9_5 .C_ON=1'b1;
    defparam \POWERLED.count_off_5_LC_5_9_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_5_LC_5_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_5_LC_5_9_5  (
            .in0(N__12065),
            .in1(N__12148),
            .in2(_gnd_net_),
            .in3(N__11789),
            .lcout(\POWERLED.count_offZ0Z_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_4 ),
            .carryout(\POWERLED.un1_count_off_1_cry_5 ),
            .clk(N__20585),
            .ce(N__19797),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_6_LC_5_9_6 .C_ON=1'b1;
    defparam \POWERLED.count_off_6_LC_5_9_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_6_LC_5_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_6_LC_5_9_6  (
            .in0(N__12064),
            .in1(N__12178),
            .in2(_gnd_net_),
            .in3(N__11786),
            .lcout(\POWERLED.count_offZ0Z_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_5 ),
            .carryout(\POWERLED.un1_count_off_1_cry_6 ),
            .clk(N__20585),
            .ce(N__19797),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_7_LC_5_9_7 .C_ON=1'b1;
    defparam \POWERLED.count_off_7_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_7_LC_5_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_7_LC_5_9_7  (
            .in0(N__12118),
            .in1(N__13354),
            .in2(_gnd_net_),
            .in3(N__11783),
            .lcout(\POWERLED.count_offZ0Z_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_6 ),
            .carryout(\POWERLED.un1_count_off_1_cry_7 ),
            .clk(N__20585),
            .ce(N__19797),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_8_LC_5_10_0 .C_ON=1'b1;
    defparam \POWERLED.count_off_8_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_8_LC_5_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_8_LC_5_10_0  (
            .in0(N__12111),
            .in1(N__12193),
            .in2(_gnd_net_),
            .in3(N__11780),
            .lcout(\POWERLED.count_offZ0Z_8 ),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\POWERLED.un1_count_off_1_cry_8 ),
            .clk(N__20604),
            .ce(N__19807),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_9_LC_5_10_1 .C_ON=1'b1;
    defparam \POWERLED.count_off_9_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_9_LC_5_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_9_LC_5_10_1  (
            .in0(N__12114),
            .in1(N__12163),
            .in2(_gnd_net_),
            .in3(N__11930),
            .lcout(\POWERLED.count_offZ0Z_9 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_8 ),
            .carryout(\POWERLED.un1_count_off_1_cry_9 ),
            .clk(N__20604),
            .ce(N__19807),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_10_LC_5_10_2 .C_ON=1'b1;
    defparam \POWERLED.count_off_10_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_10_LC_5_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_10_LC_5_10_2  (
            .in0(N__12108),
            .in1(N__11813),
            .in2(_gnd_net_),
            .in3(N__11927),
            .lcout(\POWERLED.count_offZ0Z_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_9 ),
            .carryout(\POWERLED.un1_count_off_1_cry_10 ),
            .clk(N__20604),
            .ce(N__19807),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_11_LC_5_10_3 .C_ON=1'b1;
    defparam \POWERLED.count_off_11_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_11_LC_5_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_11_LC_5_10_3  (
            .in0(N__12112),
            .in1(N__11855),
            .in2(_gnd_net_),
            .in3(N__11924),
            .lcout(\POWERLED.count_offZ0Z_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_10 ),
            .carryout(\POWERLED.un1_count_off_1_cry_11 ),
            .clk(N__20604),
            .ce(N__19807),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_12_LC_5_10_4 .C_ON=1'b1;
    defparam \POWERLED.count_off_12_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_12_LC_5_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_12_LC_5_10_4  (
            .in0(N__12109),
            .in1(N__11909),
            .in2(_gnd_net_),
            .in3(N__11921),
            .lcout(\POWERLED.count_offZ0Z_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_11 ),
            .carryout(\POWERLED.un1_count_off_1_cry_12 ),
            .clk(N__20604),
            .ce(N__19807),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_13_LC_5_10_5 .C_ON=1'b1;
    defparam \POWERLED.count_off_13_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_13_LC_5_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_13_LC_5_10_5  (
            .in0(N__12113),
            .in1(N__11897),
            .in2(_gnd_net_),
            .in3(N__11918),
            .lcout(\POWERLED.count_offZ0Z_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_12 ),
            .carryout(\POWERLED.un1_count_off_1_cry_13 ),
            .clk(N__20604),
            .ce(N__19807),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_14_LC_5_10_6 .C_ON=1'b1;
    defparam \POWERLED.count_off_14_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_14_LC_5_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_14_LC_5_10_6  (
            .in0(N__12110),
            .in1(N__11827),
            .in2(_gnd_net_),
            .in3(N__11915),
            .lcout(\POWERLED.count_offZ0Z_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_13 ),
            .carryout(\POWERLED.un1_count_off_1_cry_14 ),
            .clk(N__20604),
            .ce(N__19807),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_15_LC_5_10_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_15_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_15_LC_5_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \POWERLED.count_off_15_LC_5_10_7  (
            .in0(N__12115),
            .in1(N__11884),
            .in2(_gnd_net_),
            .in3(N__11912),
            .lcout(\POWERLED.count_offZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20604),
            .ce(N__19807),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIAJ6S_15_LC_5_11_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIAJ6S_15_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIAJ6S_15_LC_5_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNIAJ6S_15_LC_5_11_0  (
            .in0(N__11908),
            .in1(N__11896),
            .in2(N__11885),
            .in3(N__11870),
            .lcout(\POWERLED.func_state_ns_0_a2_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI4D6S_10_LC_5_11_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI4D6S_10_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI4D6S_10_LC_5_11_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI4D6S_10_LC_5_11_1  (
            .in0(N__11854),
            .in1(N__11843),
            .in2(N__11828),
            .in3(N__11812),
            .lcout(\POWERLED.func_state_ns_0_a2_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI8GP11_5_LC_5_11_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI8GP11_5_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI8GP11_5_LC_5_11_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.count_off_RNI8GP11_5_LC_5_11_2  (
            .in0(N__12194),
            .in1(N__12179),
            .in2(N__12164),
            .in3(N__12149),
            .lcout(),
            .ltout(\POWERLED.func_state_ns_0_a2_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIIKVR3_10_LC_5_11_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIIKVR3_10_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIIKVR3_10_LC_5_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.count_off_RNIIKVR3_10_LC_5_11_3  (
            .in0(N__12134),
            .in1(N__12128),
            .in2(N__12122),
            .in3(N__13313),
            .lcout(\POWERLED.count_off_RNIIKVR3Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIHPO9A_0_LC_5_11_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIHPO9A_0_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIHPO9A_0_LC_5_11_5 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \POWERLED.func_state_RNIHPO9A_0_LC_5_11_5  (
            .in0(N__13698),
            .in1(N__14901),
            .in2(_gnd_net_),
            .in3(N__13521),
            .lcout(\POWERLED.count_off_0_sqmuxa ),
            .ltout(\POWERLED.count_off_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI9LL3G_1_LC_5_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI9LL3G_1_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI9LL3G_1_LC_5_11_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \POWERLED.func_state_RNI9LL3G_1_LC_5_11_6  (
            .in0(N__14933),
            .in1(_gnd_net_),
            .in2(N__12068),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_85_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_LC_5_12_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_1_LC_5_12_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \POWERLED.func_state_1_LC_5_12_1  (
            .in0(N__13712),
            .in1(N__13528),
            .in2(N__13643),
            .in3(N__14906),
            .lcout(\POWERLED.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20605),
            .ce(N__19808),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_1_cry_1_c_LC_5_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_1_cry_1_c_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_1_cry_1_c_LC_5_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_1_cry_1_c_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__12038),
            .in2(N__12016),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\POWERLED.un1_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_2_LC_5_14_1 .C_ON=1'b1;
    defparam \POWERLED.count_2_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_2_LC_5_14_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_2_LC_5_14_1  (
            .in0(N__20124),
            .in1(N__11986),
            .in2(_gnd_net_),
            .in3(N__11963),
            .lcout(\POWERLED.countZ0Z_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_1 ),
            .carryout(\POWERLED.un1_count_1_cry_2 ),
            .clk(N__20596),
            .ce(),
            .sr(N__12519));
    defparam \POWERLED.count_3_LC_5_14_2 .C_ON=1'b1;
    defparam \POWERLED.count_3_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_3_LC_5_14_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_3_LC_5_14_2  (
            .in0(N__20107),
            .in1(N__11956),
            .in2(_gnd_net_),
            .in3(N__11933),
            .lcout(\POWERLED.countZ0Z_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_2 ),
            .carryout(\POWERLED.un1_count_1_cry_3 ),
            .clk(N__20596),
            .ce(),
            .sr(N__12519));
    defparam \POWERLED.count_4_LC_5_14_3 .C_ON=1'b1;
    defparam \POWERLED.count_4_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_4_LC_5_14_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_4_LC_5_14_3  (
            .in0(N__20125),
            .in1(N__12472),
            .in2(_gnd_net_),
            .in3(N__12449),
            .lcout(\POWERLED.countZ0Z_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_3 ),
            .carryout(\POWERLED.un1_count_1_cry_4 ),
            .clk(N__20596),
            .ce(),
            .sr(N__12519));
    defparam \POWERLED.count_5_LC_5_14_4 .C_ON=1'b1;
    defparam \POWERLED.count_5_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_5_LC_5_14_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_5_LC_5_14_4  (
            .in0(N__20108),
            .in1(N__12442),
            .in2(_gnd_net_),
            .in3(N__12419),
            .lcout(\POWERLED.countZ0Z_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_4 ),
            .carryout(\POWERLED.un1_count_1_cry_5 ),
            .clk(N__20596),
            .ce(),
            .sr(N__12519));
    defparam \POWERLED.count_6_LC_5_14_5 .C_ON=1'b1;
    defparam \POWERLED.count_6_LC_5_14_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_6_LC_5_14_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_6_LC_5_14_5  (
            .in0(N__20126),
            .in1(N__12412),
            .in2(_gnd_net_),
            .in3(N__12389),
            .lcout(\POWERLED.countZ0Z_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_5 ),
            .carryout(\POWERLED.un1_count_1_cry_6 ),
            .clk(N__20596),
            .ce(),
            .sr(N__12519));
    defparam \POWERLED.count_7_LC_5_14_6 .C_ON=1'b1;
    defparam \POWERLED.count_7_LC_5_14_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_7_LC_5_14_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_7_LC_5_14_6  (
            .in0(N__20109),
            .in1(N__12377),
            .in2(_gnd_net_),
            .in3(N__12356),
            .lcout(\POWERLED.countZ0Z_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_6 ),
            .carryout(\POWERLED.un1_count_1_cry_7 ),
            .clk(N__20596),
            .ce(),
            .sr(N__12519));
    defparam \POWERLED.count_8_LC_5_14_7 .C_ON=1'b1;
    defparam \POWERLED.count_8_LC_5_14_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_8_LC_5_14_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_8_LC_5_14_7  (
            .in0(N__20127),
            .in1(N__12352),
            .in2(_gnd_net_),
            .in3(N__12329),
            .lcout(\POWERLED.countZ0Z_8 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_7 ),
            .carryout(\POWERLED.un1_count_1_cry_8 ),
            .clk(N__20596),
            .ce(),
            .sr(N__12519));
    defparam \POWERLED.count_9_LC_5_15_0 .C_ON=1'b1;
    defparam \POWERLED.count_9_LC_5_15_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_9_LC_5_15_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_9_LC_5_15_0  (
            .in0(N__20141),
            .in1(N__12321),
            .in2(_gnd_net_),
            .in3(N__12293),
            .lcout(\POWERLED.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\POWERLED.un1_count_1_cry_9 ),
            .clk(N__20630),
            .ce(),
            .sr(N__12515));
    defparam \POWERLED.count_10_LC_5_15_1 .C_ON=1'b1;
    defparam \POWERLED.count_10_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_10_LC_5_15_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_10_LC_5_15_1  (
            .in0(N__20150),
            .in1(N__12286),
            .in2(_gnd_net_),
            .in3(N__12263),
            .lcout(\POWERLED.countZ0Z_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_9 ),
            .carryout(\POWERLED.un1_count_1_cry_10 ),
            .clk(N__20630),
            .ce(),
            .sr(N__12515));
    defparam \POWERLED.count_11_LC_5_15_2 .C_ON=1'b1;
    defparam \POWERLED.count_11_LC_5_15_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_11_LC_5_15_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_11_LC_5_15_2  (
            .in0(N__20139),
            .in1(N__12256),
            .in2(_gnd_net_),
            .in3(N__12230),
            .lcout(\POWERLED.countZ0Z_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_10 ),
            .carryout(\POWERLED.un1_count_1_cry_11 ),
            .clk(N__20630),
            .ce(),
            .sr(N__12515));
    defparam \POWERLED.count_12_LC_5_15_3 .C_ON=1'b1;
    defparam \POWERLED.count_12_LC_5_15_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_12_LC_5_15_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_12_LC_5_15_3  (
            .in0(N__20151),
            .in1(N__12223),
            .in2(_gnd_net_),
            .in3(N__12197),
            .lcout(\POWERLED.countZ0Z_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_11 ),
            .carryout(\POWERLED.un1_count_1_cry_12 ),
            .clk(N__20630),
            .ce(),
            .sr(N__12515));
    defparam \POWERLED.count_13_LC_5_15_4 .C_ON=1'b1;
    defparam \POWERLED.count_13_LC_5_15_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_13_LC_5_15_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_13_LC_5_15_4  (
            .in0(N__20140),
            .in1(N__12622),
            .in2(_gnd_net_),
            .in3(N__12599),
            .lcout(\POWERLED.countZ0Z_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_12 ),
            .carryout(\POWERLED.un1_count_1_cry_13 ),
            .clk(N__20630),
            .ce(),
            .sr(N__12515));
    defparam \POWERLED.count_14_LC_5_15_5 .C_ON=1'b1;
    defparam \POWERLED.count_14_LC_5_15_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_14_LC_5_15_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_14_LC_5_15_5  (
            .in0(N__20152),
            .in1(N__12592),
            .in2(_gnd_net_),
            .in3(N__12566),
            .lcout(\POWERLED.countZ0Z_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_13 ),
            .carryout(\POWERLED.un1_count_1_cry_14 ),
            .clk(N__20630),
            .ce(),
            .sr(N__12515));
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_15_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(N__18301),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_14 ),
            .carryout(\POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_5_15_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_5_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__18318),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryout(\POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_esr_15_LC_5_16_0 .C_ON=1'b0;
    defparam \POWERLED.count_esr_15_LC_5_16_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_esr_15_LC_5_16_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.count_esr_15_LC_5_16_0  (
            .in0(_gnd_net_),
            .in1(N__12556),
            .in2(_gnd_net_),
            .in3(N__12563),
            .lcout(\POWERLED.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20635),
            .ce(N__12533),
            .sr(N__12520));
    defparam \HDA_STRAP.count_RNO_0_0_LC_6_1_0 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_0_LC_6_1_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_0_LC_6_1_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_0_LC_6_1_0  (
            .in0(_gnd_net_),
            .in1(N__13874),
            .in2(N__13928),
            .in3(N__13927),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_6_1_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_1_LC_6_1_1 .C_ON=1'b1;
    defparam \HDA_STRAP.count_1_LC_6_1_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_1_LC_6_1_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_1_LC_6_1_1  (
            .in0(_gnd_net_),
            .in1(N__13901),
            .in2(_gnd_net_),
            .in3(N__12482),
            .lcout(\HDA_STRAP.countZ0Z_1 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_0 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_1 ),
            .clk(N__20205),
            .ce(N__19712),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_2_LC_6_1_2 .C_ON=1'b1;
    defparam \HDA_STRAP.count_2_LC_6_1_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_2_LC_6_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_2_LC_6_1_2  (
            .in0(_gnd_net_),
            .in1(N__13913),
            .in2(_gnd_net_),
            .in3(N__12479),
            .lcout(\HDA_STRAP.countZ0Z_2 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_1 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_2 ),
            .clk(N__20205),
            .ce(N__19712),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_3_LC_6_1_3 .C_ON=1'b1;
    defparam \HDA_STRAP.count_3_LC_6_1_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_3_LC_6_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_3_LC_6_1_3  (
            .in0(_gnd_net_),
            .in1(N__13888),
            .in2(_gnd_net_),
            .in3(N__12659),
            .lcout(\HDA_STRAP.countZ0Z_3 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_2 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_3 ),
            .clk(N__20205),
            .ce(N__19712),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_4_LC_6_1_4 .C_ON=1'b1;
    defparam \HDA_STRAP.count_4_LC_6_1_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_4_LC_6_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_4_LC_6_1_4  (
            .in0(_gnd_net_),
            .in1(N__13766),
            .in2(_gnd_net_),
            .in3(N__12656),
            .lcout(\HDA_STRAP.countZ0Z_4 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_3 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_4 ),
            .clk(N__20205),
            .ce(N__19712),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_5_LC_6_1_5 .C_ON=1'b1;
    defparam \HDA_STRAP.count_5_LC_6_1_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_5_LC_6_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_5_LC_6_1_5  (
            .in0(_gnd_net_),
            .in1(N__13793),
            .in2(_gnd_net_),
            .in3(N__12653),
            .lcout(\HDA_STRAP.countZ0Z_5 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_4 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_5 ),
            .clk(N__20205),
            .ce(N__19712),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_6_LC_6_1_6 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_6_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_6_LC_6_1_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_6_LC_6_1_6  (
            .in0(_gnd_net_),
            .in1(N__15686),
            .in2(_gnd_net_),
            .in3(N__12650),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_5 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_7_LC_6_1_7 .C_ON=1'b1;
    defparam \HDA_STRAP.count_7_LC_6_1_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_7_LC_6_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_7_LC_6_1_7  (
            .in0(_gnd_net_),
            .in1(N__13805),
            .in2(_gnd_net_),
            .in3(N__12647),
            .lcout(\HDA_STRAP.countZ0Z_7 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_6 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_7 ),
            .clk(N__20205),
            .ce(N__19712),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_8_LC_6_2_0 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_8_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_8_LC_6_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_8_LC_6_2_0  (
            .in0(_gnd_net_),
            .in1(N__13958),
            .in2(_gnd_net_),
            .in3(N__12644),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_6_2_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_9_LC_6_2_1 .C_ON=1'b1;
    defparam \HDA_STRAP.count_9_LC_6_2_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_9_LC_6_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_9_LC_6_2_1  (
            .in0(_gnd_net_),
            .in1(N__13780),
            .in2(_gnd_net_),
            .in3(N__12641),
            .lcout(\HDA_STRAP.countZ0Z_9 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_8 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_9 ),
            .clk(N__20370),
            .ce(N__19741),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_10_LC_6_2_2 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_10_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_10_LC_6_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_10_LC_6_2_2  (
            .in0(_gnd_net_),
            .in1(N__14011),
            .in2(_gnd_net_),
            .in3(N__12638),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_9 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_11_LC_6_2_3 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_11_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_11_LC_6_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_11_LC_6_2_3  (
            .in0(_gnd_net_),
            .in1(N__13753),
            .in2(_gnd_net_),
            .in3(N__12629),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_10 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_12_LC_6_2_4 .C_ON=1'b1;
    defparam \HDA_STRAP.count_12_LC_6_2_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_12_LC_6_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_12_LC_6_2_4  (
            .in0(_gnd_net_),
            .in1(N__13832),
            .in2(_gnd_net_),
            .in3(N__12776),
            .lcout(\HDA_STRAP.countZ0Z_12 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_11 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_12 ),
            .clk(N__20370),
            .ce(N__19741),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_13_LC_6_2_5 .C_ON=1'b1;
    defparam \HDA_STRAP.count_13_LC_6_2_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_13_LC_6_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_13_LC_6_2_5  (
            .in0(_gnd_net_),
            .in1(N__13817),
            .in2(_gnd_net_),
            .in3(N__12773),
            .lcout(\HDA_STRAP.countZ0Z_13 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_12 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_13 ),
            .clk(N__20370),
            .ce(N__19741),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_14_LC_6_2_6 .C_ON=1'b1;
    defparam \HDA_STRAP.count_14_LC_6_2_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_14_LC_6_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_14_LC_6_2_6  (
            .in0(_gnd_net_),
            .in1(N__13859),
            .in2(_gnd_net_),
            .in3(N__12770),
            .lcout(\HDA_STRAP.countZ0Z_14 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_13 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_14 ),
            .clk(N__20370),
            .ce(N__19741),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_15_LC_6_2_7 .C_ON=1'b1;
    defparam \HDA_STRAP.count_15_LC_6_2_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_15_LC_6_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_15_LC_6_2_7  (
            .in0(_gnd_net_),
            .in1(N__13846),
            .in2(_gnd_net_),
            .in3(N__12767),
            .lcout(\HDA_STRAP.countZ0Z_15 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_14 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_15 ),
            .clk(N__20370),
            .ce(N__19741),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_16_LC_6_3_0 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_16_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_16_LC_6_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_16_LC_6_3_0  (
            .in0(_gnd_net_),
            .in1(N__13994),
            .in2(_gnd_net_),
            .in3(N__12764),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_17_LC_6_3_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNO_0_17_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_17_LC_6_3_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \HDA_STRAP.count_RNO_0_17_LC_6_3_1  (
            .in0(_gnd_net_),
            .in1(N__13976),
            .in2(_gnd_net_),
            .in3(N__12761),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIVL3D_0_LC_6_5_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNIVL3D_0_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIVL3D_0_LC_6_5_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \POWERLED.dutycycle_RNIVL3D_0_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(N__14658),
            .in2(N__14194),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_dutycycle_1_axb_0 ),
            .ltout(),
            .carryin(bfn_6_5_0_),
            .carryout(\POWERLED.un1_dutycycle_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_6_5_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_6_5_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12740),
            .in3(N__12707),
            .lcout(\POWERLED.mult1_un138_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_0 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_6_5_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_6_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_6_5_2  (
            .in0(_gnd_net_),
            .in1(N__12704),
            .in2(N__12698),
            .in3(N__12662),
            .lcout(\POWERLED.mult1_un131_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_1 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_6_5_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_6_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_6_5_3  (
            .in0(_gnd_net_),
            .in1(N__14261),
            .in2(N__14278),
            .in3(N__12986),
            .lcout(\POWERLED.mult1_un124_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_2 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_6_5_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_6_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_6_5_4  (
            .in0(_gnd_net_),
            .in1(N__14225),
            .in2(N__14243),
            .in3(N__12962),
            .lcout(\POWERLED.mult1_un117_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_3 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_6_5_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_6_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_6_5_5  (
            .in0(_gnd_net_),
            .in1(N__14219),
            .in2(N__12959),
            .in3(N__12929),
            .lcout(\POWERLED.mult1_un110_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_4 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_6_5_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_6_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_6_5_6  (
            .in0(_gnd_net_),
            .in1(N__12926),
            .in2(N__13025),
            .in3(N__12893),
            .lcout(\POWERLED.mult1_un103_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_5 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_6_5_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_6_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_6_5_7  (
            .in0(_gnd_net_),
            .in1(N__12890),
            .in2(N__13202),
            .in3(N__12851),
            .lcout(\POWERLED.mult1_un96_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_6 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_6_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_6_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__13250),
            .in2(N__13235),
            .in3(N__12821),
            .lcout(\POWERLED.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(\POWERLED.un1_dutycycle_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_6_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_6_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__13271),
            .in2(N__14315),
            .in3(N__12797),
            .lcout(\POWERLED.mult1_un82_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_8 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_6_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_6_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__13289),
            .in2(N__13301),
            .in3(N__12779),
            .lcout(\POWERLED.mult1_un75_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_6_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_6_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__13376),
            .in2(N__16493),
            .in3(N__13163),
            .lcout(\POWERLED.mult1_un68_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_6_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_6_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(N__13385),
            .in2(N__13400),
            .in3(N__13142),
            .lcout(\POWERLED.mult1_un61_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_6_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_6_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_6_6_5  (
            .in0(_gnd_net_),
            .in1(N__13481),
            .in2(N__13946),
            .in3(N__13121),
            .lcout(\POWERLED.mult1_un54_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_6_6_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_6_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(N__13277),
            .in2(N__13937),
            .in3(N__13100),
            .lcout(\POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_6_6_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_6_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_6_6_7  (
            .in0(_gnd_net_),
            .in1(N__13283),
            .in2(N__13493),
            .in3(N__13076),
            .lcout(\POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_14 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_6_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_6_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(N__16128),
            .in2(N__13265),
            .in3(N__13058),
            .lcout(\POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71 ),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(\POWERLED.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_6_7_1 .C_ON=1'b0;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_6_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.CO2_THRU_LUT4_0_LC_6_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13055),
            .lcout(\POWERLED.CO2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNI8MSK_5_LC_6_7_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNI8MSK_5_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNI8MSK_5_LC_6_7_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \POWERLED.dutycycle_fast_RNI8MSK_5_LC_6_7_2  (
            .in0(N__16066),
            .in1(N__14601),
            .in2(_gnd_net_),
            .in3(N__13043),
            .lcout(\POWERLED.dutycycle_fast_RNI8MSKZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIE4FL_9_LC_6_7_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIE4FL_9_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIE4FL_9_LC_6_7_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \POWERLED.dutycycle_RNIE4FL_9_LC_6_7_3  (
            .in0(N__16388),
            .in1(N__16237),
            .in2(_gnd_net_),
            .in3(N__16068),
            .lcout(\POWERLED.dutycycle_RNIE4FLZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI53MG_14_LC_6_7_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI53MG_14_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI53MG_14_LC_6_7_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.dutycycle_RNI53MG_14_LC_6_7_4  (
            .in0(N__16339),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16460),
            .lcout(\POWERLED.dutycycle_RNI53MGZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNI2GSK_6_LC_6_7_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNI2GSK_6_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNI2GSK_6_LC_6_7_5 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_fast_RNI2GSK_6_LC_6_7_5  (
            .in0(_gnd_net_),
            .in1(N__14644),
            .in2(N__13223),
            .in3(N__14722),
            .lcout(\POWERLED.dutycycle_fast_RNI2GSKZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI84C11_14_LC_6_7_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI84C11_14_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI84C11_14_LC_6_7_6 .LUT_INIT=16'b0100101101111000;
    LogicCell40 \POWERLED.dutycycle_RNI84C11_14_LC_6_7_6  (
            .in0(N__16458),
            .in1(N__16389),
            .in2(N__16345),
            .in3(N__16459),
            .lcout(\POWERLED.dutycycle_RNI84C11Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIB1FL_8_LC_6_7_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIB1FL_8_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIB1FL_8_LC_6_7_7 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \POWERLED.dutycycle_RNIB1FL_8_LC_6_7_7  (
            .in0(N__14393),
            .in1(N__16185),
            .in2(_gnd_net_),
            .in3(N__16067),
            .lcout(\POWERLED.dutycycle_RNIB1FLZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI75MG_15_LC_6_8_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI75MG_15_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI75MG_15_LC_6_8_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \POWERLED.dutycycle_RNI75MG_15_LC_6_8_0  (
            .in0(N__16117),
            .in1(_gnd_net_),
            .in2(N__16344),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI75MGZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIM0TE_8_LC_6_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIM0TE_8_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIM0TE_8_LC_6_8_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNIM0TE_8_LC_6_8_1  (
            .in0(_gnd_net_),
            .in1(N__16065),
            .in2(_gnd_net_),
            .in3(N__16167),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_1_34_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIUUB41_6_LC_6_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIUUB41_6_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIUUB41_6_LC_6_8_2 .LUT_INIT=16'b1110000101111000;
    LogicCell40 \POWERLED.dutycycle_RNIUUB41_6_LC_6_8_2  (
            .in0(N__16281),
            .in1(N__14445),
            .in2(N__13256),
            .in3(N__14373),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_1_axb_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJL1R1_6_LC_6_8_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJL1R1_6_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJL1R1_6_LC_6_8_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNIJL1R1_6_LC_6_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13253),
            .in3(N__13246),
            .lcout(\POWERLED.dutycycle_RNIJL1R1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNIBPSK_6_LC_6_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNIBPSK_6_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNIBPSK_6_LC_6_8_4 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \POWERLED.dutycycle_fast_RNIBPSK_6_LC_6_8_4  (
            .in0(N__16231),
            .in1(N__14523),
            .in2(_gnd_net_),
            .in3(N__13222),
            .lcout(\POWERLED.dutycycle_fast_RNIBPSKZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2V0P_10_LC_6_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2V0P_10_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2V0P_10_LC_6_8_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \POWERLED.dutycycle_RNI2V0P_10_LC_6_8_5  (
            .in0(N__16173),
            .in1(N__16330),
            .in2(_gnd_net_),
            .in3(N__16283),
            .lcout(\POWERLED.dutycycle_RNI2V0PZ0Z_10 ),
            .ltout(\POWERLED.dutycycle_RNI2V0PZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI712I1_15_LC_6_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI712I1_15_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI712I1_15_LC_6_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNI712I1_15_LC_6_8_6  (
            .in0(N__16116),
            .in1(N__16172),
            .in2(N__13388),
            .in3(N__16394),
            .lcout(\POWERLED.dutycycle_RNI712I1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQ09G1_10_LC_6_8_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQ09G1_10_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQ09G1_10_LC_6_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNIQ09G1_10_LC_6_8_7  (
            .in0(N__16489),
            .in1(N__16329),
            .in2(N__16184),
            .in3(N__16282),
            .lcout(\POWERLED.dutycycle_RNIQ09G1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_0_2_LC_6_9_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_0_2_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_0_2_LC_6_9_0 .LUT_INIT=16'b0110111011101110;
    LogicCell40 \POWERLED.dutycycle_RNO_0_2_LC_6_9_0  (
            .in0(N__15359),
            .in1(N__15098),
            .in2(N__16590),
            .in3(N__15298),
            .lcout(\POWERLED.dutycycle_lm_0_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIS3P11_2_LC_6_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIS3P11_2_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIS3P11_2_LC_6_9_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \POWERLED.count_off_RNIS3P11_2_LC_6_9_1  (
            .in0(N__13366),
            .in1(N__13355),
            .in2(N__13340),
            .in3(N__13324),
            .lcout(\POWERLED.func_state_ns_0_a2_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI1DHM_6_LC_6_9_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI1DHM_6_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI1DHM_6_LC_6_9_2 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \POWERLED.count_clk_RNI1DHM_6_LC_6_9_2  (
            .in0(N__18055),
            .in1(N__18007),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_368_0_i_i_a6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI1VLG_10_LC_6_9_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI1VLG_10_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI1VLG_10_LC_6_9_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI1VLG_10_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(N__16284),
            .in2(_gnd_net_),
            .in3(N__16448),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_1_44_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIF3561_9_LC_6_9_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIF3561_9_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIF3561_9_LC_6_9_4 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \POWERLED.dutycycle_RNIF3561_9_LC_6_9_4  (
            .in0(N__16082),
            .in1(N__16236),
            .in2(N__13304),
            .in3(N__16393),
            .lcout(\POWERLED.dutycycle_RNIF3561Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIC8C11_15_LC_6_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIC8C11_15_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIC8C11_15_LC_6_9_6 .LUT_INIT=16'b0110001101101100;
    LogicCell40 \POWERLED.dutycycle_RNIC8C11_15_LC_6_9_6  (
            .in0(N__16334),
            .in1(N__16118),
            .in2(N__16466),
            .in3(N__16335),
            .lcout(\POWERLED.dutycycle_RNIC8C11Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI73C11_15_LC_6_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI73C11_15_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI73C11_15_LC_6_9_7 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_RNI73C11_15_LC_6_9_7  (
            .in0(N__16465),
            .in1(N__16168),
            .in2(N__16402),
            .in3(N__16115),
            .lcout(\POWERLED.dutycycle_RNI73C11Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIBR4E9_6_LC_6_10_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIBR4E9_6_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIBR4E9_6_LC_6_10_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.count_clk_RNIBR4E9_6_LC_6_10_1  (
            .in0(N__16676),
            .in1(N__13606),
            .in2(N__13469),
            .in3(N__16630),
            .lcout(\POWERLED.N_177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIAA8L4_0_LC_6_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIAA8L4_0_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIAA8L4_0_LC_6_10_2 .LUT_INIT=16'b0000000000101110;
    LogicCell40 \POWERLED.func_state_RNIAA8L4_0_LC_6_10_2  (
            .in0(N__13548),
            .in1(N__15220),
            .in2(N__14306),
            .in3(N__16000),
            .lcout(\POWERLED.N_200_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIS0FM9_7_LC_6_10_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIS0FM9_7_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIS0FM9_7_LC_6_10_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \POWERLED.count_clk_RNIS0FM9_7_LC_6_10_3  (
            .in0(N__13701),
            .in1(N__16631),
            .in2(N__13442),
            .in3(N__18019),
            .lcout(),
            .ltout(\POWERLED.N_207_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI5LMRL_1_LC_6_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI5LMRL_1_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI5LMRL_1_LC_6_10_4 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \POWERLED.count_clk_RNI5LMRL_1_LC_6_10_4  (
            .in0(N__14762),
            .in1(N__16814),
            .in2(N__13460),
            .in3(N__14926),
            .lcout(\POWERLED.N_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIG4MR5_1_LC_6_10_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIG4MR5_1_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIG4MR5_1_LC_6_10_5 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \POWERLED.func_state_RNIG4MR5_1_LC_6_10_5  (
            .in0(N__15300),
            .in1(N__16652),
            .in2(_gnd_net_),
            .in3(N__15147),
            .lcout(\POWERLED.N_149 ),
            .ltout(\POWERLED.N_149_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIJ13KB_7_LC_6_10_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIJ13KB_7_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIJ13KB_7_LC_6_10_6 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \POWERLED.count_clk_RNIJ13KB_7_LC_6_10_6  (
            .in0(N__18018),
            .in1(N__15651),
            .in2(N__13433),
            .in3(N__15419),
            .lcout(\POWERLED.un2_slp_s3n_2_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5J285_5_LC_6_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5J285_5_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5J285_5_LC_6_10_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \POWERLED.dutycycle_RNI5J285_5_LC_6_10_7  (
            .in0(N__13702),
            .in1(N__16001),
            .in2(N__15446),
            .in3(N__13549),
            .lcout(\POWERLED.N_214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI0AN05_0_0_LC_6_11_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI0AN05_0_0_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI0AN05_0_0_LC_6_11_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.func_state_RNI0AN05_0_0_LC_6_11_0  (
            .in0(N__15996),
            .in1(N__13683),
            .in2(N__15223),
            .in3(N__14304),
            .lcout(\POWERLED.N_248 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_2_0_LC_6_11_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_2_0_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_2_0_LC_6_11_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.func_state_RNO_2_0_LC_6_11_1  (
            .in0(N__15282),
            .in1(N__13556),
            .in2(N__13700),
            .in3(N__15999),
            .lcout(\POWERLED.N_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI1UHM1_0_LC_6_11_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI1UHM1_0_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI1UHM1_0_LC_6_11_2 .LUT_INIT=16'b0000000011000100;
    LogicCell40 \POWERLED.func_state_RNI1UHM1_0_LC_6_11_2  (
            .in0(N__16581),
            .in1(N__15093),
            .in2(N__15224),
            .in3(N__15636),
            .lcout(\POWERLED.N_213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3T7Q4_5_LC_6_11_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3T7Q4_5_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3T7Q4_5_LC_6_11_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \POWERLED.dutycycle_RNI3T7Q4_5_LC_6_11_3  (
            .in0(N__15635),
            .in1(N__13555),
            .in2(N__15445),
            .in3(N__15997),
            .lcout(),
            .ltout(\POWERLED.N_218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNITEUV5_5_LC_6_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNITEUV5_5_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNITEUV5_5_LC_6_11_4 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \POWERLED.dutycycle_RNITEUV5_5_LC_6_11_4  (
            .in0(N__15350),
            .in1(_gnd_net_),
            .in2(N__13532),
            .in3(N__15010),
            .lcout(\POWERLED.count_clk_1_sqmuxa_5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI9HME_1_LC_6_11_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI9HME_1_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI9HME_1_LC_6_11_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.func_state_RNI9HME_1_LC_6_11_5  (
            .in0(_gnd_net_),
            .in1(N__15212),
            .in2(_gnd_net_),
            .in3(N__15258),
            .lcout(\POWERLED.N_88 ),
            .ltout(\POWERLED.N_88_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIIA93A_0_LC_6_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIIA93A_0_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIIA93A_0_LC_6_11_6 .LUT_INIT=16'b1110111111001100;
    LogicCell40 \POWERLED.func_state_RNIIA93A_0_LC_6_11_6  (
            .in0(N__15137),
            .in1(N__13517),
            .in2(N__13496),
            .in3(N__15011),
            .lcout(\POWERLED.count_clk_1_sqmuxa_5_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI0AN05_0_LC_6_11_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI0AN05_0_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI0AN05_0_LC_6_11_7 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \POWERLED.func_state_RNI0AN05_0_LC_6_11_7  (
            .in0(N__14305),
            .in1(N__15216),
            .in2(N__13699),
            .in3(N__15998),
            .lcout(\POWERLED.N_250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_1_sqmuxa_5_0_a2_LC_6_12_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_1_sqmuxa_5_0_a2_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_1_sqmuxa_5_0_a2_LC_6_12_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.count_clk_1_sqmuxa_5_0_a2_LC_6_12_0  (
            .in0(N__15002),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15355),
            .lcout(\POWERLED.N_228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_1_0_LC_6_12_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_1_0_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_1_0_LC_6_12_1 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \POWERLED.func_state_RNO_1_0_LC_6_12_1  (
            .in0(N__15356),
            .in1(N__15211),
            .in2(N__15161),
            .in3(N__15003),
            .lcout(\POWERLED.N_179 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_3_1_LC_6_12_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_3_1_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_3_1_LC_6_12_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \POWERLED.func_state_RNO_3_1_LC_6_12_2  (
            .in0(N__15091),
            .in1(N__15104),
            .in2(N__16591),
            .in3(N__15645),
            .lcout(),
            .ltout(\POWERLED.N_208_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_1_1_LC_6_12_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_1_1_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_1_1_LC_6_12_3 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \POWERLED.func_state_RNO_1_1_LC_6_12_3  (
            .in0(N__13655),
            .in1(N__16583),
            .in2(N__13715),
            .in3(N__14897),
            .lcout(\POWERLED.func_state_ns_i_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_ns_0_i_0_0_a2_0_0_LC_6_12_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_ns_0_i_0_0_a2_0_0_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_ns_0_i_0_0_a2_0_0_LC_6_12_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \POWERLED.func_state_ns_0_i_0_0_a2_0_0_LC_6_12_4  (
            .in0(N__15092),
            .in1(N__15357),
            .in2(_gnd_net_),
            .in3(N__20708),
            .lcout(\POWERLED.N_222 ),
            .ltout(\POWERLED.N_222_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_2_1_LC_6_12_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_2_1_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_2_1_LC_6_12_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \POWERLED.func_state_RNO_2_1_LC_6_12_5  (
            .in0(N__15294),
            .in1(N__15210),
            .in2(N__13658),
            .in3(N__15148),
            .lcout(),
            .ltout(\POWERLED.N_211_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_0_1_LC_6_12_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_0_1_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_0_1_LC_6_12_6 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \POWERLED.func_state_RNO_0_1_LC_6_12_6  (
            .in0(_gnd_net_),
            .in1(N__13654),
            .in2(N__13646),
            .in3(N__15374),
            .lcout(\POWERLED.func_state_ns_i_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_0_0_LC_6_12_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_0_0_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_0_0_LC_6_12_7 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \POWERLED.func_state_RNO_0_0_LC_6_12_7  (
            .in0(N__15646),
            .in1(N__15090),
            .in2(N__14902),
            .in3(N__16582),
            .lcout(\POWERLED.N_178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_LC_6_13_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_LC_6_13_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_0_LC_6_13_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.func_state_0_LC_6_13_5  (
            .in0(N__13634),
            .in1(N__13628),
            .in2(N__13622),
            .in3(N__13610),
            .lcout(\POWERLED.func_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20534),
            .ce(N__19806),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_6_14_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_14_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_14_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_1_LC_6_15_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_1_LC_6_15_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_1_LC_6_15_3 .LUT_INIT=16'b0000111100100010;
    LogicCell40 \VPP_VDDQ.curr_state_1_LC_6_15_3  (
            .in0(N__15512),
            .in1(N__15584),
            .in2(N__18881),
            .in3(N__15542),
            .lcout(\VPP_VDDQ.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20593),
            .ce(N__19811),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_0_LC_6_15_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_0_LC_6_15_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_0_LC_6_15_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \VPP_VDDQ.curr_state_0_LC_6_15_5  (
            .in0(_gnd_net_),
            .in1(N__15541),
            .in2(_gnd_net_),
            .in3(N__15583),
            .lcout(\VPP_VDDQ.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20593),
            .ce(N__19811),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIH91A_0_LC_7_1_4 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIH91A_0_LC_7_1_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIH91A_0_LC_7_1_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \HDA_STRAP.curr_state_RNIH91A_0_LC_7_1_4  (
            .in0(_gnd_net_),
            .in1(N__15879),
            .in2(_gnd_net_),
            .in3(N__15809),
            .lcout(\HDA_STRAP.curr_state_RNIH91AZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIQC821_0_LC_7_1_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIQC821_0_LC_7_1_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIQC821_0_LC_7_1_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \HDA_STRAP.count_RNIQC821_0_LC_7_1_7  (
            .in0(N__13912),
            .in1(N__13900),
            .in2(N__13889),
            .in3(N__13873),
            .lcout(\HDA_STRAP.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_7_2_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_7_2_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \HDA_STRAP.count_RNIDLB61_6_LC_7_2_1  (
            .in0(N__13858),
            .in1(N__13957),
            .in2(N__13847),
            .in3(N__15679),
            .lcout(),
            .ltout(\HDA_STRAP.un4_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIUKIR1_12_LC_7_2_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIUKIR1_12_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIUKIR1_12_LC_7_2_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \HDA_STRAP.count_RNIUKIR1_12_LC_7_2_2  (
            .in0(N__13831),
            .in1(_gnd_net_),
            .in2(N__13820),
            .in3(N__13816),
            .lcout(\HDA_STRAP.un4_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNID0921_4_LC_7_2_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNID0921_4_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNID0921_4_LC_7_2_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \HDA_STRAP.count_RNID0921_4_LC_7_2_3  (
            .in0(N__13804),
            .in1(N__13792),
            .in2(N__13781),
            .in3(N__13765),
            .lcout(\HDA_STRAP.un4_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI63EA1_17_LC_7_2_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI63EA1_17_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI63EA1_17_LC_7_2_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \HDA_STRAP.count_RNI63EA1_17_LC_7_2_4  (
            .in0(N__13993),
            .in1(N__13754),
            .in2(N__14015),
            .in3(N__13975),
            .lcout(),
            .ltout(\HDA_STRAP.un4_count_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIB5IA5_0_LC_7_2_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIB5IA5_0_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIB5IA5_0_LC_7_2_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \HDA_STRAP.count_RNIB5IA5_0_LC_7_2_5  (
            .in0(N__13739),
            .in1(N__13733),
            .in2(N__13727),
            .in3(N__13724),
            .lcout(\HDA_STRAP.count_RNIB5IA5Z0Z_0 ),
            .ltout(\HDA_STRAP.count_RNIB5IA5Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_7_2_6 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_7_2_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \HDA_STRAP.curr_state_RNO_0_2_LC_7_2_6  (
            .in0(N__15902),
            .in1(_gnd_net_),
            .in2(N__13718),
            .in3(N__15810),
            .lcout(\HDA_STRAP.curr_state_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_10_LC_7_3_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_10_LC_7_3_0 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_10_LC_7_3_0 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \HDA_STRAP.count_10_LC_7_3_0  (
            .in0(N__15811),
            .in1(N__15904),
            .in2(N__14024),
            .in3(N__15723),
            .lcout(\HDA_STRAP.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20341),
            .ce(N__19762),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_16_LC_7_3_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_16_LC_7_3_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_16_LC_7_3_1 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \HDA_STRAP.count_16_LC_7_3_1  (
            .in0(N__15722),
            .in1(N__14000),
            .in2(N__15915),
            .in3(N__15814),
            .lcout(\HDA_STRAP.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20341),
            .ce(N__19762),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_17_LC_7_3_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_17_LC_7_3_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_17_LC_7_3_2 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \HDA_STRAP.count_17_LC_7_3_2  (
            .in0(N__15812),
            .in1(N__13982),
            .in2(N__15916),
            .in3(N__15724),
            .lcout(\HDA_STRAP.countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20341),
            .ce(N__19762),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_8_LC_7_3_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_8_LC_7_3_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_8_LC_7_3_6 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \HDA_STRAP.count_8_LC_7_3_6  (
            .in0(N__15813),
            .in1(N__13964),
            .in2(N__15917),
            .in3(N__15725),
            .lcout(\HDA_STRAP.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20341),
            .ce(N__19762),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI8M7Q_2_LC_7_5_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI8M7Q_2_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI8M7Q_2_LC_7_5_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \POWERLED.dutycycle_RNI8M7Q_2_LC_7_5_1  (
            .in0(N__14726),
            .in1(N__14602),
            .in2(N__14665),
            .in3(N__14394),
            .lcout(\POWERLED.un2_slp_s3n_2_0_o2_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI31MG_0_12_LC_7_5_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI31MG_0_12_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI31MG_0_12_LC_7_5_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI31MG_0_12_LC_7_5_2  (
            .in0(_gnd_net_),
            .in1(N__16467),
            .in2(_gnd_net_),
            .in3(N__16398),
            .lcout(\POWERLED.dutycycle_RNI31MG_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI31MG_12_LC_7_5_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI31MG_12_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI31MG_12_LC_7_5_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \POWERLED.dutycycle_RNI31MG_12_LC_7_5_3  (
            .in0(N__16468),
            .in1(_gnd_net_),
            .in2(N__16403),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI31MGZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIO2TE_9_LC_7_5_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIO2TE_9_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIO2TE_9_LC_7_5_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNIO2TE_9_LC_7_5_4  (
            .in0(_gnd_net_),
            .in1(N__16243),
            .in2(_gnd_net_),
            .in3(N__16397),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_1_39_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI34C41_8_LC_7_5_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI34C41_8_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI34C41_8_LC_7_5_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI34C41_8_LC_7_5_5  (
            .in0(N__16186),
            .in1(N__14395),
            .in2(N__14318),
            .in3(N__16080),
            .lcout(\POWERLED.dutycycle_RNI34C41Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI4I7Q_5_LC_7_6_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI4I7Q_5_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI4I7Q_5_LC_7_6_0 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \POWERLED.dutycycle_RNI4I7Q_5_LC_7_6_0  (
            .in0(N__14119),
            .in1(N__14195),
            .in2(N__14543),
            .in3(N__14455),
            .lcout(\POWERLED.N_117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIK4I81_6_LC_7_6_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIK4I81_6_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIK4I81_6_LC_7_6_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNIK4I81_6_LC_7_6_2  (
            .in0(N__14645),
            .in1(N__14279),
            .in2(N__14740),
            .in3(N__14454),
            .lcout(\POWERLED.dutycycle_RNIK4I81Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_2_LC_7_6_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_2_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_2_LC_7_6_3 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \POWERLED.dutycycle_2_LC_7_6_3  (
            .in0(N__14675),
            .in1(N__16761),
            .in2(N__14255),
            .in3(N__20716),
            .lcout(\POWERLED.dutycycleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20384),
            .ce(N__19749),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQAI81_4_LC_7_6_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQAI81_4_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQAI81_4_LC_7_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNIQAI81_4_LC_7_6_5  (
            .in0(N__14239),
            .in1(N__14585),
            .in2(N__14399),
            .in3(N__14646),
            .lcout(\POWERLED.dutycycle_RNIQAI81Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOQLJ_4_LC_7_6_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOQLJ_4_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOQLJ_4_LC_7_6_6 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \POWERLED.dutycycle_RNIOQLJ_4_LC_7_6_6  (
            .in0(N__14586),
            .in1(N__14392),
            .in2(_gnd_net_),
            .in3(N__14647),
            .lcout(\POWERLED.dutycycle_RNIOQLJZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_7_7_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_7_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__15388),
            .in2(N__15392),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\POWERLED.dutycycle_cry_c_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_0_0_LC_7_7_1 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNO_0_0_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_0_0_LC_7_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNO_0_0_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__14836),
            .in2(N__14213),
            .in3(N__14132),
            .lcout(\POWERLED.dutycycle_s_0 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_c_0_THRU_CO ),
            .carryout(\POWERLED.dutycycle_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_0_1_LC_7_7_2 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNO_0_1_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_0_1_LC_7_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNO_0_1_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__14128),
            .in2(N__14853),
            .in3(N__14039),
            .lcout(\POWERLED.dutycycle_s_1 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_0 ),
            .carryout(\POWERLED.dutycycle_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_1_2_LC_7_7_3 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNO_1_2_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_1_2_LC_7_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNO_1_2_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__14840),
            .in2(N__14741),
            .in3(N__14669),
            .lcout(\POWERLED.dutycycle_s_2 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_1 ),
            .carryout(\POWERLED.dutycycle_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_3_LC_7_7_4 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_3_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_3_LC_7_7_4 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_3_LC_7_7_4  (
            .in0(N__16772),
            .in1(N__14654),
            .in2(N__14854),
            .in3(N__14609),
            .lcout(\POWERLED.dutycycleZ0Z_3 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_2 ),
            .carryout(\POWERLED.dutycycle_cry_3 ),
            .clk(N__20450),
            .ce(N__19786),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_4_LC_7_7_5 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_4_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_4_LC_7_7_5 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_4_LC_7_7_5  (
            .in0(N__16760),
            .in1(N__14844),
            .in2(N__14603),
            .in3(N__14546),
            .lcout(\POWERLED.dutycycleZ0Z_4 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_3 ),
            .carryout(\POWERLED.dutycycle_cry_4 ),
            .clk(N__20450),
            .ce(N__19786),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_cry_c_RNIV95M9_4_LC_7_7_6 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_cry_c_RNIV95M9_4_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_cry_c_RNIV95M9_4_LC_7_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_cry_c_RNIV95M9_4_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__14542),
            .in2(N__14855),
            .in3(N__14462),
            .lcout(\POWERLED.dutycycle_s_5 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_4 ),
            .carryout(\POWERLED.dutycycle_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_cry_c_RNI1C5M9_5_LC_7_7_7 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_cry_c_RNI1C5M9_5_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_cry_c_RNI1C5M9_5_LC_7_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_cry_c_RNI1C5M9_5_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(N__14848),
            .in2(N__14459),
            .in3(N__14402),
            .lcout(\POWERLED.dutycycle_s_6 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_5 ),
            .carryout(\POWERLED.dutycycle_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_7_LC_7_8_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_7_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_7_LC_7_8_0 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_7_LC_7_8_0  (
            .in0(N__16758),
            .in1(N__14820),
            .in2(N__14396),
            .in3(N__14327),
            .lcout(\POWERLED.dutycycleZ0Z_7 ),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(\POWERLED.dutycycle_cry_7 ),
            .clk(N__20473),
            .ce(N__19774),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_8_LC_7_8_1 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_8_LC_7_8_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_8_LC_7_8_1 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_8_LC_7_8_1  (
            .in0(N__16738),
            .in1(N__16073),
            .in2(N__14849),
            .in3(N__14324),
            .lcout(\POWERLED.dutycycleZ0Z_8 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_7 ),
            .carryout(\POWERLED.dutycycle_cry_8 ),
            .clk(N__20473),
            .ce(N__19774),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_9_LC_7_8_2 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_9_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_9_LC_7_8_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_9_LC_7_8_2  (
            .in0(N__16759),
            .in1(N__14824),
            .in2(N__16244),
            .in3(N__14321),
            .lcout(\POWERLED.dutycycleZ0Z_9 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_8 ),
            .carryout(\POWERLED.dutycycle_cry_9 ),
            .clk(N__20473),
            .ce(N__19774),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_10_LC_7_8_3 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_10_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_10_LC_7_8_3 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_10_LC_7_8_3  (
            .in0(N__16735),
            .in1(N__16287),
            .in2(N__14850),
            .in3(N__14870),
            .lcout(\POWERLED.dutycycleZ0Z_10 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_9 ),
            .carryout(\POWERLED.dutycycle_cry_10 ),
            .clk(N__20473),
            .ce(N__19774),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_11_LC_7_8_4 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_11_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_11_LC_7_8_4 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_11_LC_7_8_4  (
            .in0(N__16756),
            .in1(N__14828),
            .in2(N__16187),
            .in3(N__14867),
            .lcout(\POWERLED.dutycycleZ0Z_11 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_10 ),
            .carryout(\POWERLED.dutycycle_cry_11 ),
            .clk(N__20473),
            .ce(N__19774),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_12_LC_7_8_5 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_12_LC_7_8_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_12_LC_7_8_5 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_12_LC_7_8_5  (
            .in0(N__16736),
            .in1(N__16396),
            .in2(N__14851),
            .in3(N__14864),
            .lcout(\POWERLED.dutycycleZ0Z_12 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_11 ),
            .carryout(\POWERLED.dutycycle_cry_12 ),
            .clk(N__20473),
            .ce(N__19774),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_13_LC_7_8_6 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_13_LC_7_8_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_13_LC_7_8_6 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_13_LC_7_8_6  (
            .in0(N__16757),
            .in1(N__14832),
            .in2(N__16469),
            .in3(N__14861),
            .lcout(\POWERLED.dutycycleZ0Z_13 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_12 ),
            .carryout(\POWERLED.dutycycle_cry_13 ),
            .clk(N__20473),
            .ce(N__19774),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_14_LC_7_8_7 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_14_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_14_LC_7_8_7 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_14_LC_7_8_7  (
            .in0(N__16737),
            .in1(N__16343),
            .in2(N__14852),
            .in3(N__14858),
            .lcout(\POWERLED.dutycycleZ0Z_14 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_13 ),
            .carryout(\POWERLED.dutycycle_cry_14 ),
            .clk(N__20473),
            .ce(N__19774),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_15_LC_7_9_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_15_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_15_LC_7_9_0 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_15_LC_7_9_0  (
            .in0(N__16739),
            .in1(N__14804),
            .in2(N__16130),
            .in3(N__14768),
            .lcout(\POWERLED.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20451),
            .ce(N__19785),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI33DK1_1_LC_7_10_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI33DK1_1_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI33DK1_1_LC_7_10_0 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \POWERLED.func_state_RNI33DK1_1_LC_7_10_0  (
            .in0(N__15299),
            .in1(N__15222),
            .in2(N__15097),
            .in3(N__15648),
            .lcout(\POWERLED.N_246 ),
            .ltout(\POWERLED.N_246_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIS9OC3_1_LC_7_10_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIS9OC3_1_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIS9OC3_1_LC_7_10_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \POWERLED.func_state_RNIS9OC3_1_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14765),
            .in3(N__16645),
            .lcout(\POWERLED.N_203_4 ),
            .ltout(\POWERLED.N_203_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI09QT9_1_LC_7_10_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI09QT9_1_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI09QT9_1_LC_7_10_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \POWERLED.count_clk_RNI09QT9_1_LC_7_10_2  (
            .in0(N__16607),
            .in1(N__16825),
            .in2(N__14756),
            .in3(N__15162),
            .lcout(),
            .ltout(\POWERLED.N_203_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNITU0DB_1_LC_7_10_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNITU0DB_1_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNITU0DB_1_LC_7_10_3 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \POWERLED.count_clk_RNITU0DB_1_LC_7_10_3  (
            .in0(N__15650),
            .in1(N__15086),
            .in2(N__14960),
            .in3(N__16556),
            .lcout(\POWERLED.count_clk_139_tz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI2M0Q4_6_LC_7_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI2M0Q4_6_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI2M0Q4_6_LC_7_10_4 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \POWERLED.count_clk_RNI2M0Q4_6_LC_7_10_4  (
            .in0(N__18056),
            .in1(N__15649),
            .in2(N__16672),
            .in3(N__16623),
            .lcout(\POWERLED.N_251 ),
            .ltout(\POWERLED.N_251_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI01TCL_7_LC_7_10_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI01TCL_7_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI01TCL_7_LC_7_10_5 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \POWERLED.count_clk_RNI01TCL_7_LC_7_10_5  (
            .in0(N__18020),
            .in1(N__14912),
            .in2(N__14957),
            .in3(N__14954),
            .lcout(),
            .ltout(\POWERLED.un2_slp_s3n_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIOH1J11_7_LC_7_10_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIOH1J11_7_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIOH1J11_7_LC_7_10_6 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \POWERLED.count_clk_RNIOH1J11_7_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(N__14948),
            .in2(N__14942),
            .in3(N__20056),
            .lcout(\POWERLED.count_clk_RNIOH1J11Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIORSP5_1_LC_7_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIORSP5_1_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIORSP5_1_LC_7_10_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.func_state_RNIORSP5_1_LC_7_10_7  (
            .in0(N__15163),
            .in1(N__16557),
            .in2(_gnd_net_),
            .in3(N__14939),
            .lcout(\POWERLED.N_205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIA8VP_7_LC_7_11_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIA8VP_7_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIA8VP_7_LC_7_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_clk_RNIA8VP_7_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__18016),
            .in2(_gnd_net_),
            .in3(N__15372),
            .lcout(),
            .ltout(\POWERLED.un2_slp_s3n_2_0_a6_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIAIGJ4_7_LC_7_11_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIAIGJ4_7_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIAIGJ4_7_LC_7_11_1 .LUT_INIT=16'b1011101110111010;
    LogicCell40 \POWERLED.count_clk_RNIAIGJ4_7_LC_7_11_1  (
            .in0(N__15012),
            .in1(N__15643),
            .in2(N__14915),
            .in3(N__16629),
            .lcout(\POWERLED.un2_slp_s3n_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI7LE01_7_LC_7_11_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI7LE01_7_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI7LE01_7_LC_7_11_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \POWERLED.count_clk_RNI7LE01_7_LC_7_11_2  (
            .in0(N__15083),
            .in1(N__18017),
            .in2(_gnd_net_),
            .in3(N__15221),
            .lcout(\POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNINTA34_1_LC_7_11_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNINTA34_1_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNINTA34_1_LC_7_11_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \POWERLED.func_state_RNINTA34_1_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__15301),
            .in2(_gnd_net_),
            .in3(N__15157),
            .lcout(\POWERLED.N_127 ),
            .ltout(\POWERLED.N_127_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIUIEUK_1_LC_7_11_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIUIEUK_1_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIUIEUK_1_LC_7_11_4 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \POWERLED.func_state_RNIUIEUK_1_LC_7_11_4  (
            .in0(N__15644),
            .in1(N__15461),
            .in2(N__15455),
            .in3(N__15452),
            .lcout(\POWERLED.count_clk_1_sqmuxa_5_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIH2SJ1_1_LC_7_11_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIH2SJ1_1_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIH2SJ1_1_LC_7_11_5 .LUT_INIT=16'b1001100100011001;
    LogicCell40 \POWERLED.func_state_RNIH2SJ1_1_LC_7_11_5  (
            .in0(N__15351),
            .in1(N__15085),
            .in2(N__16577),
            .in3(N__15438),
            .lcout(),
            .ltout(\POWERLED.dutycycle_3_sqmuxa_1_i_0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI6KL57_0_LC_7_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI6KL57_0_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI6KL57_0_LC_7_11_6 .LUT_INIT=16'b1111010111110100;
    LogicCell40 \POWERLED.func_state_RNI6KL57_0_LC_7_11_6  (
            .in0(N__15084),
            .in1(N__15373),
            .in2(N__15422),
            .in3(N__15418),
            .lcout(\POWERLED.N_366_1 ),
            .ltout(\POWERLED.N_366_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI446AD_7_LC_7_11_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI446AD_7_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI446AD_7_LC_7_11_7 .LUT_INIT=16'b1111101111110011;
    LogicCell40 \POWERLED.count_clk_RNI446AD_7_LC_7_11_7  (
            .in0(N__15407),
            .in1(N__20704),
            .in2(N__15401),
            .in3(N__15398),
            .lcout(\POWERLED.dutycycle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI9HME_0_1_LC_7_12_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI9HME_0_1_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI9HME_0_1_LC_7_12_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.func_state_RNI9HME_0_1_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__15289),
            .in2(_gnd_net_),
            .in3(N__15208),
            .lcout(\POWERLED.N_243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.N_55_i_i_o6_LC_7_12_2 .C_ON=1'b0;
    defparam \POWERLED.N_55_i_i_o6_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.N_55_i_i_o6_LC_7_12_2 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \POWERLED.N_55_i_i_o6_LC_7_12_2  (
            .in0(N__15358),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20702),
            .lcout(N_55),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_4_1_LC_7_12_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_4_1_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_4_1_LC_7_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.func_state_RNO_4_1_LC_7_12_4  (
            .in0(N__15293),
            .in1(N__15209),
            .in2(_gnd_net_),
            .in3(N__15164),
            .lcout(\POWERLED.N_148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_EN_i_i_0_a2_LC_7_13_0 .C_ON=1'b0;
    defparam \POWERLED.VCCST_EN_i_i_0_a2_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_EN_i_i_0_a2_LC_7_13_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.VCCST_EN_i_i_0_a2_LC_7_13_0  (
            .in0(N__20703),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15057),
            .lcout(vccst_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIJKKQ_LC_7_13_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIJKKQ_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIJKKQ_LC_7_13_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNIJKKQ_LC_7_13_4  (
            .in0(N__15647),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15554),
            .lcout(vpp_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_7_14_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_7_14_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_7_14_0  (
            .in0(N__15582),
            .in1(N__15508),
            .in2(_gnd_net_),
            .in3(N__15540),
            .lcout(\VPP_VDDQ.G_127_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNIDNTT1_0_LC_7_14_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNIDNTT1_0_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNIDNTT1_0_LC_7_14_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \VPP_VDDQ.curr_state_RNIDNTT1_0_LC_7_14_1  (
            .in0(N__15507),
            .in1(N__15538),
            .in2(_gnd_net_),
            .in3(N__15581),
            .lcout(\VPP_VDDQ.N_108_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_LC_7_14_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_LC_7_14_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_LC_7_14_2  (
            .in0(N__19555),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15652),
            .lcout(\VPP_VDDQ.N_238 ),
            .ltout(\VPP_VDDQ.N_238_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNINMKE1_1_LC_7_14_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNINMKE1_1_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNINMKE1_1_LC_7_14_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \VPP_VDDQ.curr_state_RNINMKE1_1_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15566),
            .in3(N__15537),
            .lcout(\VPP_VDDQ.N_128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_7_14_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_7_14_6 .LUT_INIT=16'b0011100010101010;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_7_14_6  (
            .in0(N__15553),
            .in1(N__15509),
            .in2(N__15482),
            .in3(N__20083),
            .lcout(),
            .ltout(\VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_7_14_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_7_14_7 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_LC_7_14_7  (
            .in0(N__20084),
            .in1(_gnd_net_),
            .in2(N__15563),
            .in3(N__15560),
            .lcout(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20547),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNI8I855_0_LC_7_15_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNI8I855_0_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNI8I855_0_LC_7_15_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.curr_state_RNI8I855_0_LC_7_15_0  (
            .in0(N__15510),
            .in1(N__15539),
            .in2(_gnd_net_),
            .in3(N__18877),
            .lcout(),
            .ltout(\VPP_VDDQ.N_154_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNIGR9S7_0_LC_7_15_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNIGR9S7_0_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNIGR9S7_0_LC_7_15_1 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \VPP_VDDQ.curr_state_RNIGR9S7_0_LC_7_15_1  (
            .in0(N__15511),
            .in1(N__15475),
            .in2(N__15464),
            .in3(N__20062),
            .lcout(\VPP_VDDQ.curr_state_RNIGR9S7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_7_16_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_7_16_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \VPP_VDDQ.count_esr_RNO_0_15_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__16923),
            .in2(_gnd_net_),
            .in3(N__20078),
            .lcout(\VPP_VDDQ.N_65_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_6_LC_8_1_2 .C_ON=1'b0;
    defparam \COUNTER.counter_6_LC_8_1_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_6_LC_8_1_2 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \COUNTER.counter_6_LC_8_1_2  (
            .in0(N__19444),
            .in1(_gnd_net_),
            .in2(N__17027),
            .in3(N__17009),
            .lcout(\COUNTER.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20206),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_5_LC_8_1_3 .C_ON=1'b0;
    defparam \COUNTER.counter_5_LC_8_1_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_5_LC_8_1_3 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_5_LC_8_1_3  (
            .in0(N__17050),
            .in1(N__17036),
            .in2(_gnd_net_),
            .in3(N__19443),
            .lcout(\COUNTER.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20206),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_LC_8_1_4 .C_ON=1'b0;
    defparam \COUNTER.counter_1_LC_8_1_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_1_LC_8_1_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \COUNTER.counter_1_LC_8_1_4  (
            .in0(N__19445),
            .in1(N__16909),
            .in2(_gnd_net_),
            .in3(N__17591),
            .lcout(\COUNTER.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20206),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_RNO_LC_8_1_6 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_8_1_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \COUNTER.un4_counter_1_c_RNO_LC_8_1_6  (
            .in0(N__17022),
            .in1(N__17049),
            .in2(N__17000),
            .in3(N__16908),
            .lcout(\COUNTER.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_6_LC_8_2_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_6_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_6_LC_8_2_1 .LUT_INIT=16'b1000101010101010;
    LogicCell40 \HDA_STRAP.count_6_LC_8_2_1  (
            .in0(N__15929),
            .in1(N__15903),
            .in2(N__15818),
            .in3(N__15721),
            .lcout(\HDA_STRAP.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20377),
            .ce(N__19742),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_0_LC_8_5_0 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_0_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_0_LC_8_5_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_0_LC_8_5_0  (
            .in0(N__20118),
            .in1(N__17345),
            .in2(N__19384),
            .in3(N__19385),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_5_0_),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_0 ),
            .clk(N__20533),
            .ce(),
            .sr(N__17891));
    defparam \ALL_SYS_PWRGD.count_1_LC_8_5_1 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_1_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_1_LC_8_5_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_1_LC_8_5_1  (
            .in0(N__20103),
            .in1(N__17384),
            .in2(_gnd_net_),
            .in3(N__15668),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_0 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_1 ),
            .clk(N__20533),
            .ce(),
            .sr(N__17891));
    defparam \ALL_SYS_PWRGD.count_2_LC_8_5_2 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_2_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_2_LC_8_5_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_2_LC_8_5_2  (
            .in0(N__20119),
            .in1(N__17231),
            .in2(_gnd_net_),
            .in3(N__15665),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_1 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_2 ),
            .clk(N__20533),
            .ce(),
            .sr(N__17891));
    defparam \ALL_SYS_PWRGD.count_3_LC_8_5_3 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_3_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_3_LC_8_5_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_3_LC_8_5_3  (
            .in0(N__20104),
            .in1(N__17258),
            .in2(_gnd_net_),
            .in3(N__15662),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_2 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_3 ),
            .clk(N__20533),
            .ce(),
            .sr(N__17891));
    defparam \ALL_SYS_PWRGD.count_4_LC_8_5_4 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_4_LC_8_5_4 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_4_LC_8_5_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_4_LC_8_5_4  (
            .in0(N__20120),
            .in1(N__17462),
            .in2(_gnd_net_),
            .in3(N__15956),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_3 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_4 ),
            .clk(N__20533),
            .ce(),
            .sr(N__17891));
    defparam \ALL_SYS_PWRGD.count_5_LC_8_5_5 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_5_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_5_LC_8_5_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_5_LC_8_5_5  (
            .in0(N__20105),
            .in1(N__17270),
            .in2(_gnd_net_),
            .in3(N__15953),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_4 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_5 ),
            .clk(N__20533),
            .ce(),
            .sr(N__17891));
    defparam \ALL_SYS_PWRGD.count_6_LC_8_5_6 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_6_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_6_LC_8_5_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_6_LC_8_5_6  (
            .in0(N__20121),
            .in1(N__17476),
            .in2(_gnd_net_),
            .in3(N__15950),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_5 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_6 ),
            .clk(N__20533),
            .ce(),
            .sr(N__17891));
    defparam \ALL_SYS_PWRGD.count_7_LC_8_5_7 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_7_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_7_LC_8_5_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_7_LC_8_5_7  (
            .in0(N__20106),
            .in1(N__17501),
            .in2(_gnd_net_),
            .in3(N__15947),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_6 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_7 ),
            .clk(N__20533),
            .ce(),
            .sr(N__17891));
    defparam \ALL_SYS_PWRGD.count_8_LC_8_6_0 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_8_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_8_LC_8_6_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_8_LC_8_6_0  (
            .in0(N__20082),
            .in1(N__17489),
            .in2(_gnd_net_),
            .in3(N__15944),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_8 ),
            .clk(N__20472),
            .ce(),
            .sr(N__17890));
    defparam \ALL_SYS_PWRGD.count_9_LC_8_6_1 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_9_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_9_LC_8_6_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_9_LC_8_6_1  (
            .in0(N__20073),
            .in1(N__17372),
            .in2(_gnd_net_),
            .in3(N__15941),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_8 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_9 ),
            .clk(N__20472),
            .ce(),
            .sr(N__17890));
    defparam \ALL_SYS_PWRGD.count_10_LC_8_6_2 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_10_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_10_LC_8_6_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_10_LC_8_6_2  (
            .in0(N__20079),
            .in1(N__17359),
            .in2(_gnd_net_),
            .in3(N__15938),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_9 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_10 ),
            .clk(N__20472),
            .ce(),
            .sr(N__17890));
    defparam \ALL_SYS_PWRGD.count_11_LC_8_6_3 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_11_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_11_LC_8_6_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_11_LC_8_6_3  (
            .in0(N__20071),
            .in1(N__17245),
            .in2(_gnd_net_),
            .in3(N__15935),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_10 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_11 ),
            .clk(N__20472),
            .ce(),
            .sr(N__17890));
    defparam \ALL_SYS_PWRGD.count_12_LC_8_6_4 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_12_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_12_LC_8_6_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_12_LC_8_6_4  (
            .in0(N__20080),
            .in1(N__17411),
            .in2(_gnd_net_),
            .in3(N__15932),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_11 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_12 ),
            .clk(N__20472),
            .ce(),
            .sr(N__17890));
    defparam \ALL_SYS_PWRGD.count_13_LC_8_6_5 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_13_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_13_LC_8_6_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_13_LC_8_6_5  (
            .in0(N__20072),
            .in1(N__17425),
            .in2(_gnd_net_),
            .in3(N__16502),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_12 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_13 ),
            .clk(N__20472),
            .ce(),
            .sr(N__17890));
    defparam \ALL_SYS_PWRGD.count_14_LC_8_6_6 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_14_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_14_LC_8_6_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_14_LC_8_6_6  (
            .in0(N__20081),
            .in1(N__17450),
            .in2(_gnd_net_),
            .in3(N__16499),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_13 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_14 ),
            .clk(N__20472),
            .ce(),
            .sr(N__17890));
    defparam \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_6_7 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_6_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(N__18375),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_14 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_esr_15_LC_8_7_0 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_esr_15_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_esr_15_LC_8_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALL_SYS_PWRGD.count_esr_15_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__17438),
            .in2(_gnd_net_),
            .in3(N__16496),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20557),
            .ce(N__17858),
            .sr(N__17883));
    defparam \POWERLED.dutycycle_RNIO18N_9_LC_8_8_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIO18N_9_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIO18N_9_LC_8_8_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \POWERLED.dutycycle_RNIO18N_9_LC_8_8_0  (
            .in0(N__16235),
            .in1(N__16452),
            .in2(_gnd_net_),
            .in3(N__16285),
            .lcout(\POWERLED.dutycycle_RNIO18NZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI51C11_10_LC_8_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI51C11_10_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI51C11_10_LC_8_8_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.dutycycle_RNI51C11_10_LC_8_8_2  (
            .in0(N__16461),
            .in1(N__16395),
            .in2(N__16346),
            .in3(N__16286),
            .lcout(\POWERLED.un2_slp_s3n_2_0_o2_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIH6QT_15_LC_8_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIH6QT_15_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIH6QT_15_LC_8_8_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.dutycycle_RNIH6QT_15_LC_8_8_5  (
            .in0(N__16238),
            .in1(N__16180),
            .in2(N__16129),
            .in3(N__16072),
            .lcout(),
            .ltout(\POWERLED.un2_slp_s3n_2_0_o2_3_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIUTDP2_2_LC_8_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIUTDP2_2_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIUTDP2_2_LC_8_8_6 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \POWERLED.dutycycle_RNIUTDP2_2_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__16022),
            .in2(N__16016),
            .in3(N__16013),
            .lcout(\POWERLED.N_112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIROMF7_0_LC_8_9_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIROMF7_0_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIROMF7_0_LC_8_9_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \POWERLED.func_state_RNIROMF7_0_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__16784),
            .in2(_gnd_net_),
            .in3(N__20715),
            .lcout(\POWERLED.un1_dutycycle_4_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIPG2D1_2_LC_8_9_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIPG2D1_2_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIPG2D1_2_LC_8_9_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.count_clk_RNIPG2D1_2_LC_8_9_2  (
            .in0(N__18097),
            .in1(N__18115),
            .in2(N__17648),
            .in3(N__17950),
            .lcout(\POWERLED.N_177_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIP4HM_2_LC_8_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIP4HM_2_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIP4HM_2_LC_8_9_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \POWERLED.count_clk_RNIP4HM_2_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__18114),
            .in2(_gnd_net_),
            .in3(N__17643),
            .lcout(),
            .ltout(\POWERLED.count_clk_0_sqmuxa_5_0_o2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIP6BO1_4_LC_8_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIP6BO1_4_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIP6BO1_4_LC_8_9_5 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \POWERLED.count_clk_RNIP6BO1_4_LC_8_9_5  (
            .in0(N__17949),
            .in1(N__18044),
            .in2(N__16655),
            .in3(N__18096),
            .lcout(\POWERLED.N_141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIKKV71_12_LC_8_10_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIKKV71_12_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIKKV71_12_LC_8_10_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNIKKV71_12_LC_8_10_0  (
            .in0(N__18442),
            .in1(N__17680),
            .in2(N__18428),
            .in3(N__16598),
            .lcout(\POWERLED.N_136 ),
            .ltout(\POWERLED.N_136_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIHJP92_1_LC_8_10_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIHJP92_1_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIHJP92_1_LC_8_10_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \POWERLED.count_clk_RNIHJP92_1_LC_8_10_1  (
            .in0(N__17930),
            .in1(N__18077),
            .in2(N__16634),
            .in3(N__17666),
            .lcout(\POWERLED.N_146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIUL2D1_1_LC_8_10_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIUL2D1_1_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIUL2D1_1_LC_8_10_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.count_clk_RNIUL2D1_1_LC_8_10_2  (
            .in0(N__17667),
            .in1(N__17931),
            .in2(N__18006),
            .in3(N__18078),
            .lcout(\POWERLED.count_clk_0_sqmuxa_5_0_a6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_esr_RNO_0_15_LC_8_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_esr_RNO_0_15_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_esr_RNO_0_15_LC_8_10_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.count_clk_esr_RNO_0_15_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__18233),
            .in2(_gnd_net_),
            .in3(N__20061),
            .lcout(\POWERLED.N_65_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_esr_RNIVU6L_15_LC_8_10_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_esr_RNIVU6L_15_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_esr_RNIVU6L_15_LC_8_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_esr_RNIVU6L_15_LC_8_10_5  (
            .in0(N__18409),
            .in1(N__18457),
            .in2(N__18281),
            .in3(N__17911),
            .lcout(\POWERLED.count_clk_0_sqmuxa_5_0_o2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI3G101_5_LC_8_10_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI3G101_5_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI3G101_5_LC_8_10_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.count_clk_RNI3G101_5_LC_8_10_6  (
            .in0(N__17990),
            .in1(N__16537),
            .in2(_gnd_net_),
            .in3(N__18079),
            .lcout(),
            .ltout(\POWERLED.count_off_1_sqmuxa_i_a6_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNILEIU2_1_LC_8_10_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNILEIU2_1_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNILEIU2_1_LC_8_10_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.count_clk_RNILEIU2_1_LC_8_10_7  (
            .in0(N__17932),
            .in1(N__17668),
            .in2(N__16829),
            .in3(N__16826),
            .lcout(\POWERLED.count_off_1_sqmuxa_i_a6_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_0_LC_8_11_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_0_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_0_LC_8_11_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_0_LC_8_11_0  (
            .in0(N__20142),
            .in1(N__18167),
            .in2(N__18491),
            .in3(N__18490),
            .lcout(\RSMRST_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .clk(N__20636),
            .ce(),
            .sr(N__18530));
    defparam \RSMRST_PWRGD.count_1_LC_8_11_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_1_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_1_LC_8_11_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_1_LC_8_11_1  (
            .in0(N__20132),
            .in1(N__18551),
            .in2(_gnd_net_),
            .in3(N__16805),
            .lcout(\RSMRST_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .clk(N__20636),
            .ce(),
            .sr(N__18530));
    defparam \RSMRST_PWRGD.count_2_LC_8_11_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_2_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_2_LC_8_11_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_2_LC_8_11_2  (
            .in0(N__20143),
            .in1(N__18578),
            .in2(_gnd_net_),
            .in3(N__16802),
            .lcout(\RSMRST_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .clk(N__20636),
            .ce(),
            .sr(N__18530));
    defparam \RSMRST_PWRGD.count_3_LC_8_11_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_3_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_3_LC_8_11_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_3_LC_8_11_3  (
            .in0(N__20133),
            .in1(N__18608),
            .in2(_gnd_net_),
            .in3(N__16799),
            .lcout(\RSMRST_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .clk(N__20636),
            .ce(),
            .sr(N__18530));
    defparam \RSMRST_PWRGD.count_4_LC_8_11_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_4_LC_8_11_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_4_LC_8_11_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_4_LC_8_11_4  (
            .in0(N__20144),
            .in1(N__18590),
            .in2(_gnd_net_),
            .in3(N__16796),
            .lcout(\RSMRST_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .clk(N__20636),
            .ce(),
            .sr(N__18530));
    defparam \RSMRST_PWRGD.count_5_LC_8_11_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_5_LC_8_11_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_5_LC_8_11_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_5_LC_8_11_5  (
            .in0(N__20134),
            .in1(N__18565),
            .in2(_gnd_net_),
            .in3(N__16793),
            .lcout(\RSMRST_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .clk(N__20636),
            .ce(),
            .sr(N__18530));
    defparam \RSMRST_PWRGD.count_6_LC_8_11_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_6_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_6_LC_8_11_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_6_LC_8_11_6  (
            .in0(N__20145),
            .in1(N__18179),
            .in2(_gnd_net_),
            .in3(N__16790),
            .lcout(\RSMRST_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .clk(N__20636),
            .ce(),
            .sr(N__18530));
    defparam \RSMRST_PWRGD.count_7_LC_8_11_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_7_LC_8_11_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_7_LC_8_11_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_7_LC_8_11_7  (
            .in0(N__20135),
            .in1(N__18623),
            .in2(_gnd_net_),
            .in3(N__16787),
            .lcout(\RSMRST_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .clk(N__20636),
            .ce(),
            .sr(N__18530));
    defparam \RSMRST_PWRGD.count_8_LC_8_12_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_8_LC_8_12_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_8_LC_8_12_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_8_LC_8_12_0  (
            .in0(N__20149),
            .in1(N__18155),
            .in2(_gnd_net_),
            .in3(N__16853),
            .lcout(\RSMRST_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .clk(N__20631),
            .ce(),
            .sr(N__18529));
    defparam \RSMRST_PWRGD.count_9_LC_8_12_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_9_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_9_LC_8_12_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_9_LC_8_12_1  (
            .in0(N__20138),
            .in1(N__18142),
            .in2(_gnd_net_),
            .in3(N__16850),
            .lcout(\RSMRST_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .clk(N__20631),
            .ce(),
            .sr(N__18529));
    defparam \RSMRST_PWRGD.count_10_LC_8_12_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_10_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_10_LC_8_12_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_10_LC_8_12_2  (
            .in0(N__20146),
            .in1(N__18206),
            .in2(_gnd_net_),
            .in3(N__16847),
            .lcout(\RSMRST_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .clk(N__20631),
            .ce(),
            .sr(N__18529));
    defparam \RSMRST_PWRGD.count_11_LC_8_12_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_11_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_11_LC_8_12_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_11_LC_8_12_3  (
            .in0(N__20136),
            .in1(N__18218),
            .in2(_gnd_net_),
            .in3(N__16844),
            .lcout(\RSMRST_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .clk(N__20631),
            .ce(),
            .sr(N__18529));
    defparam \RSMRST_PWRGD.count_12_LC_8_12_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_12_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_12_LC_8_12_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_12_LC_8_12_4  (
            .in0(N__20147),
            .in1(N__18128),
            .in2(_gnd_net_),
            .in3(N__16841),
            .lcout(\RSMRST_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .clk(N__20631),
            .ce(),
            .sr(N__18529));
    defparam \RSMRST_PWRGD.count_13_LC_8_12_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_13_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_13_LC_8_12_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_13_LC_8_12_5  (
            .in0(N__20137),
            .in1(N__18193),
            .in2(_gnd_net_),
            .in3(N__16838),
            .lcout(\RSMRST_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .clk(N__20631),
            .ce(),
            .sr(N__18529));
    defparam \RSMRST_PWRGD.count_14_LC_8_12_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_14_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_14_LC_8_12_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_14_LC_8_12_6  (
            .in0(N__20148),
            .in1(N__18635),
            .in2(_gnd_net_),
            .in3(N__16835),
            .lcout(\RSMRST_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .clk(N__20631),
            .ce(),
            .sr(N__18529));
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_12_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__18337),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_15_LC_8_13_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_15_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_esr_15_LC_8_13_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \RSMRST_PWRGD.count_esr_15_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__18647),
            .in2(_gnd_net_),
            .in3(N__16832),
            .lcout(\RSMRST_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20637),
            .ce(N__18497),
            .sr(N__18522));
    defparam \VPP_VDDQ.count_0_LC_8_14_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_0_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_0_LC_8_14_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_0_LC_8_14_0  (
            .in0(N__20128),
            .in1(N__18914),
            .in2(N__16894),
            .in3(N__16895),
            .lcout(\VPP_VDDQ.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_0 ),
            .clk(N__20600),
            .ce(),
            .sr(N__16942));
    defparam \VPP_VDDQ.count_1_LC_8_14_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_1_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_1_LC_8_14_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_1_LC_8_14_1  (
            .in0(N__20110),
            .in1(N__18968),
            .in2(_gnd_net_),
            .in3(N__16877),
            .lcout(\VPP_VDDQ.countZ0Z_1 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_0 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_1 ),
            .clk(N__20600),
            .ce(),
            .sr(N__16942));
    defparam \VPP_VDDQ.count_2_LC_8_14_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_2_LC_8_14_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_LC_8_14_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_2_LC_8_14_2  (
            .in0(N__20129),
            .in1(N__18995),
            .in2(_gnd_net_),
            .in3(N__16874),
            .lcout(\VPP_VDDQ.countZ0Z_2 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_2 ),
            .clk(N__20600),
            .ce(),
            .sr(N__16942));
    defparam \VPP_VDDQ.count_3_LC_8_14_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_3_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_3_LC_8_14_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_3_LC_8_14_3  (
            .in0(N__20111),
            .in1(N__19070),
            .in2(_gnd_net_),
            .in3(N__16871),
            .lcout(\VPP_VDDQ.countZ0Z_3 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_3 ),
            .clk(N__20600),
            .ce(),
            .sr(N__16942));
    defparam \VPP_VDDQ.count_4_LC_8_14_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_4_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_4_LC_8_14_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_4_LC_8_14_4  (
            .in0(N__20130),
            .in1(N__19097),
            .in2(_gnd_net_),
            .in3(N__16868),
            .lcout(\VPP_VDDQ.countZ0Z_4 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_4 ),
            .clk(N__20600),
            .ce(),
            .sr(N__16942));
    defparam \VPP_VDDQ.count_5_LC_8_14_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_5_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_5_LC_8_14_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_5_LC_8_14_5  (
            .in0(N__20112),
            .in1(N__18470),
            .in2(_gnd_net_),
            .in3(N__16865),
            .lcout(\VPP_VDDQ.countZ0Z_5 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_5 ),
            .clk(N__20600),
            .ce(),
            .sr(N__16942));
    defparam \VPP_VDDQ.count_6_LC_8_14_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_6_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_6_LC_8_14_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_6_LC_8_14_6  (
            .in0(N__20131),
            .in1(N__19007),
            .in2(_gnd_net_),
            .in3(N__16862),
            .lcout(\VPP_VDDQ.countZ0Z_6 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_6 ),
            .clk(N__20600),
            .ce(),
            .sr(N__16942));
    defparam \VPP_VDDQ.count_7_LC_8_14_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_7_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_7_LC_8_14_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_7_LC_8_14_7  (
            .in0(N__20113),
            .in1(N__19084),
            .in2(_gnd_net_),
            .in3(N__16859),
            .lcout(\VPP_VDDQ.countZ0Z_7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_7 ),
            .clk(N__20600),
            .ce(),
            .sr(N__16942));
    defparam \VPP_VDDQ.count_8_LC_8_15_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_8_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_8_LC_8_15_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_8_LC_8_15_0  (
            .in0(N__20159),
            .in1(N__18941),
            .in2(_gnd_net_),
            .in3(N__16856),
            .lcout(\VPP_VDDQ.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_8 ),
            .clk(N__20641),
            .ce(),
            .sr(N__16930));
    defparam \VPP_VDDQ.count_9_LC_8_15_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_9_LC_8_15_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_9_LC_8_15_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_9_LC_8_15_1  (
            .in0(N__20155),
            .in1(N__18955),
            .in2(_gnd_net_),
            .in3(N__16976),
            .lcout(\VPP_VDDQ.countZ0Z_9 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_8 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_9 ),
            .clk(N__20641),
            .ce(),
            .sr(N__16930));
    defparam \VPP_VDDQ.count_10_LC_8_15_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_10_LC_8_15_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_10_LC_8_15_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_10_LC_8_15_2  (
            .in0(N__20156),
            .in1(N__18982),
            .in2(_gnd_net_),
            .in3(N__16973),
            .lcout(\VPP_VDDQ.countZ0Z_10 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_10 ),
            .clk(N__20641),
            .ce(),
            .sr(N__16930));
    defparam \VPP_VDDQ.count_11_LC_8_15_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_11_LC_8_15_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_11_LC_8_15_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_11_LC_8_15_3  (
            .in0(N__20153),
            .in1(N__18928),
            .in2(_gnd_net_),
            .in3(N__16970),
            .lcout(\VPP_VDDQ.countZ0Z_11 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_11 ),
            .clk(N__20641),
            .ce(),
            .sr(N__16930));
    defparam \VPP_VDDQ.count_12_LC_8_15_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_12_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_12_LC_8_15_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_12_LC_8_15_4  (
            .in0(N__20157),
            .in1(N__19019),
            .in2(_gnd_net_),
            .in3(N__16967),
            .lcout(\VPP_VDDQ.countZ0Z_12 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_12 ),
            .clk(N__20641),
            .ce(),
            .sr(N__16930));
    defparam \VPP_VDDQ.count_13_LC_8_15_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_13_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_13_LC_8_15_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_13_LC_8_15_5  (
            .in0(N__20154),
            .in1(N__19033),
            .in2(_gnd_net_),
            .in3(N__16964),
            .lcout(\VPP_VDDQ.countZ0Z_13 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_13 ),
            .clk(N__20641),
            .ce(),
            .sr(N__16930));
    defparam \VPP_VDDQ.count_14_LC_8_15_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_14_LC_8_15_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_14_LC_8_15_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_14_LC_8_15_6  (
            .in0(N__20158),
            .in1(N__19058),
            .in2(_gnd_net_),
            .in3(N__16961),
            .lcout(\VPP_VDDQ.countZ0Z_14 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14 ),
            .clk(N__20641),
            .ce(),
            .sr(N__16930));
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_15_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(N__18336),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_14 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_15_LC_8_16_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_15_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_esr_15_LC_8_16_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \VPP_VDDQ.count_esr_15_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__19046),
            .in2(_gnd_net_),
            .in3(N__16958),
            .lcout(\VPP_VDDQ.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20642),
            .ce(N__16955),
            .sr(N__16946));
    defparam \COUNTER.counter_1_cry_1_c_LC_9_1_0 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_c_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_c_LC_9_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.counter_1_cry_1_c_LC_9_1_0  (
            .in0(_gnd_net_),
            .in1(N__16910),
            .in2(N__17590),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_1_0_),
            .carryout(\COUNTER.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_9_1_1 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_9_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_9_1_1  (
            .in0(_gnd_net_),
            .in1(N__17552),
            .in2(_gnd_net_),
            .in3(N__17060),
            .lcout(\COUNTER.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_1 ),
            .carryout(\COUNTER.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_9_1_2 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_9_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_9_1_2  (
            .in0(_gnd_net_),
            .in1(N__17522),
            .in2(_gnd_net_),
            .in3(N__17057),
            .lcout(\COUNTER.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_2 ),
            .carryout(\COUNTER.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_9_1_3 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_9_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_9_1_3  (
            .in0(_gnd_net_),
            .in1(N__17612),
            .in2(_gnd_net_),
            .in3(N__17054),
            .lcout(\COUNTER.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_3 ),
            .carryout(\COUNTER.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_9_1_4 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_9_1_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_9_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_9_1_4  (
            .in0(_gnd_net_),
            .in1(N__17051),
            .in2(_gnd_net_),
            .in3(N__17030),
            .lcout(\COUNTER.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_4 ),
            .carryout(\COUNTER.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_9_1_5 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_9_1_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_9_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_9_1_5  (
            .in0(_gnd_net_),
            .in1(N__17026),
            .in2(_gnd_net_),
            .in3(N__17003),
            .lcout(\COUNTER.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_5 ),
            .carryout(\COUNTER.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_7_LC_9_1_6 .C_ON=1'b1;
    defparam \COUNTER.counter_7_LC_9_1_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_7_LC_9_1_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_7_LC_9_1_6  (
            .in0(_gnd_net_),
            .in1(N__16999),
            .in2(_gnd_net_),
            .in3(N__16985),
            .lcout(\COUNTER.counterZ0Z_7 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_6 ),
            .carryout(\COUNTER.counter_1_cry_7 ),
            .clk(N__20407),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_8_LC_9_1_7 .C_ON=1'b1;
    defparam \COUNTER.counter_8_LC_9_1_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_8_LC_9_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_8_LC_9_1_7  (
            .in0(_gnd_net_),
            .in1(N__18670),
            .in2(_gnd_net_),
            .in3(N__16982),
            .lcout(\COUNTER.counterZ0Z_8 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_7 ),
            .carryout(\COUNTER.counter_1_cry_8 ),
            .clk(N__20407),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_9_LC_9_2_0 .C_ON=1'b1;
    defparam \COUNTER.counter_9_LC_9_2_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_9_LC_9_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_9_LC_9_2_0  (
            .in0(_gnd_net_),
            .in1(N__18709),
            .in2(_gnd_net_),
            .in3(N__16979),
            .lcout(\COUNTER.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_9_2_0_),
            .carryout(\COUNTER.counter_1_cry_9 ),
            .clk(N__20465),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_10_LC_9_2_1 .C_ON=1'b1;
    defparam \COUNTER.counter_10_LC_9_2_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_10_LC_9_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_10_LC_9_2_1  (
            .in0(_gnd_net_),
            .in1(N__18727),
            .in2(_gnd_net_),
            .in3(N__17087),
            .lcout(\COUNTER.counterZ0Z_10 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_9 ),
            .carryout(\COUNTER.counter_1_cry_10 ),
            .clk(N__20465),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_11_LC_9_2_2 .C_ON=1'b1;
    defparam \COUNTER.counter_11_LC_9_2_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_11_LC_9_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_11_LC_9_2_2  (
            .in0(_gnd_net_),
            .in1(N__18688),
            .in2(_gnd_net_),
            .in3(N__17084),
            .lcout(\COUNTER.counterZ0Z_11 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_10 ),
            .carryout(\COUNTER.counter_1_cry_11 ),
            .clk(N__20465),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_12_LC_9_2_3 .C_ON=1'b1;
    defparam \COUNTER.counter_12_LC_9_2_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_12_LC_9_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_12_LC_9_2_3  (
            .in0(_gnd_net_),
            .in1(N__18811),
            .in2(_gnd_net_),
            .in3(N__17081),
            .lcout(\COUNTER.counterZ0Z_12 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_11 ),
            .carryout(\COUNTER.counter_1_cry_12 ),
            .clk(N__20465),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_13_LC_9_2_4 .C_ON=1'b1;
    defparam \COUNTER.counter_13_LC_9_2_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_13_LC_9_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_13_LC_9_2_4  (
            .in0(_gnd_net_),
            .in1(N__18844),
            .in2(_gnd_net_),
            .in3(N__17078),
            .lcout(\COUNTER.counterZ0Z_13 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_12 ),
            .carryout(\COUNTER.counter_1_cry_13 ),
            .clk(N__20465),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_14_LC_9_2_5 .C_ON=1'b1;
    defparam \COUNTER.counter_14_LC_9_2_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_14_LC_9_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_14_LC_9_2_5  (
            .in0(_gnd_net_),
            .in1(N__18859),
            .in2(_gnd_net_),
            .in3(N__17075),
            .lcout(\COUNTER.counterZ0Z_14 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_13 ),
            .carryout(\COUNTER.counter_1_cry_14 ),
            .clk(N__20465),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_15_LC_9_2_6 .C_ON=1'b1;
    defparam \COUNTER.counter_15_LC_9_2_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_15_LC_9_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_15_LC_9_2_6  (
            .in0(_gnd_net_),
            .in1(N__18826),
            .in2(_gnd_net_),
            .in3(N__17072),
            .lcout(\COUNTER.counterZ0Z_15 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_14 ),
            .carryout(\COUNTER.counter_1_cry_15 ),
            .clk(N__20465),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_16_LC_9_2_7 .C_ON=1'b1;
    defparam \COUNTER.counter_16_LC_9_2_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_16_LC_9_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_16_LC_9_2_7  (
            .in0(_gnd_net_),
            .in1(N__18745),
            .in2(_gnd_net_),
            .in3(N__17069),
            .lcout(\COUNTER.counterZ0Z_16 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_15 ),
            .carryout(\COUNTER.counter_1_cry_16 ),
            .clk(N__20465),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_17_LC_9_3_0 .C_ON=1'b1;
    defparam \COUNTER.counter_17_LC_9_3_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_17_LC_9_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_17_LC_9_3_0  (
            .in0(_gnd_net_),
            .in1(N__18781),
            .in2(_gnd_net_),
            .in3(N__17066),
            .lcout(\COUNTER.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_9_3_0_),
            .carryout(\COUNTER.counter_1_cry_17 ),
            .clk(N__20408),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_18_LC_9_3_1 .C_ON=1'b1;
    defparam \COUNTER.counter_18_LC_9_3_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_18_LC_9_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_18_LC_9_3_1  (
            .in0(_gnd_net_),
            .in1(N__18796),
            .in2(_gnd_net_),
            .in3(N__17063),
            .lcout(\COUNTER.counterZ0Z_18 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_17 ),
            .carryout(\COUNTER.counter_1_cry_18 ),
            .clk(N__20408),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_19_LC_9_3_2 .C_ON=1'b1;
    defparam \COUNTER.counter_19_LC_9_3_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_19_LC_9_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_19_LC_9_3_2  (
            .in0(_gnd_net_),
            .in1(N__18766),
            .in2(_gnd_net_),
            .in3(N__17114),
            .lcout(\COUNTER.counterZ0Z_19 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_18 ),
            .carryout(\COUNTER.counter_1_cry_19 ),
            .clk(N__20408),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_20_LC_9_3_3 .C_ON=1'b1;
    defparam \COUNTER.counter_20_LC_9_3_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_20_LC_9_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_20_LC_9_3_3  (
            .in0(_gnd_net_),
            .in1(N__17282),
            .in2(_gnd_net_),
            .in3(N__17111),
            .lcout(\COUNTER.counterZ0Z_20 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_19 ),
            .carryout(\COUNTER.counter_1_cry_20 ),
            .clk(N__20408),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_21_LC_9_3_4 .C_ON=1'b1;
    defparam \COUNTER.counter_21_LC_9_3_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_21_LC_9_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_21_LC_9_3_4  (
            .in0(_gnd_net_),
            .in1(N__17309),
            .in2(_gnd_net_),
            .in3(N__17108),
            .lcout(\COUNTER.counterZ0Z_21 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_20 ),
            .carryout(\COUNTER.counter_1_cry_21 ),
            .clk(N__20408),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_22_LC_9_3_5 .C_ON=1'b1;
    defparam \COUNTER.counter_22_LC_9_3_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_22_LC_9_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_22_LC_9_3_5  (
            .in0(_gnd_net_),
            .in1(N__17321),
            .in2(_gnd_net_),
            .in3(N__17105),
            .lcout(\COUNTER.counterZ0Z_22 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_21 ),
            .carryout(\COUNTER.counter_1_cry_22 ),
            .clk(N__20408),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_23_LC_9_3_6 .C_ON=1'b1;
    defparam \COUNTER.counter_23_LC_9_3_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_23_LC_9_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_23_LC_9_3_6  (
            .in0(_gnd_net_),
            .in1(N__17296),
            .in2(_gnd_net_),
            .in3(N__17102),
            .lcout(\COUNTER.counterZ0Z_23 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_22 ),
            .carryout(\COUNTER.counter_1_cry_23 ),
            .clk(N__20408),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_24_LC_9_3_7 .C_ON=1'b1;
    defparam \COUNTER.counter_24_LC_9_3_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_24_LC_9_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_24_LC_9_3_7  (
            .in0(_gnd_net_),
            .in1(N__17179),
            .in2(_gnd_net_),
            .in3(N__17099),
            .lcout(\COUNTER.counterZ0Z_24 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_23 ),
            .carryout(\COUNTER.counter_1_cry_24 ),
            .clk(N__20408),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_25_LC_9_4_0 .C_ON=1'b1;
    defparam \COUNTER.counter_25_LC_9_4_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_25_LC_9_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_25_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(N__17207),
            .in2(_gnd_net_),
            .in3(N__17096),
            .lcout(\COUNTER.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_9_4_0_),
            .carryout(\COUNTER.counter_1_cry_25 ),
            .clk(N__20491),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_26_LC_9_4_1 .C_ON=1'b1;
    defparam \COUNTER.counter_26_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_26_LC_9_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_26_LC_9_4_1  (
            .in0(_gnd_net_),
            .in1(N__17219),
            .in2(_gnd_net_),
            .in3(N__17093),
            .lcout(\COUNTER.counterZ0Z_26 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_25 ),
            .carryout(\COUNTER.counter_1_cry_26 ),
            .clk(N__20491),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_27_LC_9_4_2 .C_ON=1'b1;
    defparam \COUNTER.counter_27_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_27_LC_9_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_27_LC_9_4_2  (
            .in0(_gnd_net_),
            .in1(N__17194),
            .in2(_gnd_net_),
            .in3(N__17090),
            .lcout(\COUNTER.counterZ0Z_27 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_26 ),
            .carryout(\COUNTER.counter_1_cry_27 ),
            .clk(N__20491),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_28_LC_9_4_3 .C_ON=1'b1;
    defparam \COUNTER.counter_28_LC_9_4_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_28_LC_9_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_28_LC_9_4_3  (
            .in0(_gnd_net_),
            .in1(N__17153),
            .in2(_gnd_net_),
            .in3(N__17333),
            .lcout(\COUNTER.counterZ0Z_28 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_27 ),
            .carryout(\COUNTER.counter_1_cry_28 ),
            .clk(N__20491),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_29_LC_9_4_4 .C_ON=1'b1;
    defparam \COUNTER.counter_29_LC_9_4_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_29_LC_9_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_29_LC_9_4_4  (
            .in0(_gnd_net_),
            .in1(N__17140),
            .in2(_gnd_net_),
            .in3(N__17330),
            .lcout(\COUNTER.counterZ0Z_29 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_28 ),
            .carryout(\COUNTER.counter_1_cry_29 ),
            .clk(N__20491),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_30_LC_9_4_5 .C_ON=1'b1;
    defparam \COUNTER.counter_30_LC_9_4_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_30_LC_9_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_30_LC_9_4_5  (
            .in0(_gnd_net_),
            .in1(N__17165),
            .in2(_gnd_net_),
            .in3(N__17327),
            .lcout(\COUNTER.counterZ0Z_30 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_29 ),
            .carryout(\COUNTER.counter_1_cry_30 ),
            .clk(N__20491),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_31_LC_9_4_6 .C_ON=1'b0;
    defparam \COUNTER.counter_31_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_31_LC_9_4_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.counter_31_LC_9_4_6  (
            .in0(_gnd_net_),
            .in1(N__17126),
            .in2(_gnd_net_),
            .in3(N__17324),
            .lcout(\COUNTER.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20491),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_RNO_LC_9_4_7 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_9_4_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_5_c_RNO_LC_9_4_7  (
            .in0(N__17320),
            .in1(N__17308),
            .in2(N__17297),
            .in3(N__17281),
            .lcout(\COUNTER.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_RNI027U_11_LC_9_5_0 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_RNI027U_11_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_RNI027U_11_LC_9_5_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ALL_SYS_PWRGD.count_RNI027U_11_LC_9_5_0  (
            .in0(N__17269),
            .in1(N__17257),
            .in2(N__17246),
            .in3(N__17230),
            .lcout(\ALL_SYS_PWRGD.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_0_LC_9_5_1 .C_ON=1'b0;
    defparam \COUNTER.counter_0_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_0_LC_9_5_1 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \COUNTER.counter_0_LC_9_5_1  (
            .in0(N__19435),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17577),
            .lcout(\COUNTER.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20458),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_RNO_LC_9_5_2 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_9_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_6_c_RNO_LC_9_5_2  (
            .in0(N__17218),
            .in1(N__17206),
            .in2(N__17195),
            .in3(N__17180),
            .lcout(\COUNTER.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_RNO_LC_9_5_3 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_9_5_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_7_c_RNO_LC_9_5_3  (
            .in0(N__17164),
            .in1(N__17152),
            .in2(N__17141),
            .in3(N__17125),
            .lcout(\COUNTER.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_4_LC_9_5_4 .C_ON=1'b0;
    defparam \COUNTER.counter_4_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_4_LC_9_5_4 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_4_LC_9_5_4  (
            .in0(N__17624),
            .in1(N__17607),
            .in2(_gnd_net_),
            .in3(N__19434),
            .lcout(\COUNTER.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20458),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_RNO_LC_9_5_5 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_9_5_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_RNO_LC_9_5_5  (
            .in0(N__17514),
            .in1(N__17544),
            .in2(N__17611),
            .in3(N__17576),
            .lcout(\COUNTER.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_2_LC_9_5_6 .C_ON=1'b0;
    defparam \COUNTER.counter_2_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_2_LC_9_5_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_2_LC_9_5_6  (
            .in0(N__17545),
            .in1(N__17561),
            .in2(_gnd_net_),
            .in3(N__19432),
            .lcout(\COUNTER.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20458),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_3_LC_9_5_7 .C_ON=1'b0;
    defparam \COUNTER.counter_3_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_3_LC_9_5_7 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \COUNTER.counter_3_LC_9_5_7  (
            .in0(N__19433),
            .in1(_gnd_net_),
            .in2(N__17521),
            .in3(N__17531),
            .lcout(\COUNTER.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20458),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_9_6_1 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_9_6_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_9_6_1  (
            .in0(N__17500),
            .in1(N__17488),
            .in2(N__17477),
            .in3(N__17461),
            .lcout(\ALL_SYS_PWRGD.un4_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_9_6_4 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_9_6_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_9_6_4  (
            .in0(N__17449),
            .in1(N__17437),
            .in2(N__17426),
            .in3(N__17410),
            .lcout(),
            .ltout(\ALL_SYS_PWRGD.un4_count_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_9_6_5 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_9_6_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_9_6_5  (
            .in0(N__17399),
            .in1(N__17897),
            .in2(N__17393),
            .in3(N__17390),
            .lcout(\ALL_SYS_PWRGD.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_RNIV07U_10_LC_9_6_7 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_RNIV07U_10_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_RNIV07U_10_LC_9_6_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \ALL_SYS_PWRGD.count_RNIV07U_10_LC_9_6_7  (
            .in0(N__17383),
            .in1(N__17371),
            .in2(N__17360),
            .in3(N__17344),
            .lcout(\ALL_SYS_PWRGD.un4_count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_RNIKNST6_0_LC_9_7_1 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_RNIKNST6_0_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_RNIKNST6_0_LC_9_7_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_RNIKNST6_0_LC_9_7_1  (
            .in0(N__19337),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20057),
            .lcout(\ALL_SYS_PWRGD.curr_state_RNIKNST6Z0Z_0 ),
            .ltout(\ALL_SYS_PWRGD.curr_state_RNIKNST6Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_9_7_2 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_9_7_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_9_7_2  (
            .in0(N__20058),
            .in1(_gnd_net_),
            .in2(N__17861),
            .in3(_gnd_net_),
            .lcout(\ALL_SYS_PWRGD.N_65_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_9_7_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_9_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_9_7_3  (
            .in0(N__17841),
            .in1(N__17819),
            .in2(N__17804),
            .in3(N__17776),
            .lcout(rsmrst_pwrgd_signal),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_LC_9_7_4 .C_ON=1'b0;
    defparam \COUNTER.tmp_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_LC_9_7_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \COUNTER.tmp_LC_9_7_4  (
            .in0(N__19431),
            .in1(_gnd_net_),
            .in2(N__17750),
            .in3(_gnd_net_),
            .lcout(\COUNTER.tmp_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20495),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_RNIRH3P_LC_9_7_5 .C_ON=1'b0;
    defparam \COUNTER.tmp_RNIRH3P_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_RNIRH3P_LC_9_7_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \COUNTER.tmp_RNIRH3P_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__17746),
            .in2(_gnd_net_),
            .in3(N__19430),
            .lcout(tmp_RNIRH3P),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_0_LC_9_9_0 .C_ON=1'b1;
    defparam \POWERLED.count_clk_0_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_0_LC_9_9_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_0_LC_9_9_0  (
            .in0(N__20092),
            .in1(N__17681),
            .in2(N__17702),
            .in3(N__17701),
            .lcout(\POWERLED.count_clkZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\POWERLED.un1_count_clk_1_cry_0 ),
            .clk(N__20558),
            .ce(),
            .sr(N__18251));
    defparam \POWERLED.count_clk_1_LC_9_9_1 .C_ON=1'b1;
    defparam \POWERLED.count_clk_1_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_1_LC_9_9_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_1_LC_9_9_1  (
            .in0(N__20085),
            .in1(N__17669),
            .in2(_gnd_net_),
            .in3(N__17651),
            .lcout(\POWERLED.count_clkZ0Z_1 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_0 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_1 ),
            .clk(N__20558),
            .ce(),
            .sr(N__18251));
    defparam \POWERLED.count_clk_2_LC_9_9_2 .C_ON=1'b1;
    defparam \POWERLED.count_clk_2_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_2_LC_9_9_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_2_LC_9_9_2  (
            .in0(N__20093),
            .in1(N__17647),
            .in2(_gnd_net_),
            .in3(N__17627),
            .lcout(\POWERLED.count_clkZ0Z_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_1 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_2 ),
            .clk(N__20558),
            .ce(),
            .sr(N__18251));
    defparam \POWERLED.count_clk_3_LC_9_9_3 .C_ON=1'b1;
    defparam \POWERLED.count_clk_3_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_3_LC_9_9_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_3_LC_9_9_3  (
            .in0(N__20086),
            .in1(N__18116),
            .in2(_gnd_net_),
            .in3(N__18101),
            .lcout(\POWERLED.count_clkZ0Z_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_2 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_3 ),
            .clk(N__20558),
            .ce(),
            .sr(N__18251));
    defparam \POWERLED.count_clk_4_LC_9_9_4 .C_ON=1'b1;
    defparam \POWERLED.count_clk_4_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_4_LC_9_9_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_4_LC_9_9_4  (
            .in0(N__20094),
            .in1(N__18098),
            .in2(_gnd_net_),
            .in3(N__18083),
            .lcout(\POWERLED.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_3 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_4 ),
            .clk(N__20558),
            .ce(),
            .sr(N__18251));
    defparam \POWERLED.count_clk_5_LC_9_9_5 .C_ON=1'b1;
    defparam \POWERLED.count_clk_5_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_5_LC_9_9_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_5_LC_9_9_5  (
            .in0(N__20087),
            .in1(N__18080),
            .in2(_gnd_net_),
            .in3(N__18059),
            .lcout(\POWERLED.count_clkZ0Z_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_4 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_5 ),
            .clk(N__20558),
            .ce(),
            .sr(N__18251));
    defparam \POWERLED.count_clk_6_LC_9_9_6 .C_ON=1'b1;
    defparam \POWERLED.count_clk_6_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_6_LC_9_9_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_6_LC_9_9_6  (
            .in0(N__20095),
            .in1(N__18051),
            .in2(_gnd_net_),
            .in3(N__18023),
            .lcout(\POWERLED.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_5 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_6 ),
            .clk(N__20558),
            .ce(),
            .sr(N__18251));
    defparam \POWERLED.count_clk_7_LC_9_9_7 .C_ON=1'b1;
    defparam \POWERLED.count_clk_7_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_7_LC_9_9_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_7_LC_9_9_7  (
            .in0(N__20088),
            .in1(N__18000),
            .in2(_gnd_net_),
            .in3(N__17954),
            .lcout(\POWERLED.count_clkZ0Z_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_6 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_7 ),
            .clk(N__20558),
            .ce(),
            .sr(N__18251));
    defparam \POWERLED.count_clk_8_LC_9_10_0 .C_ON=1'b1;
    defparam \POWERLED.count_clk_8_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_8_LC_9_10_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_8_LC_9_10_0  (
            .in0(N__20099),
            .in1(N__17951),
            .in2(_gnd_net_),
            .in3(N__17936),
            .lcout(\POWERLED.count_clkZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\POWERLED.un1_count_clk_1_cry_8 ),
            .clk(N__20543),
            .ce(),
            .sr(N__18243));
    defparam \POWERLED.count_clk_9_LC_9_10_1 .C_ON=1'b1;
    defparam \POWERLED.count_clk_9_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_9_LC_9_10_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_9_LC_9_10_1  (
            .in0(N__20091),
            .in1(N__17933),
            .in2(_gnd_net_),
            .in3(N__17915),
            .lcout(\POWERLED.count_clkZ0Z_9 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_8 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_9 ),
            .clk(N__20543),
            .ce(),
            .sr(N__18243));
    defparam \POWERLED.count_clk_10_LC_9_10_2 .C_ON=1'b1;
    defparam \POWERLED.count_clk_10_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_10_LC_9_10_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_10_LC_9_10_2  (
            .in0(N__20096),
            .in1(N__17912),
            .in2(_gnd_net_),
            .in3(N__17900),
            .lcout(\POWERLED.count_clkZ0Z_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_9 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_10 ),
            .clk(N__20543),
            .ce(),
            .sr(N__18243));
    defparam \POWERLED.count_clk_11_LC_9_10_3 .C_ON=1'b1;
    defparam \POWERLED.count_clk_11_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_11_LC_9_10_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_11_LC_9_10_3  (
            .in0(N__20089),
            .in1(N__18458),
            .in2(_gnd_net_),
            .in3(N__18446),
            .lcout(\POWERLED.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_10 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_11 ),
            .clk(N__20543),
            .ce(),
            .sr(N__18243));
    defparam \POWERLED.count_clk_12_LC_9_10_4 .C_ON=1'b1;
    defparam \POWERLED.count_clk_12_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_12_LC_9_10_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_12_LC_9_10_4  (
            .in0(N__20097),
            .in1(N__18443),
            .in2(_gnd_net_),
            .in3(N__18431),
            .lcout(\POWERLED.count_clkZ0Z_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_11 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_12 ),
            .clk(N__20543),
            .ce(),
            .sr(N__18243));
    defparam \POWERLED.count_clk_13_LC_9_10_5 .C_ON=1'b1;
    defparam \POWERLED.count_clk_13_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_13_LC_9_10_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_13_LC_9_10_5  (
            .in0(N__20090),
            .in1(N__18427),
            .in2(_gnd_net_),
            .in3(N__18413),
            .lcout(\POWERLED.count_clkZ0Z_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_12 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_13 ),
            .clk(N__20543),
            .ce(),
            .sr(N__18243));
    defparam \POWERLED.count_clk_14_LC_9_10_6 .C_ON=1'b1;
    defparam \POWERLED.count_clk_14_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_14_LC_9_10_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_14_LC_9_10_6  (
            .in0(N__20098),
            .in1(N__18410),
            .in2(_gnd_net_),
            .in3(N__18398),
            .lcout(\POWERLED.count_clkZ0Z_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_13 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_14 ),
            .clk(N__20543),
            .ce(),
            .sr(N__18243));
    defparam \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_9_10_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_9_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__18356),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_14 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_esr_15_LC_9_11_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_esr_15_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_esr_15_LC_9_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.count_clk_esr_15_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__18280),
            .in2(_gnd_net_),
            .in3(N__18284),
            .lcout(\POWERLED.count_clkZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20559),
            .ce(N__18266),
            .sr(N__18250));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_11_LC_9_12_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_11_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_11_LC_9_12_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_11_LC_9_12_1  (
            .in0(N__18217),
            .in1(N__18205),
            .in2(N__18194),
            .in3(N__18178),
            .lcout(\RSMRST_PWRGD.m4_i_i_a2_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_9_LC_9_12_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_9_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_9_LC_9_12_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_9_LC_9_12_3  (
            .in0(N__18166),
            .in1(N__18154),
            .in2(N__18143),
            .in3(N__18127),
            .lcout(),
            .ltout(\RSMRST_PWRGD.m4_i_i_a2_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_LC_9_12_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_LC_9_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_LC_9_12_4  (
            .in0(N__18656),
            .in1(N__18539),
            .in2(N__18650),
            .in3(N__18596),
            .lcout(\RSMRST_PWRGD.N_241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_7_LC_9_12_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_7_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_7_LC_9_12_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_7_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__18646),
            .in2(_gnd_net_),
            .in3(N__18634),
            .lcout(),
            .ltout(\RSMRST_PWRGD.m4_i_i_a2_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_12_LC_9_12_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_12_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_12_LC_9_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_12_LC_9_12_6  (
            .in0(N__18622),
            .in1(N__19229),
            .in2(N__18611),
            .in3(N__18607),
            .lcout(\RSMRST_PWRGD.m4_i_i_a2_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_10_LC_9_12_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_10_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_10_LC_9_12_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_10_LC_9_12_7  (
            .in0(N__18589),
            .in1(N__18577),
            .in2(N__18566),
            .in3(N__18550),
            .lcout(\RSMRST_PWRGD.m4_i_i_a2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_9_13_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_9_13_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_9_13_0  (
            .in0(N__19524),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19227),
            .lcout(\RSMRST_PWRGD.N_240 ),
            .ltout(\RSMRST_PWRGD.N_240_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNIJULM7_0_LC_9_13_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNIJULM7_0_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNIJULM7_0_LC_9_13_1 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNIJULM7_0_LC_9_13_1  (
            .in0(N__19186),
            .in1(N__20747),
            .in2(N__18533),
            .in3(N__20064),
            .lcout(\RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0 ),
            .ltout(\RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_13_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_13_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_13_2  (
            .in0(N__20065),
            .in1(_gnd_net_),
            .in2(N__18500),
            .in3(_gnd_net_),
            .lcout(\RSMRST_PWRGD.N_65_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_13_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_13_6 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_13_6  (
            .in0(N__19525),
            .in1(N__20746),
            .in2(_gnd_net_),
            .in3(N__19226),
            .lcout(\RSMRST_PWRGD.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_9_14_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_9_14_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_RNIVJP51_3_LC_9_14_1  (
            .in0(N__18469),
            .in1(N__19096),
            .in2(N__19085),
            .in3(N__19069),
            .lcout(\VPP_VDDQ.un6_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_15_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_15_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_15_3  (
            .in0(N__19057),
            .in1(N__19045),
            .in2(N__19034),
            .in3(N__19018),
            .lcout(\VPP_VDDQ.un6_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI63141_10_LC_9_15_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_9_15_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_RNI63141_10_LC_9_15_5  (
            .in0(N__19006),
            .in1(N__18994),
            .in2(N__18983),
            .in3(N__18967),
            .lcout(\VPP_VDDQ.un6_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_9_15_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_9_15_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \VPP_VDDQ.count_RNIFC141_11_LC_9_15_6  (
            .in0(N__18956),
            .in1(N__18940),
            .in2(N__18929),
            .in3(N__18913),
            .lcout(),
            .ltout(\VPP_VDDQ.un6_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_15_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_15_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_15_7  (
            .in0(N__18902),
            .in1(N__18896),
            .in2(N__18890),
            .in3(N__18887),
            .lcout(\VPP_VDDQ.count_esr_RNIRFM64Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_RNO_LC_11_2_1 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_11_2_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_3_c_RNO_LC_11_2_1  (
            .in0(N__18860),
            .in1(N__18845),
            .in2(N__18830),
            .in3(N__18812),
            .lcout(\COUNTER.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_RNO_LC_11_3_3 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_11_3_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_4_c_RNO_LC_11_3_3  (
            .in0(N__18797),
            .in1(N__18782),
            .in2(N__18767),
            .in3(N__18749),
            .lcout(\COUNTER.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_RNO_LC_11_3_5 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_11_3_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_2_c_RNO_LC_11_3_5  (
            .in0(N__18731),
            .in1(N__18713),
            .in2(N__18695),
            .in3(N__18674),
            .lcout(\COUNTER.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_LC_11_5_0 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_0_c_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_LC_11_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_LC_11_5_0  (
            .in0(_gnd_net_),
            .in1(N__19175),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(\COUNTER.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_LC_11_5_1 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_1_c_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_LC_11_5_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_1_c_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__19166),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_0 ),
            .carryout(\COUNTER.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_LC_11_5_2 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_2_c_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_LC_11_5_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_2_c_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(N__19154),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_1 ),
            .carryout(\COUNTER.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_LC_11_5_3 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_3_c_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_LC_11_5_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_3_c_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__19145),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_2 ),
            .carryout(\COUNTER.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_LC_11_5_4 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_4_c_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_LC_11_5_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_4_c_LC_11_5_4  (
            .in0(_gnd_net_),
            .in1(N__19136),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_3 ),
            .carryout(\COUNTER.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_LC_11_5_5 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_5_c_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_LC_11_5_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_5_c_LC_11_5_5  (
            .in0(_gnd_net_),
            .in1(N__19127),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_4 ),
            .carryout(\COUNTER.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_LC_11_5_6 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_6_c_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_LC_11_5_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_6_c_LC_11_5_6  (
            .in0(_gnd_net_),
            .in1(N__19115),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_5 ),
            .carryout(\COUNTER.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_LC_11_5_7 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_7_c_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_LC_11_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_7_c_LC_11_5_7  (
            .in0(_gnd_net_),
            .in1(N__19106),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_6 ),
            .carryout(\COUNTER.un4_counter_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_THRU_LUT4_0_LC_11_6_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_THRU_LUT4_0_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_THRU_LUT4_0_LC_11_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.un4_counter_7_THRU_LUT4_0_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19448),
            .lcout(\COUNTER.un4_counter_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_LC_11_7_2 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_LC_11_7_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_LC_11_7_2  (
            .in0(N__19304),
            .in1(N__19470),
            .in2(_gnd_net_),
            .in3(N__19325),
            .lcout(),
            .ltout(\ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_0_LC_11_7_3 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_0_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.curr_state_0_LC_11_7_3 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_0_LC_11_7_3  (
            .in0(N__19328),
            .in1(N__19360),
            .in2(N__19388),
            .in3(N__19307),
            .lcout(\ALL_SYS_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20538),
            .ce(N__19802),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_RNIUU4I2_0_LC_11_7_4 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_RNIUU4I2_0_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_RNIUU4I2_0_LC_11_7_4 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_RNIUU4I2_0_LC_11_7_4  (
            .in0(N__19303),
            .in1(N__19471),
            .in2(_gnd_net_),
            .in3(N__19324),
            .lcout(\ALL_SYS_PWRGD.un1_curr_state10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_1_LC_11_7_5 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_1_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.curr_state_1_LC_11_7_5 .LUT_INIT=16'b0000010101000100;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_1_LC_11_7_5  (
            .in0(N__19327),
            .in1(N__19466),
            .in2(N__19361),
            .in3(N__19306),
            .lcout(\ALL_SYS_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20538),
            .ce(N__19802),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_RNIP5P46_0_LC_11_7_6 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_RNIP5P46_0_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_RNIP5P46_0_LC_11_7_6 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_RNIP5P46_0_LC_11_7_6  (
            .in0(N__19302),
            .in1(N__19323),
            .in2(N__19472),
            .in3(N__19356),
            .lcout(\ALL_SYS_PWRGD.N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_11_7_7 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_11_7_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_11_7_7  (
            .in0(N__19326),
            .in1(N__19465),
            .in2(_gnd_net_),
            .in3(N__19305),
            .lcout(vccst_pwrgd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20538),
            .ce(N__19802),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_1_LC_11_13_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_1_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_1_LC_11_13_5 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \RSMRST_PWRGD.curr_state_1_LC_11_13_5  (
            .in0(N__20743),
            .in1(N__19532),
            .in2(N__19228),
            .in3(N__19195),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20594),
            .ce(N__19810),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_0_LC_11_13_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_0_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_0_LC_11_13_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \RSMRST_PWRGD.curr_state_0_LC_11_13_7  (
            .in0(N__20744),
            .in1(N__20764),
            .in2(_gnd_net_),
            .in3(N__19196),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20594),
            .ce(N__19810),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_LC_11_14_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_LC_11_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__20768),
            .in2(_gnd_net_),
            .in3(N__20745),
            .lcout(rsmrstn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20595),
            .ce(N__19809),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_1_LC_12_7_3 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_1_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_1_LC_12_7_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_1_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(N__19562),
            .in2(_gnd_net_),
            .in3(N__19538),
            .lcout(),
            .ltout(\ALL_SYS_PWRGD.m4_0_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_LC_12_7_4 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_LC_12_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_LC_12_7_4  (
            .in0(N__19523),
            .in1(N__19499),
            .in2(N__19487),
            .in3(N__19484),
            .lcout(\ALL_SYS_PWRGD.N_245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TOP
