// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 11 2022 18:27:59

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VCCST_ENn,
    GPIO_FPGA_PM_3,
    GPIO_FPGA_PCH_2,
    VR_READY_VCCINAUX,
    VCCST_OK,
    VCCIO_EN,
    V33A_ENn,
    V1P8A_EN,
    GPIO_FPGA_SV_4,
    GPIO_FPGA_PM_4,
    VDDQ_EN,
    V5S_OK,
    SLP_S3n,
    GPIO_FPGA_PCH_4,
    VCCIO_OK,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    SLP_SUSn,
    MAIN_12V_MON,
    GPIO_FPGA_SV_3,
    GPIO_FPGA_HDR_3,
    V33DSW_OK,
    TPM_GPIO,
    PLTRSTn,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    GPIO_FPGA_SV_1,
    GPIO_FPGA_HDR_1,
    FPGA_OSC,
    VCCST_PWRGD,
    V105A_EN,
    SYS_PWROK,
    GPIO_FPGA_PM_2,
    GPIO_FPGA_PCH_1,
    HDA_SDO_FPGA,
    VPP_EN,
    VDDQ_OK,
    SLP_S4n,
    GPIO_FPGA_PCH_3,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    V1P8_OK,
    DSW_PWROK,
    PM_PWROK,
    GPIO_FPGA_SV_2,
    GPIO_FPGA_PCH_5,
    V5A_EN,
    FPGA_GPIO_WD,
    VPP_OK,
    VCCIN_EN,
    V105A_OK,
    SLP_S5n,
    GPIO_FPGA_HDR_2,
    FP_RSTn,
    GPIO_FPGA_PM_1,
    V33A_OK,
    PCH_PWROK);

    output VCCST_ENn;
    input GPIO_FPGA_PM_3;
    input GPIO_FPGA_PCH_2;
    input VR_READY_VCCINAUX;
    input VCCST_OK;
    output VCCIO_EN;
    output V33A_ENn;
    output V1P8A_EN;
    input GPIO_FPGA_SV_4;
    input GPIO_FPGA_PM_4;
    output VDDQ_EN;
    input V5S_OK;
    input SLP_S3n;
    input GPIO_FPGA_PCH_4;
    input VCCIO_OK;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input SLP_SUSn;
    input MAIN_12V_MON;
    input GPIO_FPGA_SV_3;
    input GPIO_FPGA_HDR_3;
    input V33DSW_OK;
    input TPM_GPIO;
    input PLTRSTn;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input GPIO_FPGA_SV_1;
    input GPIO_FPGA_HDR_1;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output V105A_EN;
    output SYS_PWROK;
    input GPIO_FPGA_PM_2;
    input GPIO_FPGA_PCH_1;
    output HDA_SDO_FPGA;
    output VPP_EN;
    input VDDQ_OK;
    input SLP_S4n;
    input GPIO_FPGA_PCH_3;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input V1P8_OK;
    output DSW_PWROK;
    input PM_PWROK;
    input GPIO_FPGA_SV_2;
    input GPIO_FPGA_PCH_5;
    output V5A_EN;
    input FPGA_GPIO_WD;
    input VPP_OK;
    output VCCIN_EN;
    input V105A_OK;
    input SLP_S5n;
    input GPIO_FPGA_HDR_2;
    input FP_RSTn;
    input GPIO_FPGA_PM_1;
    input V33A_OK;
    output PCH_PWROK;

    wire N__35653;
    wire N__35652;
    wire N__35651;
    wire N__35642;
    wire N__35641;
    wire N__35640;
    wire N__35633;
    wire N__35632;
    wire N__35631;
    wire N__35624;
    wire N__35623;
    wire N__35622;
    wire N__35615;
    wire N__35614;
    wire N__35613;
    wire N__35606;
    wire N__35605;
    wire N__35604;
    wire N__35597;
    wire N__35596;
    wire N__35595;
    wire N__35588;
    wire N__35587;
    wire N__35586;
    wire N__35579;
    wire N__35578;
    wire N__35577;
    wire N__35570;
    wire N__35569;
    wire N__35568;
    wire N__35561;
    wire N__35560;
    wire N__35559;
    wire N__35552;
    wire N__35551;
    wire N__35550;
    wire N__35543;
    wire N__35542;
    wire N__35541;
    wire N__35534;
    wire N__35533;
    wire N__35532;
    wire N__35525;
    wire N__35524;
    wire N__35523;
    wire N__35516;
    wire N__35515;
    wire N__35514;
    wire N__35507;
    wire N__35506;
    wire N__35505;
    wire N__35498;
    wire N__35497;
    wire N__35496;
    wire N__35489;
    wire N__35488;
    wire N__35487;
    wire N__35480;
    wire N__35479;
    wire N__35478;
    wire N__35471;
    wire N__35470;
    wire N__35469;
    wire N__35462;
    wire N__35461;
    wire N__35460;
    wire N__35453;
    wire N__35452;
    wire N__35451;
    wire N__35444;
    wire N__35443;
    wire N__35442;
    wire N__35435;
    wire N__35434;
    wire N__35433;
    wire N__35426;
    wire N__35425;
    wire N__35424;
    wire N__35417;
    wire N__35416;
    wire N__35415;
    wire N__35408;
    wire N__35407;
    wire N__35406;
    wire N__35399;
    wire N__35398;
    wire N__35397;
    wire N__35390;
    wire N__35389;
    wire N__35388;
    wire N__35381;
    wire N__35380;
    wire N__35379;
    wire N__35372;
    wire N__35371;
    wire N__35370;
    wire N__35363;
    wire N__35362;
    wire N__35361;
    wire N__35354;
    wire N__35353;
    wire N__35352;
    wire N__35345;
    wire N__35344;
    wire N__35343;
    wire N__35336;
    wire N__35335;
    wire N__35334;
    wire N__35327;
    wire N__35326;
    wire N__35325;
    wire N__35308;
    wire N__35307;
    wire N__35304;
    wire N__35301;
    wire N__35298;
    wire N__35297;
    wire N__35296;
    wire N__35295;
    wire N__35294;
    wire N__35293;
    wire N__35292;
    wire N__35291;
    wire N__35290;
    wire N__35285;
    wire N__35280;
    wire N__35279;
    wire N__35278;
    wire N__35277;
    wire N__35276;
    wire N__35275;
    wire N__35274;
    wire N__35273;
    wire N__35272;
    wire N__35271;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35255;
    wire N__35250;
    wire N__35239;
    wire N__35234;
    wire N__35229;
    wire N__35228;
    wire N__35227;
    wire N__35226;
    wire N__35225;
    wire N__35224;
    wire N__35223;
    wire N__35222;
    wire N__35219;
    wire N__35214;
    wire N__35211;
    wire N__35206;
    wire N__35205;
    wire N__35204;
    wire N__35203;
    wire N__35202;
    wire N__35201;
    wire N__35196;
    wire N__35193;
    wire N__35186;
    wire N__35179;
    wire N__35178;
    wire N__35175;
    wire N__35168;
    wire N__35157;
    wire N__35154;
    wire N__35147;
    wire N__35144;
    wire N__35131;
    wire N__35130;
    wire N__35127;
    wire N__35126;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35095;
    wire N__35094;
    wire N__35093;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35083;
    wire N__35080;
    wire N__35077;
    wire N__35074;
    wire N__35071;
    wire N__35062;
    wire N__35059;
    wire N__35058;
    wire N__35055;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35042;
    wire N__35039;
    wire N__35036;
    wire N__35033;
    wire N__35026;
    wire N__35025;
    wire N__35022;
    wire N__35021;
    wire N__35020;
    wire N__35017;
    wire N__35016;
    wire N__35013;
    wire N__35008;
    wire N__35005;
    wire N__35002;
    wire N__34999;
    wire N__34996;
    wire N__34987;
    wire N__34984;
    wire N__34981;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34963;
    wire N__34960;
    wire N__34959;
    wire N__34954;
    wire N__34951;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34941;
    wire N__34940;
    wire N__34939;
    wire N__34938;
    wire N__34937;
    wire N__34936;
    wire N__34935;
    wire N__34930;
    wire N__34929;
    wire N__34928;
    wire N__34917;
    wire N__34916;
    wire N__34915;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34905;
    wire N__34904;
    wire N__34903;
    wire N__34900;
    wire N__34897;
    wire N__34896;
    wire N__34895;
    wire N__34894;
    wire N__34891;
    wire N__34886;
    wire N__34881;
    wire N__34872;
    wire N__34869;
    wire N__34862;
    wire N__34849;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34837;
    wire N__34836;
    wire N__34831;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34819;
    wire N__34816;
    wire N__34815;
    wire N__34812;
    wire N__34809;
    wire N__34804;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34794;
    wire N__34789;
    wire N__34786;
    wire N__34783;
    wire N__34780;
    wire N__34777;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34756;
    wire N__34755;
    wire N__34754;
    wire N__34753;
    wire N__34744;
    wire N__34743;
    wire N__34740;
    wire N__34737;
    wire N__34732;
    wire N__34729;
    wire N__34726;
    wire N__34723;
    wire N__34720;
    wire N__34717;
    wire N__34716;
    wire N__34713;
    wire N__34710;
    wire N__34707;
    wire N__34704;
    wire N__34699;
    wire N__34696;
    wire N__34693;
    wire N__34690;
    wire N__34689;
    wire N__34688;
    wire N__34687;
    wire N__34686;
    wire N__34685;
    wire N__34684;
    wire N__34683;
    wire N__34682;
    wire N__34681;
    wire N__34680;
    wire N__34679;
    wire N__34678;
    wire N__34677;
    wire N__34676;
    wire N__34675;
    wire N__34674;
    wire N__34673;
    wire N__34672;
    wire N__34671;
    wire N__34670;
    wire N__34669;
    wire N__34668;
    wire N__34667;
    wire N__34666;
    wire N__34665;
    wire N__34664;
    wire N__34663;
    wire N__34662;
    wire N__34661;
    wire N__34660;
    wire N__34659;
    wire N__34658;
    wire N__34657;
    wire N__34656;
    wire N__34655;
    wire N__34654;
    wire N__34653;
    wire N__34652;
    wire N__34651;
    wire N__34650;
    wire N__34649;
    wire N__34648;
    wire N__34647;
    wire N__34646;
    wire N__34645;
    wire N__34644;
    wire N__34643;
    wire N__34642;
    wire N__34641;
    wire N__34640;
    wire N__34639;
    wire N__34638;
    wire N__34637;
    wire N__34636;
    wire N__34635;
    wire N__34634;
    wire N__34633;
    wire N__34632;
    wire N__34631;
    wire N__34630;
    wire N__34629;
    wire N__34628;
    wire N__34627;
    wire N__34626;
    wire N__34625;
    wire N__34624;
    wire N__34623;
    wire N__34622;
    wire N__34621;
    wire N__34620;
    wire N__34619;
    wire N__34618;
    wire N__34617;
    wire N__34616;
    wire N__34615;
    wire N__34614;
    wire N__34613;
    wire N__34612;
    wire N__34611;
    wire N__34610;
    wire N__34609;
    wire N__34608;
    wire N__34441;
    wire N__34438;
    wire N__34435;
    wire N__34434;
    wire N__34431;
    wire N__34430;
    wire N__34429;
    wire N__34428;
    wire N__34427;
    wire N__34426;
    wire N__34425;
    wire N__34422;
    wire N__34421;
    wire N__34420;
    wire N__34419;
    wire N__34418;
    wire N__34417;
    wire N__34416;
    wire N__34415;
    wire N__34414;
    wire N__34411;
    wire N__34408;
    wire N__34405;
    wire N__34396;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34382;
    wire N__34373;
    wire N__34372;
    wire N__34371;
    wire N__34370;
    wire N__34369;
    wire N__34368;
    wire N__34365;
    wire N__34358;
    wire N__34353;
    wire N__34350;
    wire N__34347;
    wire N__34346;
    wire N__34345;
    wire N__34342;
    wire N__34333;
    wire N__34330;
    wire N__34325;
    wire N__34318;
    wire N__34313;
    wire N__34310;
    wire N__34305;
    wire N__34294;
    wire N__34291;
    wire N__34288;
    wire N__34285;
    wire N__34284;
    wire N__34279;
    wire N__34276;
    wire N__34273;
    wire N__34270;
    wire N__34267;
    wire N__34264;
    wire N__34263;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34249;
    wire N__34246;
    wire N__34243;
    wire N__34242;
    wire N__34239;
    wire N__34236;
    wire N__34231;
    wire N__34230;
    wire N__34227;
    wire N__34224;
    wire N__34219;
    wire N__34216;
    wire N__34215;
    wire N__34214;
    wire N__34209;
    wire N__34206;
    wire N__34201;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34189;
    wire N__34188;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34174;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34162;
    wire N__34161;
    wire N__34156;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34146;
    wire N__34145;
    wire N__34142;
    wire N__34139;
    wire N__34136;
    wire N__34129;
    wire N__34126;
    wire N__34123;
    wire N__34120;
    wire N__34117;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34092;
    wire N__34091;
    wire N__34090;
    wire N__34089;
    wire N__34088;
    wire N__34087;
    wire N__34086;
    wire N__34085;
    wire N__34080;
    wire N__34079;
    wire N__34078;
    wire N__34077;
    wire N__34076;
    wire N__34075;
    wire N__34074;
    wire N__34073;
    wire N__34072;
    wire N__34071;
    wire N__34070;
    wire N__34069;
    wire N__34066;
    wire N__34065;
    wire N__34064;
    wire N__34061;
    wire N__34060;
    wire N__34059;
    wire N__34058;
    wire N__34057;
    wire N__34056;
    wire N__34055;
    wire N__34054;
    wire N__34053;
    wire N__34052;
    wire N__34051;
    wire N__34050;
    wire N__34041;
    wire N__34038;
    wire N__34037;
    wire N__34036;
    wire N__34033;
    wire N__34024;
    wire N__34017;
    wire N__34012;
    wire N__34007;
    wire N__34006;
    wire N__34003;
    wire N__33998;
    wire N__33995;
    wire N__33994;
    wire N__33991;
    wire N__33986;
    wire N__33983;
    wire N__33974;
    wire N__33967;
    wire N__33964;
    wire N__33957;
    wire N__33952;
    wire N__33949;
    wire N__33946;
    wire N__33943;
    wire N__33940;
    wire N__33933;
    wire N__33930;
    wire N__33929;
    wire N__33924;
    wire N__33919;
    wire N__33912;
    wire N__33907;
    wire N__33906;
    wire N__33905;
    wire N__33904;
    wire N__33899;
    wire N__33896;
    wire N__33891;
    wire N__33888;
    wire N__33885;
    wire N__33880;
    wire N__33877;
    wire N__33870;
    wire N__33863;
    wire N__33850;
    wire N__33849;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33831;
    wire N__33830;
    wire N__33823;
    wire N__33822;
    wire N__33821;
    wire N__33818;
    wire N__33813;
    wire N__33808;
    wire N__33807;
    wire N__33806;
    wire N__33805;
    wire N__33804;
    wire N__33803;
    wire N__33802;
    wire N__33797;
    wire N__33794;
    wire N__33785;
    wire N__33778;
    wire N__33777;
    wire N__33774;
    wire N__33771;
    wire N__33770;
    wire N__33769;
    wire N__33768;
    wire N__33767;
    wire N__33764;
    wire N__33759;
    wire N__33752;
    wire N__33749;
    wire N__33746;
    wire N__33743;
    wire N__33738;
    wire N__33735;
    wire N__33730;
    wire N__33727;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33717;
    wire N__33716;
    wire N__33715;
    wire N__33714;
    wire N__33713;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33698;
    wire N__33693;
    wire N__33690;
    wire N__33689;
    wire N__33688;
    wire N__33687;
    wire N__33686;
    wire N__33685;
    wire N__33684;
    wire N__33683;
    wire N__33682;
    wire N__33681;
    wire N__33680;
    wire N__33679;
    wire N__33678;
    wire N__33675;
    wire N__33672;
    wire N__33669;
    wire N__33666;
    wire N__33631;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33613;
    wire N__33610;
    wire N__33609;
    wire N__33608;
    wire N__33605;
    wire N__33604;
    wire N__33599;
    wire N__33596;
    wire N__33595;
    wire N__33594;
    wire N__33593;
    wire N__33592;
    wire N__33591;
    wire N__33590;
    wire N__33587;
    wire N__33586;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33570;
    wire N__33561;
    wire N__33558;
    wire N__33547;
    wire N__33544;
    wire N__33541;
    wire N__33538;
    wire N__33535;
    wire N__33532;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33522;
    wire N__33517;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33487;
    wire N__33484;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33472;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33460;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33450;
    wire N__33445;
    wire N__33444;
    wire N__33441;
    wire N__33438;
    wire N__33433;
    wire N__33430;
    wire N__33427;
    wire N__33424;
    wire N__33421;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33409;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33397;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33387;
    wire N__33382;
    wire N__33381;
    wire N__33378;
    wire N__33375;
    wire N__33370;
    wire N__33367;
    wire N__33364;
    wire N__33361;
    wire N__33358;
    wire N__33355;
    wire N__33354;
    wire N__33351;
    wire N__33348;
    wire N__33343;
    wire N__33342;
    wire N__33339;
    wire N__33336;
    wire N__33331;
    wire N__33330;
    wire N__33327;
    wire N__33324;
    wire N__33321;
    wire N__33316;
    wire N__33315;
    wire N__33312;
    wire N__33309;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33292;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33280;
    wire N__33279;
    wire N__33276;
    wire N__33273;
    wire N__33268;
    wire N__33267;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33253;
    wire N__33252;
    wire N__33249;
    wire N__33246;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33225;
    wire N__33222;
    wire N__33219;
    wire N__33214;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33202;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33187;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33148;
    wire N__33147;
    wire N__33144;
    wire N__33141;
    wire N__33138;
    wire N__33133;
    wire N__33130;
    wire N__33129;
    wire N__33126;
    wire N__33123;
    wire N__33120;
    wire N__33115;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33081;
    wire N__33078;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33066;
    wire N__33063;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33049;
    wire N__33046;
    wire N__33045;
    wire N__33044;
    wire N__33041;
    wire N__33038;
    wire N__33035;
    wire N__33028;
    wire N__33027;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32986;
    wire N__32985;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32970;
    wire N__32967;
    wire N__32964;
    wire N__32959;
    wire N__32956;
    wire N__32955;
    wire N__32954;
    wire N__32953;
    wire N__32952;
    wire N__32951;
    wire N__32950;
    wire N__32949;
    wire N__32948;
    wire N__32947;
    wire N__32946;
    wire N__32943;
    wire N__32932;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32908;
    wire N__32905;
    wire N__32904;
    wire N__32901;
    wire N__32898;
    wire N__32893;
    wire N__32892;
    wire N__32889;
    wire N__32886;
    wire N__32885;
    wire N__32884;
    wire N__32883;
    wire N__32882;
    wire N__32881;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32870;
    wire N__32869;
    wire N__32868;
    wire N__32867;
    wire N__32866;
    wire N__32865;
    wire N__32862;
    wire N__32861;
    wire N__32858;
    wire N__32855;
    wire N__32852;
    wire N__32849;
    wire N__32842;
    wire N__32841;
    wire N__32840;
    wire N__32839;
    wire N__32836;
    wire N__32835;
    wire N__32834;
    wire N__32833;
    wire N__32832;
    wire N__32829;
    wire N__32828;
    wire N__32825;
    wire N__32822;
    wire N__32819;
    wire N__32810;
    wire N__32809;
    wire N__32808;
    wire N__32807;
    wire N__32806;
    wire N__32805;
    wire N__32804;
    wire N__32803;
    wire N__32802;
    wire N__32799;
    wire N__32794;
    wire N__32791;
    wire N__32786;
    wire N__32779;
    wire N__32772;
    wire N__32765;
    wire N__32762;
    wire N__32757;
    wire N__32752;
    wire N__32747;
    wire N__32742;
    wire N__32737;
    wire N__32730;
    wire N__32725;
    wire N__32720;
    wire N__32707;
    wire N__32704;
    wire N__32701;
    wire N__32698;
    wire N__32695;
    wire N__32686;
    wire N__32683;
    wire N__32682;
    wire N__32681;
    wire N__32680;
    wire N__32679;
    wire N__32678;
    wire N__32675;
    wire N__32668;
    wire N__32665;
    wire N__32664;
    wire N__32661;
    wire N__32660;
    wire N__32659;
    wire N__32652;
    wire N__32651;
    wire N__32650;
    wire N__32649;
    wire N__32648;
    wire N__32647;
    wire N__32646;
    wire N__32645;
    wire N__32644;
    wire N__32643;
    wire N__32642;
    wire N__32641;
    wire N__32638;
    wire N__32637;
    wire N__32636;
    wire N__32635;
    wire N__32634;
    wire N__32633;
    wire N__32632;
    wire N__32631;
    wire N__32626;
    wire N__32623;
    wire N__32620;
    wire N__32615;
    wire N__32608;
    wire N__32599;
    wire N__32596;
    wire N__32589;
    wire N__32584;
    wire N__32581;
    wire N__32574;
    wire N__32571;
    wire N__32556;
    wire N__32553;
    wire N__32548;
    wire N__32547;
    wire N__32546;
    wire N__32543;
    wire N__32540;
    wire N__32535;
    wire N__32530;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32512;
    wire N__32509;
    wire N__32506;
    wire N__32505;
    wire N__32504;
    wire N__32501;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32491;
    wire N__32488;
    wire N__32485;
    wire N__32482;
    wire N__32473;
    wire N__32470;
    wire N__32469;
    wire N__32466;
    wire N__32463;
    wire N__32460;
    wire N__32455;
    wire N__32452;
    wire N__32449;
    wire N__32446;
    wire N__32443;
    wire N__32442;
    wire N__32441;
    wire N__32438;
    wire N__32433;
    wire N__32430;
    wire N__32425;
    wire N__32424;
    wire N__32419;
    wire N__32416;
    wire N__32415;
    wire N__32414;
    wire N__32407;
    wire N__32404;
    wire N__32401;
    wire N__32398;
    wire N__32397;
    wire N__32396;
    wire N__32393;
    wire N__32390;
    wire N__32387;
    wire N__32384;
    wire N__32377;
    wire N__32374;
    wire N__32371;
    wire N__32368;
    wire N__32367;
    wire N__32362;
    wire N__32359;
    wire N__32358;
    wire N__32357;
    wire N__32350;
    wire N__32347;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32335;
    wire N__32332;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32320;
    wire N__32317;
    wire N__32314;
    wire N__32311;
    wire N__32308;
    wire N__32305;
    wire N__32302;
    wire N__32299;
    wire N__32298;
    wire N__32297;
    wire N__32294;
    wire N__32289;
    wire N__32284;
    wire N__32283;
    wire N__32278;
    wire N__32275;
    wire N__32272;
    wire N__32269;
    wire N__32266;
    wire N__32263;
    wire N__32260;
    wire N__32259;
    wire N__32254;
    wire N__32251;
    wire N__32248;
    wire N__32245;
    wire N__32242;
    wire N__32241;
    wire N__32238;
    wire N__32237;
    wire N__32236;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32222;
    wire N__32215;
    wire N__32214;
    wire N__32209;
    wire N__32208;
    wire N__32207;
    wire N__32206;
    wire N__32205;
    wire N__32202;
    wire N__32201;
    wire N__32200;
    wire N__32199;
    wire N__32198;
    wire N__32197;
    wire N__32196;
    wire N__32195;
    wire N__32194;
    wire N__32193;
    wire N__32190;
    wire N__32183;
    wire N__32182;
    wire N__32181;
    wire N__32180;
    wire N__32179;
    wire N__32178;
    wire N__32177;
    wire N__32174;
    wire N__32167;
    wire N__32160;
    wire N__32153;
    wire N__32148;
    wire N__32147;
    wire N__32146;
    wire N__32145;
    wire N__32144;
    wire N__32143;
    wire N__32140;
    wire N__32137;
    wire N__32128;
    wire N__32125;
    wire N__32116;
    wire N__32105;
    wire N__32092;
    wire N__32089;
    wire N__32088;
    wire N__32087;
    wire N__32086;
    wire N__32085;
    wire N__32084;
    wire N__32083;
    wire N__32082;
    wire N__32081;
    wire N__32080;
    wire N__32077;
    wire N__32066;
    wire N__32057;
    wire N__32056;
    wire N__32055;
    wire N__32054;
    wire N__32053;
    wire N__32052;
    wire N__32051;
    wire N__32048;
    wire N__32043;
    wire N__32042;
    wire N__32039;
    wire N__32038;
    wire N__32035;
    wire N__32034;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32021;
    wire N__32018;
    wire N__32015;
    wire N__32008;
    wire N__32001;
    wire N__31984;
    wire N__31981;
    wire N__31978;
    wire N__31977;
    wire N__31976;
    wire N__31975;
    wire N__31974;
    wire N__31971;
    wire N__31970;
    wire N__31967;
    wire N__31966;
    wire N__31965;
    wire N__31964;
    wire N__31963;
    wire N__31962;
    wire N__31961;
    wire N__31960;
    wire N__31959;
    wire N__31958;
    wire N__31955;
    wire N__31946;
    wire N__31943;
    wire N__31936;
    wire N__31935;
    wire N__31934;
    wire N__31933;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31921;
    wire N__31916;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31908;
    wire N__31907;
    wire N__31904;
    wire N__31901;
    wire N__31892;
    wire N__31889;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31873;
    wire N__31868;
    wire N__31863;
    wire N__31860;
    wire N__31855;
    wire N__31840;
    wire N__31837;
    wire N__31836;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31828;
    wire N__31827;
    wire N__31824;
    wire N__31819;
    wire N__31816;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31804;
    wire N__31801;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31789;
    wire N__31786;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31770;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31750;
    wire N__31747;
    wire N__31744;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31732;
    wire N__31731;
    wire N__31726;
    wire N__31723;
    wire N__31720;
    wire N__31717;
    wire N__31716;
    wire N__31711;
    wire N__31708;
    wire N__31705;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31697;
    wire N__31694;
    wire N__31689;
    wire N__31684;
    wire N__31681;
    wire N__31680;
    wire N__31675;
    wire N__31672;
    wire N__31669;
    wire N__31666;
    wire N__31663;
    wire N__31660;
    wire N__31657;
    wire N__31656;
    wire N__31651;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31635;
    wire N__31634;
    wire N__31633;
    wire N__31630;
    wire N__31625;
    wire N__31622;
    wire N__31615;
    wire N__31612;
    wire N__31611;
    wire N__31608;
    wire N__31605;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31588;
    wire N__31585;
    wire N__31582;
    wire N__31581;
    wire N__31576;
    wire N__31573;
    wire N__31570;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31552;
    wire N__31549;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31534;
    wire N__31531;
    wire N__31530;
    wire N__31525;
    wire N__31522;
    wire N__31519;
    wire N__31516;
    wire N__31513;
    wire N__31510;
    wire N__31507;
    wire N__31506;
    wire N__31501;
    wire N__31498;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31488;
    wire N__31485;
    wire N__31484;
    wire N__31481;
    wire N__31478;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31466;
    wire N__31459;
    wire N__31456;
    wire N__31455;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31443;
    wire N__31440;
    wire N__31435;
    wire N__31434;
    wire N__31429;
    wire N__31426;
    wire N__31423;
    wire N__31420;
    wire N__31417;
    wire N__31414;
    wire N__31411;
    wire N__31410;
    wire N__31407;
    wire N__31406;
    wire N__31403;
    wire N__31398;
    wire N__31395;
    wire N__31390;
    wire N__31387;
    wire N__31384;
    wire N__31381;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31371;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31359;
    wire N__31354;
    wire N__31351;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31332;
    wire N__31327;
    wire N__31324;
    wire N__31321;
    wire N__31318;
    wire N__31315;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31296;
    wire N__31291;
    wire N__31288;
    wire N__31285;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31273;
    wire N__31270;
    wire N__31267;
    wire N__31264;
    wire N__31261;
    wire N__31258;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31240;
    wire N__31237;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31213;
    wire N__31210;
    wire N__31207;
    wire N__31204;
    wire N__31201;
    wire N__31198;
    wire N__31195;
    wire N__31192;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31171;
    wire N__31168;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31153;
    wire N__31150;
    wire N__31147;
    wire N__31144;
    wire N__31141;
    wire N__31140;
    wire N__31137;
    wire N__31136;
    wire N__31133;
    wire N__31130;
    wire N__31127;
    wire N__31120;
    wire N__31117;
    wire N__31114;
    wire N__31113;
    wire N__31112;
    wire N__31109;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31099;
    wire N__31096;
    wire N__31087;
    wire N__31084;
    wire N__31083;
    wire N__31080;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31070;
    wire N__31063;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31051;
    wire N__31048;
    wire N__31045;
    wire N__31044;
    wire N__31043;
    wire N__31040;
    wire N__31037;
    wire N__31034;
    wire N__31031;
    wire N__31028;
    wire N__31021;
    wire N__31018;
    wire N__31015;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31005;
    wire N__31002;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30985;
    wire N__30982;
    wire N__30979;
    wire N__30976;
    wire N__30973;
    wire N__30970;
    wire N__30967;
    wire N__30966;
    wire N__30965;
    wire N__30962;
    wire N__30957;
    wire N__30952;
    wire N__30949;
    wire N__30946;
    wire N__30943;
    wire N__30940;
    wire N__30937;
    wire N__30934;
    wire N__30933;
    wire N__30930;
    wire N__30929;
    wire N__30926;
    wire N__30923;
    wire N__30918;
    wire N__30913;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30891;
    wire N__30888;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30868;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30847;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30819;
    wire N__30818;
    wire N__30811;
    wire N__30808;
    wire N__30805;
    wire N__30802;
    wire N__30799;
    wire N__30796;
    wire N__30793;
    wire N__30792;
    wire N__30789;
    wire N__30786;
    wire N__30783;
    wire N__30780;
    wire N__30775;
    wire N__30774;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30757;
    wire N__30754;
    wire N__30753;
    wire N__30748;
    wire N__30745;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30724;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30712;
    wire N__30709;
    wire N__30706;
    wire N__30703;
    wire N__30702;
    wire N__30701;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30669;
    wire N__30666;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30656;
    wire N__30653;
    wire N__30646;
    wire N__30643;
    wire N__30640;
    wire N__30639;
    wire N__30634;
    wire N__30633;
    wire N__30632;
    wire N__30631;
    wire N__30630;
    wire N__30629;
    wire N__30628;
    wire N__30627;
    wire N__30626;
    wire N__30625;
    wire N__30624;
    wire N__30623;
    wire N__30622;
    wire N__30619;
    wire N__30610;
    wire N__30609;
    wire N__30606;
    wire N__30605;
    wire N__30604;
    wire N__30603;
    wire N__30602;
    wire N__30599;
    wire N__30598;
    wire N__30589;
    wire N__30586;
    wire N__30583;
    wire N__30578;
    wire N__30575;
    wire N__30574;
    wire N__30573;
    wire N__30572;
    wire N__30571;
    wire N__30568;
    wire N__30567;
    wire N__30564;
    wire N__30561;
    wire N__30556;
    wire N__30553;
    wire N__30550;
    wire N__30547;
    wire N__30538;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30515;
    wire N__30512;
    wire N__30503;
    wire N__30498;
    wire N__30493;
    wire N__30490;
    wire N__30487;
    wire N__30482;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30442;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30417;
    wire N__30412;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30402;
    wire N__30399;
    wire N__30396;
    wire N__30393;
    wire N__30390;
    wire N__30389;
    wire N__30388;
    wire N__30385;
    wire N__30382;
    wire N__30379;
    wire N__30376;
    wire N__30373;
    wire N__30364;
    wire N__30361;
    wire N__30358;
    wire N__30357;
    wire N__30354;
    wire N__30353;
    wire N__30350;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30340;
    wire N__30337;
    wire N__30336;
    wire N__30335;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30316;
    wire N__30307;
    wire N__30306;
    wire N__30303;
    wire N__30302;
    wire N__30301;
    wire N__30300;
    wire N__30299;
    wire N__30298;
    wire N__30295;
    wire N__30282;
    wire N__30279;
    wire N__30276;
    wire N__30273;
    wire N__30270;
    wire N__30265;
    wire N__30262;
    wire N__30259;
    wire N__30258;
    wire N__30257;
    wire N__30256;
    wire N__30253;
    wire N__30246;
    wire N__30241;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30174;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30135;
    wire N__30132;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30118;
    wire N__30117;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30085;
    wire N__30084;
    wire N__30081;
    wire N__30078;
    wire N__30073;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30060;
    wire N__30059;
    wire N__30052;
    wire N__30049;
    wire N__30046;
    wire N__30043;
    wire N__30042;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30028;
    wire N__30027;
    wire N__30024;
    wire N__30021;
    wire N__30016;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29980;
    wire N__29977;
    wire N__29974;
    wire N__29971;
    wire N__29968;
    wire N__29967;
    wire N__29964;
    wire N__29963;
    wire N__29960;
    wire N__29957;
    wire N__29954;
    wire N__29951;
    wire N__29944;
    wire N__29941;
    wire N__29940;
    wire N__29937;
    wire N__29934;
    wire N__29931;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29913;
    wire N__29910;
    wire N__29909;
    wire N__29906;
    wire N__29905;
    wire N__29900;
    wire N__29897;
    wire N__29894;
    wire N__29887;
    wire N__29884;
    wire N__29883;
    wire N__29880;
    wire N__29877;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29859;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29842;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29825;
    wire N__29818;
    wire N__29817;
    wire N__29814;
    wire N__29811;
    wire N__29810;
    wire N__29807;
    wire N__29804;
    wire N__29801;
    wire N__29798;
    wire N__29791;
    wire N__29788;
    wire N__29785;
    wire N__29782;
    wire N__29779;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29752;
    wire N__29749;
    wire N__29746;
    wire N__29745;
    wire N__29742;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29722;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29710;
    wire N__29707;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29697;
    wire N__29694;
    wire N__29691;
    wire N__29686;
    wire N__29685;
    wire N__29682;
    wire N__29679;
    wire N__29678;
    wire N__29673;
    wire N__29672;
    wire N__29671;
    wire N__29670;
    wire N__29667;
    wire N__29664;
    wire N__29661;
    wire N__29660;
    wire N__29659;
    wire N__29658;
    wire N__29655;
    wire N__29654;
    wire N__29653;
    wire N__29652;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29639;
    wire N__29638;
    wire N__29635;
    wire N__29634;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29620;
    wire N__29619;
    wire N__29616;
    wire N__29615;
    wire N__29612;
    wire N__29609;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29590;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29566;
    wire N__29553;
    wire N__29542;
    wire N__29539;
    wire N__29536;
    wire N__29535;
    wire N__29534;
    wire N__29533;
    wire N__29532;
    wire N__29529;
    wire N__29520;
    wire N__29515;
    wire N__29514;
    wire N__29513;
    wire N__29512;
    wire N__29511;
    wire N__29510;
    wire N__29507;
    wire N__29506;
    wire N__29505;
    wire N__29502;
    wire N__29493;
    wire N__29486;
    wire N__29479;
    wire N__29476;
    wire N__29475;
    wire N__29474;
    wire N__29473;
    wire N__29472;
    wire N__29471;
    wire N__29466;
    wire N__29457;
    wire N__29452;
    wire N__29449;
    wire N__29446;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29431;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29419;
    wire N__29416;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29404;
    wire N__29401;
    wire N__29398;
    wire N__29395;
    wire N__29392;
    wire N__29389;
    wire N__29386;
    wire N__29383;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29364;
    wire N__29363;
    wire N__29362;
    wire N__29355;
    wire N__29354;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29328;
    wire N__29325;
    wire N__29318;
    wire N__29315;
    wire N__29314;
    wire N__29311;
    wire N__29308;
    wire N__29305;
    wire N__29302;
    wire N__29293;
    wire N__29290;
    wire N__29287;
    wire N__29286;
    wire N__29285;
    wire N__29284;
    wire N__29281;
    wire N__29278;
    wire N__29277;
    wire N__29274;
    wire N__29273;
    wire N__29272;
    wire N__29269;
    wire N__29268;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29251;
    wire N__29250;
    wire N__29249;
    wire N__29248;
    wire N__29247;
    wire N__29246;
    wire N__29243;
    wire N__29240;
    wire N__29239;
    wire N__29238;
    wire N__29237;
    wire N__29236;
    wire N__29235;
    wire N__29228;
    wire N__29223;
    wire N__29222;
    wire N__29221;
    wire N__29218;
    wire N__29217;
    wire N__29216;
    wire N__29215;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29202;
    wire N__29201;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29191;
    wire N__29186;
    wire N__29183;
    wire N__29180;
    wire N__29175;
    wire N__29164;
    wire N__29147;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29119;
    wire N__29116;
    wire N__29113;
    wire N__29112;
    wire N__29111;
    wire N__29108;
    wire N__29103;
    wire N__29100;
    wire N__29099;
    wire N__29096;
    wire N__29095;
    wire N__29094;
    wire N__29093;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29085;
    wire N__29082;
    wire N__29079;
    wire N__29076;
    wire N__29073;
    wire N__29072;
    wire N__29071;
    wire N__29068;
    wire N__29063;
    wire N__29060;
    wire N__29055;
    wire N__29050;
    wire N__29047;
    wire N__29044;
    wire N__29037;
    wire N__29034;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28995;
    wire N__28994;
    wire N__28993;
    wire N__28992;
    wire N__28991;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28978;
    wire N__28975;
    wire N__28974;
    wire N__28973;
    wire N__28972;
    wire N__28971;
    wire N__28966;
    wire N__28963;
    wire N__28962;
    wire N__28959;
    wire N__28958;
    wire N__28957;
    wire N__28956;
    wire N__28955;
    wire N__28954;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28944;
    wire N__28941;
    wire N__28940;
    wire N__28937;
    wire N__28936;
    wire N__28935;
    wire N__28934;
    wire N__28931;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28918;
    wire N__28915;
    wire N__28910;
    wire N__28901;
    wire N__28896;
    wire N__28893;
    wire N__28888;
    wire N__28879;
    wire N__28876;
    wire N__28873;
    wire N__28866;
    wire N__28863;
    wire N__28856;
    wire N__28837;
    wire N__28836;
    wire N__28833;
    wire N__28832;
    wire N__28831;
    wire N__28830;
    wire N__28829;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28773;
    wire N__28762;
    wire N__28761;
    wire N__28756;
    wire N__28753;
    wire N__28752;
    wire N__28751;
    wire N__28748;
    wire N__28747;
    wire N__28746;
    wire N__28745;
    wire N__28744;
    wire N__28741;
    wire N__28740;
    wire N__28739;
    wire N__28736;
    wire N__28733;
    wire N__28732;
    wire N__28731;
    wire N__28728;
    wire N__28725;
    wire N__28722;
    wire N__28717;
    wire N__28712;
    wire N__28709;
    wire N__28708;
    wire N__28707;
    wire N__28706;
    wire N__28705;
    wire N__28702;
    wire N__28697;
    wire N__28692;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28678;
    wire N__28675;
    wire N__28674;
    wire N__28669;
    wire N__28668;
    wire N__28663;
    wire N__28654;
    wire N__28651;
    wire N__28648;
    wire N__28645;
    wire N__28642;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28625;
    wire N__28620;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28606;
    wire N__28597;
    wire N__28594;
    wire N__28593;
    wire N__28592;
    wire N__28591;
    wire N__28588;
    wire N__28583;
    wire N__28582;
    wire N__28581;
    wire N__28578;
    wire N__28577;
    wire N__28576;
    wire N__28575;
    wire N__28574;
    wire N__28573;
    wire N__28572;
    wire N__28567;
    wire N__28564;
    wire N__28561;
    wire N__28560;
    wire N__28559;
    wire N__28556;
    wire N__28553;
    wire N__28550;
    wire N__28549;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28529;
    wire N__28524;
    wire N__28519;
    wire N__28516;
    wire N__28511;
    wire N__28504;
    wire N__28501;
    wire N__28496;
    wire N__28489;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28462;
    wire N__28461;
    wire N__28460;
    wire N__28459;
    wire N__28458;
    wire N__28457;
    wire N__28456;
    wire N__28455;
    wire N__28454;
    wire N__28447;
    wire N__28440;
    wire N__28435;
    wire N__28434;
    wire N__28433;
    wire N__28430;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28413;
    wire N__28412;
    wire N__28409;
    wire N__28406;
    wire N__28405;
    wire N__28404;
    wire N__28403;
    wire N__28396;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28378;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28348;
    wire N__28347;
    wire N__28346;
    wire N__28345;
    wire N__28344;
    wire N__28343;
    wire N__28340;
    wire N__28337;
    wire N__28336;
    wire N__28333;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28322;
    wire N__28317;
    wire N__28312;
    wire N__28311;
    wire N__28310;
    wire N__28309;
    wire N__28308;
    wire N__28307;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28293;
    wire N__28292;
    wire N__28291;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28277;
    wire N__28276;
    wire N__28273;
    wire N__28270;
    wire N__28265;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28253;
    wire N__28252;
    wire N__28249;
    wire N__28244;
    wire N__28241;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28223;
    wire N__28220;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28203;
    wire N__28196;
    wire N__28193;
    wire N__28188;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28168;
    wire N__28167;
    wire N__28166;
    wire N__28165;
    wire N__28164;
    wire N__28163;
    wire N__28160;
    wire N__28159;
    wire N__28158;
    wire N__28157;
    wire N__28154;
    wire N__28153;
    wire N__28148;
    wire N__28143;
    wire N__28142;
    wire N__28141;
    wire N__28140;
    wire N__28137;
    wire N__28130;
    wire N__28127;
    wire N__28124;
    wire N__28119;
    wire N__28118;
    wire N__28117;
    wire N__28114;
    wire N__28111;
    wire N__28108;
    wire N__28107;
    wire N__28102;
    wire N__28097;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28068;
    wire N__28063;
    wire N__28056;
    wire N__28053;
    wire N__28048;
    wire N__28039;
    wire N__28036;
    wire N__28033;
    wire N__28032;
    wire N__28031;
    wire N__28030;
    wire N__28029;
    wire N__28028;
    wire N__28025;
    wire N__28024;
    wire N__28021;
    wire N__28020;
    wire N__28019;
    wire N__28018;
    wire N__28017;
    wire N__28016;
    wire N__28015;
    wire N__28014;
    wire N__28013;
    wire N__28012;
    wire N__28011;
    wire N__28010;
    wire N__28003;
    wire N__28000;
    wire N__27999;
    wire N__27996;
    wire N__27991;
    wire N__27988;
    wire N__27987;
    wire N__27986;
    wire N__27985;
    wire N__27982;
    wire N__27975;
    wire N__27972;
    wire N__27969;
    wire N__27966;
    wire N__27965;
    wire N__27958;
    wire N__27957;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27942;
    wire N__27939;
    wire N__27936;
    wire N__27931;
    wire N__27928;
    wire N__27921;
    wire N__27916;
    wire N__27913;
    wire N__27912;
    wire N__27909;
    wire N__27906;
    wire N__27897;
    wire N__27890;
    wire N__27883;
    wire N__27880;
    wire N__27877;
    wire N__27862;
    wire N__27859;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27843;
    wire N__27840;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27826;
    wire N__27823;
    wire N__27820;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27780;
    wire N__27779;
    wire N__27778;
    wire N__27777;
    wire N__27776;
    wire N__27773;
    wire N__27772;
    wire N__27771;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27760;
    wire N__27759;
    wire N__27758;
    wire N__27755;
    wire N__27754;
    wire N__27753;
    wire N__27752;
    wire N__27751;
    wire N__27750;
    wire N__27747;
    wire N__27742;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27728;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27699;
    wire N__27696;
    wire N__27695;
    wire N__27694;
    wire N__27693;
    wire N__27692;
    wire N__27689;
    wire N__27686;
    wire N__27681;
    wire N__27676;
    wire N__27667;
    wire N__27664;
    wire N__27661;
    wire N__27654;
    wire N__27645;
    wire N__27642;
    wire N__27637;
    wire N__27628;
    wire N__27625;
    wire N__27624;
    wire N__27621;
    wire N__27620;
    wire N__27619;
    wire N__27618;
    wire N__27617;
    wire N__27614;
    wire N__27611;
    wire N__27610;
    wire N__27607;
    wire N__27606;
    wire N__27605;
    wire N__27604;
    wire N__27603;
    wire N__27600;
    wire N__27599;
    wire N__27598;
    wire N__27597;
    wire N__27596;
    wire N__27595;
    wire N__27594;
    wire N__27593;
    wire N__27588;
    wire N__27587;
    wire N__27582;
    wire N__27575;
    wire N__27570;
    wire N__27567;
    wire N__27564;
    wire N__27561;
    wire N__27558;
    wire N__27551;
    wire N__27550;
    wire N__27549;
    wire N__27548;
    wire N__27547;
    wire N__27546;
    wire N__27545;
    wire N__27540;
    wire N__27537;
    wire N__27536;
    wire N__27535;
    wire N__27532;
    wire N__27529;
    wire N__27524;
    wire N__27521;
    wire N__27514;
    wire N__27511;
    wire N__27504;
    wire N__27499;
    wire N__27496;
    wire N__27493;
    wire N__27490;
    wire N__27485;
    wire N__27482;
    wire N__27467;
    wire N__27464;
    wire N__27451;
    wire N__27450;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27435;
    wire N__27432;
    wire N__27429;
    wire N__27428;
    wire N__27427;
    wire N__27426;
    wire N__27423;
    wire N__27418;
    wire N__27417;
    wire N__27414;
    wire N__27413;
    wire N__27410;
    wire N__27409;
    wire N__27408;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27391;
    wire N__27390;
    wire N__27389;
    wire N__27386;
    wire N__27383;
    wire N__27382;
    wire N__27379;
    wire N__27374;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27346;
    wire N__27331;
    wire N__27330;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27318;
    wire N__27317;
    wire N__27316;
    wire N__27315;
    wire N__27314;
    wire N__27313;
    wire N__27312;
    wire N__27311;
    wire N__27308;
    wire N__27307;
    wire N__27306;
    wire N__27305;
    wire N__27304;
    wire N__27303;
    wire N__27302;
    wire N__27297;
    wire N__27296;
    wire N__27295;
    wire N__27294;
    wire N__27293;
    wire N__27292;
    wire N__27289;
    wire N__27284;
    wire N__27279;
    wire N__27276;
    wire N__27275;
    wire N__27274;
    wire N__27271;
    wire N__27266;
    wire N__27263;
    wire N__27262;
    wire N__27259;
    wire N__27258;
    wire N__27257;
    wire N__27252;
    wire N__27249;
    wire N__27240;
    wire N__27237;
    wire N__27236;
    wire N__27235;
    wire N__27234;
    wire N__27233;
    wire N__27232;
    wire N__27231;
    wire N__27230;
    wire N__27229;
    wire N__27228;
    wire N__27221;
    wire N__27218;
    wire N__27213;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27195;
    wire N__27188;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27168;
    wire N__27163;
    wire N__27160;
    wire N__27153;
    wire N__27148;
    wire N__27141;
    wire N__27124;
    wire N__27121;
    wire N__27118;
    wire N__27115;
    wire N__27112;
    wire N__27109;
    wire N__27108;
    wire N__27107;
    wire N__27104;
    wire N__27103;
    wire N__27098;
    wire N__27093;
    wire N__27092;
    wire N__27091;
    wire N__27090;
    wire N__27089;
    wire N__27088;
    wire N__27087;
    wire N__27084;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27071;
    wire N__27070;
    wire N__27065;
    wire N__27062;
    wire N__27053;
    wire N__27050;
    wire N__27045;
    wire N__27034;
    wire N__27031;
    wire N__27030;
    wire N__27029;
    wire N__27028;
    wire N__27027;
    wire N__27026;
    wire N__27025;
    wire N__27022;
    wire N__27021;
    wire N__27016;
    wire N__27013;
    wire N__27008;
    wire N__27005;
    wire N__27004;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26990;
    wire N__26987;
    wire N__26984;
    wire N__26971;
    wire N__26968;
    wire N__26965;
    wire N__26964;
    wire N__26961;
    wire N__26960;
    wire N__26959;
    wire N__26956;
    wire N__26955;
    wire N__26954;
    wire N__26951;
    wire N__26946;
    wire N__26943;
    wire N__26942;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26927;
    wire N__26926;
    wire N__26925;
    wire N__26924;
    wire N__26923;
    wire N__26920;
    wire N__26917;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26899;
    wire N__26896;
    wire N__26881;
    wire N__26880;
    wire N__26879;
    wire N__26878;
    wire N__26877;
    wire N__26874;
    wire N__26873;
    wire N__26868;
    wire N__26867;
    wire N__26866;
    wire N__26863;
    wire N__26860;
    wire N__26855;
    wire N__26852;
    wire N__26851;
    wire N__26850;
    wire N__26849;
    wire N__26848;
    wire N__26845;
    wire N__26844;
    wire N__26843;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26831;
    wire N__26828;
    wire N__26827;
    wire N__26822;
    wire N__26811;
    wire N__26806;
    wire N__26801;
    wire N__26798;
    wire N__26795;
    wire N__26782;
    wire N__26781;
    wire N__26780;
    wire N__26779;
    wire N__26776;
    wire N__26773;
    wire N__26770;
    wire N__26767;
    wire N__26766;
    wire N__26765;
    wire N__26764;
    wire N__26761;
    wire N__26758;
    wire N__26757;
    wire N__26754;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26732;
    wire N__26729;
    wire N__26724;
    wire N__26721;
    wire N__26718;
    wire N__26713;
    wire N__26708;
    wire N__26703;
    wire N__26692;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26668;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26656;
    wire N__26653;
    wire N__26650;
    wire N__26649;
    wire N__26646;
    wire N__26643;
    wire N__26642;
    wire N__26639;
    wire N__26638;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26610;
    wire N__26607;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26597;
    wire N__26594;
    wire N__26587;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26566;
    wire N__26563;
    wire N__26560;
    wire N__26559;
    wire N__26556;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26536;
    wire N__26535;
    wire N__26532;
    wire N__26531;
    wire N__26528;
    wire N__26525;
    wire N__26522;
    wire N__26519;
    wire N__26518;
    wire N__26517;
    wire N__26512;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26494;
    wire N__26491;
    wire N__26490;
    wire N__26489;
    wire N__26488;
    wire N__26487;
    wire N__26486;
    wire N__26485;
    wire N__26484;
    wire N__26483;
    wire N__26482;
    wire N__26481;
    wire N__26480;
    wire N__26479;
    wire N__26470;
    wire N__26465;
    wire N__26464;
    wire N__26463;
    wire N__26462;
    wire N__26455;
    wire N__26446;
    wire N__26441;
    wire N__26440;
    wire N__26433;
    wire N__26428;
    wire N__26425;
    wire N__26422;
    wire N__26413;
    wire N__26410;
    wire N__26407;
    wire N__26404;
    wire N__26403;
    wire N__26400;
    wire N__26397;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26380;
    wire N__26379;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26329;
    wire N__26328;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26314;
    wire N__26311;
    wire N__26308;
    wire N__26307;
    wire N__26306;
    wire N__26305;
    wire N__26302;
    wire N__26301;
    wire N__26298;
    wire N__26289;
    wire N__26284;
    wire N__26283;
    wire N__26282;
    wire N__26279;
    wire N__26274;
    wire N__26269;
    wire N__26266;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26241;
    wire N__26236;
    wire N__26235;
    wire N__26234;
    wire N__26233;
    wire N__26232;
    wire N__26231;
    wire N__26230;
    wire N__26225;
    wire N__26224;
    wire N__26223;
    wire N__26220;
    wire N__26219;
    wire N__26216;
    wire N__26215;
    wire N__26214;
    wire N__26213;
    wire N__26212;
    wire N__26211;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26203;
    wire N__26200;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26190;
    wire N__26189;
    wire N__26188;
    wire N__26187;
    wire N__26184;
    wire N__26181;
    wire N__26180;
    wire N__26179;
    wire N__26178;
    wire N__26175;
    wire N__26168;
    wire N__26163;
    wire N__26160;
    wire N__26157;
    wire N__26148;
    wire N__26145;
    wire N__26142;
    wire N__26139;
    wire N__26134;
    wire N__26131;
    wire N__26126;
    wire N__26119;
    wire N__26112;
    wire N__26105;
    wire N__26086;
    wire N__26085;
    wire N__26080;
    wire N__26077;
    wire N__26074;
    wire N__26071;
    wire N__26070;
    wire N__26067;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26047;
    wire N__26044;
    wire N__26043;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26025;
    wire N__26022;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26002;
    wire N__26001;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25983;
    wire N__25980;
    wire N__25979;
    wire N__25976;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25960;
    wire N__25959;
    wire N__25954;
    wire N__25951;
    wire N__25948;
    wire N__25945;
    wire N__25942;
    wire N__25939;
    wire N__25936;
    wire N__25933;
    wire N__25930;
    wire N__25927;
    wire N__25924;
    wire N__25921;
    wire N__25920;
    wire N__25919;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25899;
    wire N__25894;
    wire N__25893;
    wire N__25890;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25870;
    wire N__25867;
    wire N__25866;
    wire N__25863;
    wire N__25862;
    wire N__25859;
    wire N__25856;
    wire N__25853;
    wire N__25846;
    wire N__25843;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25826;
    wire N__25819;
    wire N__25816;
    wire N__25815;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25789;
    wire N__25788;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25765;
    wire N__25762;
    wire N__25759;
    wire N__25758;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25738;
    wire N__25735;
    wire N__25732;
    wire N__25731;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25711;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25701;
    wire N__25700;
    wire N__25697;
    wire N__25696;
    wire N__25693;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25663;
    wire N__25662;
    wire N__25657;
    wire N__25656;
    wire N__25655;
    wire N__25654;
    wire N__25653;
    wire N__25652;
    wire N__25649;
    wire N__25646;
    wire N__25637;
    wire N__25634;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25620;
    wire N__25617;
    wire N__25616;
    wire N__25613;
    wire N__25610;
    wire N__25607;
    wire N__25604;
    wire N__25597;
    wire N__25596;
    wire N__25595;
    wire N__25594;
    wire N__25591;
    wire N__25590;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25571;
    wire N__25570;
    wire N__25567;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25552;
    wire N__25551;
    wire N__25550;
    wire N__25549;
    wire N__25548;
    wire N__25545;
    wire N__25540;
    wire N__25537;
    wire N__25534;
    wire N__25531;
    wire N__25528;
    wire N__25525;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25468;
    wire N__25467;
    wire N__25466;
    wire N__25465;
    wire N__25464;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25444;
    wire N__25443;
    wire N__25440;
    wire N__25439;
    wire N__25432;
    wire N__25429;
    wire N__25426;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25392;
    wire N__25391;
    wire N__25390;
    wire N__25389;
    wire N__25386;
    wire N__25385;
    wire N__25384;
    wire N__25383;
    wire N__25380;
    wire N__25379;
    wire N__25376;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25364;
    wire N__25361;
    wire N__25360;
    wire N__25355;
    wire N__25352;
    wire N__25347;
    wire N__25346;
    wire N__25341;
    wire N__25338;
    wire N__25337;
    wire N__25334;
    wire N__25333;
    wire N__25330;
    wire N__25327;
    wire N__25322;
    wire N__25319;
    wire N__25318;
    wire N__25315;
    wire N__25312;
    wire N__25309;
    wire N__25308;
    wire N__25305;
    wire N__25300;
    wire N__25293;
    wire N__25290;
    wire N__25285;
    wire N__25282;
    wire N__25279;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25243;
    wire N__25240;
    wire N__25237;
    wire N__25234;
    wire N__25231;
    wire N__25230;
    wire N__25225;
    wire N__25222;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25210;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25197;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25156;
    wire N__25153;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25141;
    wire N__25138;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25116;
    wire N__25111;
    wire N__25108;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25086;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25078;
    wire N__25077;
    wire N__25074;
    wire N__25073;
    wire N__25068;
    wire N__25067;
    wire N__25066;
    wire N__25065;
    wire N__25056;
    wire N__25055;
    wire N__25052;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25022;
    wire N__25019;
    wire N__25016;
    wire N__25013;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24976;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24954;
    wire N__24951;
    wire N__24948;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24918;
    wire N__24917;
    wire N__24912;
    wire N__24909;
    wire N__24904;
    wire N__24903;
    wire N__24898;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24883;
    wire N__24880;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24868;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24845;
    wire N__24838;
    wire N__24835;
    wire N__24832;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24820;
    wire N__24819;
    wire N__24818;
    wire N__24817;
    wire N__24816;
    wire N__24813;
    wire N__24812;
    wire N__24809;
    wire N__24808;
    wire N__24807;
    wire N__24802;
    wire N__24799;
    wire N__24796;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24782;
    wire N__24781;
    wire N__24780;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24754;
    wire N__24749;
    wire N__24746;
    wire N__24741;
    wire N__24724;
    wire N__24723;
    wire N__24722;
    wire N__24717;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24702;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24690;
    wire N__24689;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24677;
    wire N__24676;
    wire N__24675;
    wire N__24672;
    wire N__24669;
    wire N__24664;
    wire N__24661;
    wire N__24652;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24642;
    wire N__24639;
    wire N__24636;
    wire N__24633;
    wire N__24628;
    wire N__24625;
    wire N__24624;
    wire N__24621;
    wire N__24618;
    wire N__24615;
    wire N__24610;
    wire N__24607;
    wire N__24604;
    wire N__24601;
    wire N__24600;
    wire N__24595;
    wire N__24592;
    wire N__24589;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24564;
    wire N__24559;
    wire N__24556;
    wire N__24553;
    wire N__24552;
    wire N__24547;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24537;
    wire N__24534;
    wire N__24531;
    wire N__24526;
    wire N__24525;
    wire N__24522;
    wire N__24519;
    wire N__24516;
    wire N__24513;
    wire N__24512;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24500;
    wire N__24493;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24483;
    wire N__24482;
    wire N__24481;
    wire N__24478;
    wire N__24473;
    wire N__24470;
    wire N__24469;
    wire N__24468;
    wire N__24465;
    wire N__24464;
    wire N__24461;
    wire N__24456;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24441;
    wire N__24436;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24394;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24382;
    wire N__24379;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24365;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24353;
    wire N__24348;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24334;
    wire N__24331;
    wire N__24328;
    wire N__24325;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24317;
    wire N__24316;
    wire N__24315;
    wire N__24314;
    wire N__24313;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24301;
    wire N__24298;
    wire N__24295;
    wire N__24292;
    wire N__24291;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24279;
    wire N__24278;
    wire N__24277;
    wire N__24274;
    wire N__24269;
    wire N__24266;
    wire N__24259;
    wire N__24252;
    wire N__24247;
    wire N__24238;
    wire N__24237;
    wire N__24236;
    wire N__24233;
    wire N__24232;
    wire N__24231;
    wire N__24228;
    wire N__24227;
    wire N__24224;
    wire N__24221;
    wire N__24218;
    wire N__24215;
    wire N__24214;
    wire N__24211;
    wire N__24210;
    wire N__24207;
    wire N__24204;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24187;
    wire N__24184;
    wire N__24179;
    wire N__24176;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24164;
    wire N__24163;
    wire N__24162;
    wire N__24161;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24151;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24139;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24109;
    wire N__24106;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24096;
    wire N__24093;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24083;
    wire N__24082;
    wire N__24079;
    wire N__24076;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24062;
    wire N__24059;
    wire N__24058;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24046;
    wire N__24037;
    wire N__24034;
    wire N__24031;
    wire N__24028;
    wire N__24027;
    wire N__24022;
    wire N__24019;
    wire N__24018;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__24001;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23983;
    wire N__23980;
    wire N__23977;
    wire N__23974;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23949;
    wire N__23946;
    wire N__23943;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23922;
    wire N__23917;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23905;
    wire N__23904;
    wire N__23901;
    wire N__23898;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23874;
    wire N__23873;
    wire N__23872;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23854;
    wire N__23851;
    wire N__23848;
    wire N__23847;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23826;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23814;
    wire N__23811;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23796;
    wire N__23791;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23775;
    wire N__23770;
    wire N__23767;
    wire N__23764;
    wire N__23763;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23743;
    wire N__23740;
    wire N__23737;
    wire N__23734;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23722;
    wire N__23719;
    wire N__23718;
    wire N__23715;
    wire N__23714;
    wire N__23713;
    wire N__23710;
    wire N__23709;
    wire N__23702;
    wire N__23699;
    wire N__23696;
    wire N__23689;
    wire N__23688;
    wire N__23685;
    wire N__23684;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23619;
    wire N__23616;
    wire N__23615;
    wire N__23614;
    wire N__23613;
    wire N__23610;
    wire N__23603;
    wire N__23600;
    wire N__23593;
    wire N__23592;
    wire N__23589;
    wire N__23588;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23569;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23512;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23473;
    wire N__23470;
    wire N__23467;
    wire N__23466;
    wire N__23463;
    wire N__23460;
    wire N__23455;
    wire N__23452;
    wire N__23449;
    wire N__23448;
    wire N__23443;
    wire N__23440;
    wire N__23439;
    wire N__23436;
    wire N__23431;
    wire N__23428;
    wire N__23427;
    wire N__23424;
    wire N__23423;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23415;
    wire N__23414;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23398;
    wire N__23395;
    wire N__23386;
    wire N__23383;
    wire N__23382;
    wire N__23379;
    wire N__23378;
    wire N__23377;
    wire N__23376;
    wire N__23375;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23360;
    wire N__23355;
    wire N__23352;
    wire N__23347;
    wire N__23344;
    wire N__23343;
    wire N__23342;
    wire N__23341;
    wire N__23340;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23320;
    wire N__23317;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23286;
    wire N__23285;
    wire N__23284;
    wire N__23281;
    wire N__23278;
    wire N__23275;
    wire N__23272;
    wire N__23269;
    wire N__23264;
    wire N__23261;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23238;
    wire N__23235;
    wire N__23232;
    wire N__23231;
    wire N__23226;
    wire N__23223;
    wire N__23220;
    wire N__23217;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23205;
    wire N__23204;
    wire N__23201;
    wire N__23196;
    wire N__23193;
    wire N__23188;
    wire N__23185;
    wire N__23184;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23176;
    wire N__23175;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23157;
    wire N__23154;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23127;
    wire N__23122;
    wire N__23121;
    wire N__23118;
    wire N__23115;
    wire N__23114;
    wire N__23113;
    wire N__23112;
    wire N__23111;
    wire N__23110;
    wire N__23109;
    wire N__23108;
    wire N__23103;
    wire N__23100;
    wire N__23093;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23077;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23055;
    wire N__23054;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23044;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22983;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22971;
    wire N__22968;
    wire N__22965;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22941;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22929;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22894;
    wire N__22893;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22824;
    wire N__22819;
    wire N__22816;
    wire N__22813;
    wire N__22810;
    wire N__22809;
    wire N__22804;
    wire N__22801;
    wire N__22800;
    wire N__22797;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22785;
    wire N__22784;
    wire N__22783;
    wire N__22780;
    wire N__22779;
    wire N__22778;
    wire N__22777;
    wire N__22776;
    wire N__22775;
    wire N__22774;
    wire N__22773;
    wire N__22772;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22764;
    wire N__22763;
    wire N__22762;
    wire N__22761;
    wire N__22758;
    wire N__22755;
    wire N__22750;
    wire N__22743;
    wire N__22738;
    wire N__22735;
    wire N__22734;
    wire N__22733;
    wire N__22730;
    wire N__22729;
    wire N__22728;
    wire N__22727;
    wire N__22726;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22711;
    wire N__22708;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22692;
    wire N__22681;
    wire N__22674;
    wire N__22669;
    wire N__22664;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22593;
    wire N__22592;
    wire N__22589;
    wire N__22588;
    wire N__22587;
    wire N__22586;
    wire N__22585;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22577;
    wire N__22574;
    wire N__22567;
    wire N__22562;
    wire N__22557;
    wire N__22554;
    wire N__22553;
    wire N__22550;
    wire N__22547;
    wire N__22542;
    wire N__22537;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22497;
    wire N__22494;
    wire N__22493;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22401;
    wire N__22400;
    wire N__22397;
    wire N__22396;
    wire N__22393;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22366;
    wire N__22363;
    wire N__22362;
    wire N__22361;
    wire N__22360;
    wire N__22359;
    wire N__22356;
    wire N__22355;
    wire N__22354;
    wire N__22351;
    wire N__22350;
    wire N__22349;
    wire N__22348;
    wire N__22347;
    wire N__22346;
    wire N__22345;
    wire N__22342;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22324;
    wire N__22321;
    wire N__22318;
    wire N__22311;
    wire N__22310;
    wire N__22309;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22295;
    wire N__22288;
    wire N__22287;
    wire N__22284;
    wire N__22279;
    wire N__22276;
    wire N__22269;
    wire N__22266;
    wire N__22255;
    wire N__22254;
    wire N__22253;
    wire N__22250;
    wire N__22245;
    wire N__22244;
    wire N__22243;
    wire N__22242;
    wire N__22241;
    wire N__22240;
    wire N__22239;
    wire N__22238;
    wire N__22233;
    wire N__22228;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22199;
    wire N__22194;
    wire N__22191;
    wire N__22188;
    wire N__22181;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22072;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22024;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21988;
    wire N__21985;
    wire N__21982;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21958;
    wire N__21955;
    wire N__21952;
    wire N__21949;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21901;
    wire N__21898;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21855;
    wire N__21854;
    wire N__21853;
    wire N__21846;
    wire N__21843;
    wire N__21838;
    wire N__21835;
    wire N__21832;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21824;
    wire N__21823;
    wire N__21822;
    wire N__21819;
    wire N__21812;
    wire N__21809;
    wire N__21802;
    wire N__21801;
    wire N__21798;
    wire N__21797;
    wire N__21796;
    wire N__21793;
    wire N__21788;
    wire N__21785;
    wire N__21778;
    wire N__21775;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21745;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21721;
    wire N__21718;
    wire N__21717;
    wire N__21714;
    wire N__21713;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21627;
    wire N__21624;
    wire N__21623;
    wire N__21620;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21600;
    wire N__21599;
    wire N__21598;
    wire N__21597;
    wire N__21592;
    wire N__21591;
    wire N__21586;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21563;
    wire N__21560;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21492;
    wire N__21489;
    wire N__21486;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21453;
    wire N__21448;
    wire N__21445;
    wire N__21442;
    wire N__21441;
    wire N__21440;
    wire N__21437;
    wire N__21436;
    wire N__21435;
    wire N__21434;
    wire N__21433;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21417;
    wire N__21416;
    wire N__21415;
    wire N__21410;
    wire N__21409;
    wire N__21406;
    wire N__21399;
    wire N__21396;
    wire N__21395;
    wire N__21394;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21373;
    wire N__21368;
    wire N__21355;
    wire N__21354;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21336;
    wire N__21335;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21325;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21314;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21265;
    wire N__21264;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21246;
    wire N__21245;
    wire N__21244;
    wire N__21241;
    wire N__21240;
    wire N__21235;
    wire N__21232;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21224;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21214;
    wire N__21211;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21187;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21169;
    wire N__21166;
    wire N__21163;
    wire N__21160;
    wire N__21157;
    wire N__21156;
    wire N__21155;
    wire N__21154;
    wire N__21153;
    wire N__21150;
    wire N__21149;
    wire N__21144;
    wire N__21141;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21123;
    wire N__21120;
    wire N__21109;
    wire N__21106;
    wire N__21105;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21064;
    wire N__21063;
    wire N__21058;
    wire N__21055;
    wire N__21052;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21034;
    wire N__21031;
    wire N__21028;
    wire N__21025;
    wire N__21022;
    wire N__21019;
    wire N__21016;
    wire N__21015;
    wire N__21014;
    wire N__21013;
    wire N__21012;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20998;
    wire N__20997;
    wire N__20996;
    wire N__20995;
    wire N__20994;
    wire N__20989;
    wire N__20986;
    wire N__20983;
    wire N__20980;
    wire N__20977;
    wire N__20976;
    wire N__20971;
    wire N__20968;
    wire N__20963;
    wire N__20960;
    wire N__20959;
    wire N__20958;
    wire N__20957;
    wire N__20956;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20934;
    wire N__20925;
    wire N__20914;
    wire N__20911;
    wire N__20910;
    wire N__20905;
    wire N__20902;
    wire N__20899;
    wire N__20896;
    wire N__20893;
    wire N__20892;
    wire N__20891;
    wire N__20890;
    wire N__20887;
    wire N__20884;
    wire N__20881;
    wire N__20880;
    wire N__20877;
    wire N__20876;
    wire N__20875;
    wire N__20874;
    wire N__20871;
    wire N__20866;
    wire N__20863;
    wire N__20860;
    wire N__20853;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20815;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20800;
    wire N__20799;
    wire N__20798;
    wire N__20797;
    wire N__20788;
    wire N__20785;
    wire N__20782;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20742;
    wire N__20737;
    wire N__20734;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20722;
    wire N__20719;
    wire N__20718;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20700;
    wire N__20695;
    wire N__20692;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20680;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20662;
    wire N__20659;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20629;
    wire N__20628;
    wire N__20627;
    wire N__20626;
    wire N__20619;
    wire N__20616;
    wire N__20613;
    wire N__20610;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20593;
    wire N__20592;
    wire N__20589;
    wire N__20586;
    wire N__20581;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20557;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20544;
    wire N__20543;
    wire N__20542;
    wire N__20541;
    wire N__20540;
    wire N__20537;
    wire N__20526;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20493;
    wire N__20490;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20388;
    wire N__20385;
    wire N__20384;
    wire N__20383;
    wire N__20380;
    wire N__20375;
    wire N__20372;
    wire N__20365;
    wire N__20362;
    wire N__20359;
    wire N__20358;
    wire N__20353;
    wire N__20350;
    wire N__20347;
    wire N__20346;
    wire N__20345;
    wire N__20344;
    wire N__20343;
    wire N__20342;
    wire N__20341;
    wire N__20340;
    wire N__20339;
    wire N__20336;
    wire N__20331;
    wire N__20326;
    wire N__20319;
    wire N__20316;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20290;
    wire N__20287;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20274;
    wire N__20273;
    wire N__20272;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20264;
    wire N__20263;
    wire N__20256;
    wire N__20253;
    wire N__20248;
    wire N__20245;
    wire N__20236;
    wire N__20233;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20221;
    wire N__20218;
    wire N__20215;
    wire N__20212;
    wire N__20209;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20176;
    wire N__20175;
    wire N__20172;
    wire N__20171;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20157;
    wire N__20154;
    wire N__20153;
    wire N__20150;
    wire N__20149;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20137;
    wire N__20134;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20118;
    wire N__20115;
    wire N__20114;
    wire N__20111;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20097;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20080;
    wire N__20077;
    wire N__20076;
    wire N__20073;
    wire N__20070;
    wire N__20069;
    wire N__20068;
    wire N__20065;
    wire N__20060;
    wire N__20057;
    wire N__20050;
    wire N__20049;
    wire N__20046;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20038;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20011;
    wire N__20008;
    wire N__20007;
    wire N__20004;
    wire N__20001;
    wire N__20000;
    wire N__19999;
    wire N__19996;
    wire N__19991;
    wire N__19988;
    wire N__19981;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19930;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19914;
    wire N__19911;
    wire N__19908;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19884;
    wire N__19881;
    wire N__19878;
    wire N__19877;
    wire N__19876;
    wire N__19873;
    wire N__19868;
    wire N__19865;
    wire N__19858;
    wire N__19855;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19825;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19813;
    wire N__19810;
    wire N__19807;
    wire N__19804;
    wire N__19801;
    wire N__19798;
    wire N__19797;
    wire N__19794;
    wire N__19793;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19761;
    wire N__19758;
    wire N__19757;
    wire N__19750;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19729;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19714;
    wire N__19711;
    wire N__19708;
    wire N__19705;
    wire N__19702;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19669;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire N__19641;
    wire N__19638;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19609;
    wire N__19606;
    wire N__19605;
    wire N__19602;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19590;
    wire N__19585;
    wire N__19582;
    wire N__19581;
    wire N__19580;
    wire N__19579;
    wire N__19576;
    wire N__19575;
    wire N__19574;
    wire N__19573;
    wire N__19572;
    wire N__19571;
    wire N__19570;
    wire N__19569;
    wire N__19568;
    wire N__19567;
    wire N__19566;
    wire N__19565;
    wire N__19564;
    wire N__19563;
    wire N__19562;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19542;
    wire N__19541;
    wire N__19532;
    wire N__19523;
    wire N__19520;
    wire N__19519;
    wire N__19518;
    wire N__19517;
    wire N__19516;
    wire N__19515;
    wire N__19508;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19481;
    wire N__19478;
    wire N__19473;
    wire N__19472;
    wire N__19471;
    wire N__19470;
    wire N__19469;
    wire N__19468;
    wire N__19467;
    wire N__19466;
    wire N__19459;
    wire N__19454;
    wire N__19439;
    wire N__19432;
    wire N__19431;
    wire N__19430;
    wire N__19429;
    wire N__19428;
    wire N__19423;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19407;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19344;
    wire N__19341;
    wire N__19340;
    wire N__19339;
    wire N__19338;
    wire N__19337;
    wire N__19334;
    wire N__19333;
    wire N__19332;
    wire N__19329;
    wire N__19328;
    wire N__19323;
    wire N__19320;
    wire N__19319;
    wire N__19318;
    wire N__19313;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19297;
    wire N__19292;
    wire N__19279;
    wire N__19276;
    wire N__19273;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19258;
    wire N__19255;
    wire N__19252;
    wire N__19249;
    wire N__19246;
    wire N__19243;
    wire N__19240;
    wire N__19239;
    wire N__19236;
    wire N__19231;
    wire N__19228;
    wire N__19227;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19201;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19183;
    wire N__19180;
    wire N__19177;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19155;
    wire N__19154;
    wire N__19151;
    wire N__19150;
    wire N__19147;
    wire N__19144;
    wire N__19143;
    wire N__19142;
    wire N__19141;
    wire N__19140;
    wire N__19139;
    wire N__19134;
    wire N__19125;
    wire N__19118;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19057;
    wire N__19054;
    wire N__19051;
    wire N__19048;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19011;
    wire N__19008;
    wire N__19005;
    wire N__19002;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18951;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18937;
    wire N__18934;
    wire N__18931;
    wire N__18928;
    wire N__18927;
    wire N__18926;
    wire N__18925;
    wire N__18922;
    wire N__18915;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18897;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18879;
    wire N__18874;
    wire N__18871;
    wire N__18868;
    wire N__18865;
    wire N__18862;
    wire N__18859;
    wire N__18858;
    wire N__18855;
    wire N__18852;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18832;
    wire N__18829;
    wire N__18826;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18807;
    wire N__18804;
    wire N__18801;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18784;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18772;
    wire N__18769;
    wire N__18766;
    wire N__18763;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18741;
    wire N__18738;
    wire N__18735;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18694;
    wire N__18691;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18672;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18655;
    wire N__18652;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18622;
    wire N__18619;
    wire N__18618;
    wire N__18615;
    wire N__18614;
    wire N__18609;
    wire N__18606;
    wire N__18601;
    wire N__18598;
    wire N__18597;
    wire N__18594;
    wire N__18593;
    wire N__18590;
    wire N__18583;
    wire N__18580;
    wire N__18577;
    wire N__18574;
    wire N__18571;
    wire N__18568;
    wire N__18565;
    wire N__18562;
    wire N__18559;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18541;
    wire N__18538;
    wire N__18535;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18523;
    wire N__18520;
    wire N__18517;
    wire N__18514;
    wire N__18511;
    wire N__18508;
    wire N__18505;
    wire N__18502;
    wire N__18501;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18439;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18409;
    wire N__18408;
    wire N__18405;
    wire N__18404;
    wire N__18397;
    wire N__18394;
    wire N__18391;
    wire N__18388;
    wire N__18385;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18373;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18361;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18351;
    wire N__18350;
    wire N__18349;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18331;
    wire N__18328;
    wire N__18327;
    wire N__18326;
    wire N__18319;
    wire N__18316;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18304;
    wire N__18301;
    wire N__18298;
    wire N__18295;
    wire N__18292;
    wire N__18289;
    wire N__18286;
    wire N__18283;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18259;
    wire N__18256;
    wire N__18253;
    wire N__18250;
    wire N__18247;
    wire N__18244;
    wire N__18241;
    wire N__18238;
    wire N__18235;
    wire N__18234;
    wire N__18231;
    wire N__18230;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18208;
    wire N__18205;
    wire N__18202;
    wire N__18199;
    wire N__18196;
    wire N__18193;
    wire N__18190;
    wire N__18189;
    wire N__18186;
    wire N__18185;
    wire N__18178;
    wire N__18175;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18163;
    wire N__18162;
    wire N__18159;
    wire N__18158;
    wire N__18157;
    wire N__18156;
    wire N__18155;
    wire N__18154;
    wire N__18153;
    wire N__18152;
    wire N__18151;
    wire N__18144;
    wire N__18143;
    wire N__18140;
    wire N__18139;
    wire N__18138;
    wire N__18137;
    wire N__18136;
    wire N__18135;
    wire N__18134;
    wire N__18133;
    wire N__18132;
    wire N__18131;
    wire N__18130;
    wire N__18127;
    wire N__18120;
    wire N__18115;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18103;
    wire N__18102;
    wire N__18101;
    wire N__18100;
    wire N__18097;
    wire N__18094;
    wire N__18083;
    wire N__18078;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18057;
    wire N__18050;
    wire N__18047;
    wire N__18042;
    wire N__18039;
    wire N__18038;
    wire N__18037;
    wire N__18034;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18018;
    wire N__18011;
    wire N__18008;
    wire N__17999;
    wire N__17986;
    wire N__17983;
    wire N__17980;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17965;
    wire N__17962;
    wire N__17959;
    wire N__17958;
    wire N__17955;
    wire N__17954;
    wire N__17953;
    wire N__17952;
    wire N__17949;
    wire N__17944;
    wire N__17941;
    wire N__17938;
    wire N__17929;
    wire N__17926;
    wire N__17923;
    wire N__17920;
    wire N__17917;
    wire N__17914;
    wire N__17911;
    wire N__17910;
    wire N__17907;
    wire N__17904;
    wire N__17901;
    wire N__17898;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17883;
    wire N__17878;
    wire N__17875;
    wire N__17872;
    wire N__17869;
    wire N__17866;
    wire N__17863;
    wire N__17862;
    wire N__17859;
    wire N__17856;
    wire N__17853;
    wire N__17852;
    wire N__17849;
    wire N__17846;
    wire N__17845;
    wire N__17842;
    wire N__17837;
    wire N__17832;
    wire N__17827;
    wire N__17824;
    wire N__17821;
    wire N__17818;
    wire N__17815;
    wire N__17812;
    wire N__17811;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17799;
    wire N__17796;
    wire N__17793;
    wire N__17790;
    wire N__17787;
    wire N__17784;
    wire N__17781;
    wire N__17776;
    wire N__17773;
    wire N__17772;
    wire N__17769;
    wire N__17766;
    wire N__17761;
    wire N__17758;
    wire N__17755;
    wire N__17752;
    wire N__17751;
    wire N__17746;
    wire N__17743;
    wire N__17740;
    wire N__17737;
    wire N__17734;
    wire N__17733;
    wire N__17728;
    wire N__17725;
    wire N__17722;
    wire N__17719;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17692;
    wire N__17689;
    wire N__17686;
    wire N__17683;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17673;
    wire N__17672;
    wire N__17671;
    wire N__17662;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17640;
    wire N__17637;
    wire N__17634;
    wire N__17629;
    wire N__17626;
    wire N__17625;
    wire N__17622;
    wire N__17619;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17605;
    wire N__17604;
    wire N__17599;
    wire N__17596;
    wire N__17595;
    wire N__17592;
    wire N__17589;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17575;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17565;
    wire N__17562;
    wire N__17559;
    wire N__17554;
    wire N__17551;
    wire N__17548;
    wire N__17545;
    wire N__17542;
    wire N__17539;
    wire N__17538;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17527;
    wire N__17526;
    wire N__17525;
    wire N__17524;
    wire N__17523;
    wire N__17520;
    wire N__17515;
    wire N__17512;
    wire N__17511;
    wire N__17508;
    wire N__17501;
    wire N__17500;
    wire N__17499;
    wire N__17496;
    wire N__17495;
    wire N__17494;
    wire N__17489;
    wire N__17486;
    wire N__17485;
    wire N__17484;
    wire N__17483;
    wire N__17482;
    wire N__17481;
    wire N__17480;
    wire N__17477;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17467;
    wire N__17466;
    wire N__17463;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17447;
    wire N__17438;
    wire N__17433;
    wire N__17430;
    wire N__17423;
    wire N__17418;
    wire N__17401;
    wire N__17398;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17373;
    wire N__17370;
    wire N__17367;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17341;
    wire N__17338;
    wire N__17335;
    wire N__17332;
    wire N__17329;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17307;
    wire N__17304;
    wire N__17301;
    wire N__17296;
    wire N__17295;
    wire N__17290;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17236;
    wire N__17233;
    wire N__17230;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17212;
    wire N__17209;
    wire N__17206;
    wire N__17205;
    wire N__17202;
    wire N__17201;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17187;
    wire N__17184;
    wire N__17183;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17161;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17092;
    wire N__17089;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17049;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17026;
    wire N__17023;
    wire N__17020;
    wire N__17017;
    wire N__17014;
    wire N__17011;
    wire N__17010;
    wire N__17005;
    wire N__17002;
    wire N__17001;
    wire N__16998;
    wire N__16995;
    wire N__16990;
    wire N__16987;
    wire N__16984;
    wire N__16981;
    wire N__16978;
    wire N__16975;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16962;
    wire N__16959;
    wire N__16956;
    wire N__16953;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16938;
    wire N__16933;
    wire N__16930;
    wire N__16927;
    wire N__16924;
    wire N__16923;
    wire N__16920;
    wire N__16917;
    wire N__16914;
    wire N__16911;
    wire N__16906;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16887;
    wire N__16884;
    wire N__16881;
    wire N__16876;
    wire N__16873;
    wire N__16870;
    wire N__16869;
    wire N__16866;
    wire N__16863;
    wire N__16860;
    wire N__16855;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16842;
    wire N__16837;
    wire N__16834;
    wire N__16831;
    wire N__16828;
    wire N__16825;
    wire N__16824;
    wire N__16819;
    wire N__16816;
    wire N__16813;
    wire N__16810;
    wire N__16807;
    wire N__16804;
    wire N__16801;
    wire N__16798;
    wire N__16795;
    wire N__16794;
    wire N__16789;
    wire N__16786;
    wire N__16783;
    wire N__16780;
    wire N__16777;
    wire N__16774;
    wire N__16771;
    wire N__16770;
    wire N__16765;
    wire N__16762;
    wire N__16759;
    wire N__16756;
    wire N__16753;
    wire N__16752;
    wire N__16749;
    wire N__16746;
    wire N__16743;
    wire N__16740;
    wire N__16735;
    wire N__16732;
    wire N__16731;
    wire N__16726;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16714;
    wire N__16713;
    wire N__16712;
    wire N__16709;
    wire N__16704;
    wire N__16701;
    wire N__16696;
    wire N__16693;
    wire N__16692;
    wire N__16691;
    wire N__16690;
    wire N__16687;
    wire N__16680;
    wire N__16677;
    wire N__16672;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16662;
    wire N__16657;
    wire N__16654;
    wire N__16651;
    wire N__16648;
    wire N__16645;
    wire N__16642;
    wire N__16641;
    wire N__16638;
    wire N__16635;
    wire N__16630;
    wire N__16627;
    wire N__16624;
    wire N__16621;
    wire N__16618;
    wire N__16617;
    wire N__16614;
    wire N__16613;
    wire N__16612;
    wire N__16611;
    wire N__16610;
    wire N__16607;
    wire N__16606;
    wire N__16605;
    wire N__16604;
    wire N__16603;
    wire N__16602;
    wire N__16601;
    wire N__16600;
    wire N__16599;
    wire N__16596;
    wire N__16595;
    wire N__16594;
    wire N__16593;
    wire N__16582;
    wire N__16573;
    wire N__16566;
    wire N__16565;
    wire N__16564;
    wire N__16561;
    wire N__16558;
    wire N__16551;
    wire N__16544;
    wire N__16543;
    wire N__16542;
    wire N__16535;
    wire N__16530;
    wire N__16527;
    wire N__16522;
    wire N__16513;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16489;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16479;
    wire N__16474;
    wire N__16471;
    wire N__16468;
    wire N__16467;
    wire N__16462;
    wire N__16459;
    wire N__16456;
    wire N__16453;
    wire N__16450;
    wire N__16447;
    wire N__16444;
    wire N__16441;
    wire N__16440;
    wire N__16439;
    wire N__16432;
    wire N__16431;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16421;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16405;
    wire N__16402;
    wire N__16399;
    wire N__16398;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16385;
    wire N__16378;
    wire N__16377;
    wire N__16372;
    wire N__16369;
    wire N__16366;
    wire N__16365;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16345;
    wire N__16342;
    wire N__16339;
    wire N__16336;
    wire N__16335;
    wire N__16334;
    wire N__16331;
    wire N__16326;
    wire N__16323;
    wire N__16318;
    wire N__16315;
    wire N__16314;
    wire N__16313;
    wire N__16310;
    wire N__16305;
    wire N__16302;
    wire N__16297;
    wire N__16296;
    wire N__16293;
    wire N__16290;
    wire N__16289;
    wire N__16286;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16270;
    wire N__16269;
    wire N__16268;
    wire N__16265;
    wire N__16260;
    wire N__16255;
    wire N__16254;
    wire N__16253;
    wire N__16248;
    wire N__16245;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16233;
    wire N__16232;
    wire N__16231;
    wire N__16228;
    wire N__16221;
    wire N__16218;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16200;
    wire N__16195;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16183;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16173;
    wire N__16168;
    wire N__16165;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16150;
    wire N__16147;
    wire N__16146;
    wire N__16143;
    wire N__16140;
    wire N__16137;
    wire N__16132;
    wire N__16129;
    wire N__16126;
    wire N__16125;
    wire N__16120;
    wire N__16117;
    wire N__16116;
    wire N__16113;
    wire N__16110;
    wire N__16107;
    wire N__16102;
    wire N__16101;
    wire N__16096;
    wire N__16093;
    wire N__16090;
    wire N__16087;
    wire N__16086;
    wire N__16083;
    wire N__16080;
    wire N__16075;
    wire N__16074;
    wire N__16069;
    wire N__16066;
    wire N__16063;
    wire N__16062;
    wire N__16059;
    wire N__16056;
    wire N__16051;
    wire N__16048;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16026;
    wire N__16023;
    wire N__16020;
    wire N__16015;
    wire N__16014;
    wire N__16009;
    wire N__16006;
    wire N__16003;
    wire N__16000;
    wire N__15997;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15985;
    wire N__15982;
    wire N__15981;
    wire N__15976;
    wire N__15973;
    wire N__15970;
    wire N__15969;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15952;
    wire N__15949;
    wire N__15948;
    wire N__15945;
    wire N__15942;
    wire N__15937;
    wire N__15936;
    wire N__15933;
    wire N__15930;
    wire N__15925;
    wire N__15922;
    wire N__15921;
    wire N__15918;
    wire N__15915;
    wire N__15910;
    wire N__15907;
    wire N__15906;
    wire N__15903;
    wire N__15900;
    wire N__15895;
    wire N__15892;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15880;
    wire N__15877;
    wire N__15876;
    wire N__15871;
    wire N__15868;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15858;
    wire N__15853;
    wire N__15850;
    wire N__15847;
    wire N__15844;
    wire N__15843;
    wire N__15840;
    wire N__15837;
    wire N__15832;
    wire N__15829;
    wire N__15828;
    wire N__15823;
    wire N__15820;
    wire N__15817;
    wire N__15814;
    wire N__15813;
    wire N__15810;
    wire N__15807;
    wire N__15804;
    wire N__15801;
    wire N__15796;
    wire N__15795;
    wire N__15790;
    wire N__15787;
    wire N__15784;
    wire N__15781;
    wire N__15780;
    wire N__15777;
    wire N__15774;
    wire N__15769;
    wire N__15768;
    wire N__15763;
    wire N__15760;
    wire N__15757;
    wire N__15756;
    wire N__15753;
    wire N__15750;
    wire N__15745;
    wire N__15744;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15720;
    wire N__15719;
    wire N__15718;
    wire N__15717;
    wire N__15716;
    wire N__15715;
    wire N__15714;
    wire N__15713;
    wire N__15712;
    wire N__15711;
    wire N__15710;
    wire N__15709;
    wire N__15708;
    wire N__15707;
    wire N__15706;
    wire N__15705;
    wire N__15704;
    wire N__15701;
    wire N__15696;
    wire N__15689;
    wire N__15680;
    wire N__15671;
    wire N__15662;
    wire N__15661;
    wire N__15660;
    wire N__15659;
    wire N__15658;
    wire N__15657;
    wire N__15656;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15638;
    wire N__15613;
    wire N__15610;
    wire N__15607;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15586;
    wire N__15585;
    wire N__15582;
    wire N__15579;
    wire N__15574;
    wire N__15573;
    wire N__15568;
    wire N__15565;
    wire N__15562;
    wire N__15561;
    wire N__15558;
    wire N__15555;
    wire N__15550;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15540;
    wire N__15535;
    wire N__15532;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15520;
    wire N__15519;
    wire N__15514;
    wire N__15511;
    wire N__15508;
    wire N__15505;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15493;
    wire N__15492;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15480;
    wire N__15477;
    wire N__15474;
    wire N__15469;
    wire N__15468;
    wire N__15463;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15427;
    wire N__15424;
    wire N__15421;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15403;
    wire N__15400;
    wire N__15397;
    wire N__15396;
    wire N__15391;
    wire N__15388;
    wire N__15385;
    wire N__15382;
    wire N__15381;
    wire N__15380;
    wire N__15379;
    wire N__15378;
    wire N__15377;
    wire N__15372;
    wire N__15369;
    wire N__15362;
    wire N__15355;
    wire N__15352;
    wire N__15349;
    wire N__15346;
    wire N__15345;
    wire N__15342;
    wire N__15339;
    wire N__15334;
    wire N__15333;
    wire N__15328;
    wire N__15325;
    wire N__15322;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15301;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15289;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15277;
    wire N__15274;
    wire N__15271;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15250;
    wire N__15247;
    wire N__15244;
    wire N__15241;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15229;
    wire N__15226;
    wire N__15223;
    wire N__15222;
    wire N__15221;
    wire N__15218;
    wire N__15213;
    wire N__15210;
    wire N__15205;
    wire N__15204;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15192;
    wire N__15189;
    wire N__15186;
    wire N__15183;
    wire N__15180;
    wire N__15175;
    wire N__15172;
    wire N__15171;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15159;
    wire N__15154;
    wire N__15151;
    wire N__15150;
    wire N__15147;
    wire N__15144;
    wire N__15139;
    wire N__15136;
    wire N__15133;
    wire N__15130;
    wire N__15127;
    wire N__15124;
    wire N__15121;
    wire N__15118;
    wire N__15115;
    wire N__15112;
    wire N__15109;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15088;
    wire N__15085;
    wire N__15082;
    wire N__15079;
    wire N__15078;
    wire N__15073;
    wire N__15070;
    wire N__15067;
    wire N__15066;
    wire N__15061;
    wire N__15058;
    wire N__15057;
    wire N__15052;
    wire N__15049;
    wire N__15046;
    wire N__15043;
    wire N__15040;
    wire N__15037;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15024;
    wire N__15019;
    wire N__15016;
    wire N__15013;
    wire N__15010;
    wire N__15007;
    wire N__15004;
    wire N__15001;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14980;
    wire N__14977;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14967;
    wire N__14962;
    wire N__14959;
    wire N__14956;
    wire N__14953;
    wire N__14950;
    wire N__14949;
    wire N__14946;
    wire N__14943;
    wire N__14940;
    wire N__14935;
    wire N__14934;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14917;
    wire N__14914;
    wire N__14911;
    wire N__14908;
    wire N__14907;
    wire N__14902;
    wire N__14899;
    wire N__14896;
    wire N__14893;
    wire N__14890;
    wire N__14887;
    wire N__14884;
    wire N__14883;
    wire N__14878;
    wire N__14875;
    wire N__14872;
    wire N__14869;
    wire N__14868;
    wire N__14865;
    wire N__14862;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14850;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14836;
    wire N__14833;
    wire N__14832;
    wire N__14829;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14815;
    wire N__14812;
    wire N__14811;
    wire N__14808;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14790;
    wire N__14785;
    wire N__14782;
    wire N__14779;
    wire N__14776;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14754;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14740;
    wire N__14737;
    wire N__14734;
    wire N__14731;
    wire N__14728;
    wire N__14725;
    wire N__14722;
    wire N__14719;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14707;
    wire N__14704;
    wire N__14701;
    wire N__14698;
    wire N__14695;
    wire N__14692;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14668;
    wire N__14665;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14607;
    wire N__14602;
    wire N__14599;
    wire N__14596;
    wire N__14593;
    wire N__14592;
    wire N__14587;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14577;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14535;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14514;
    wire N__14511;
    wire N__14508;
    wire N__14503;
    wire N__14502;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14490;
    wire N__14487;
    wire N__14484;
    wire N__14479;
    wire N__14476;
    wire N__14473;
    wire N__14472;
    wire N__14469;
    wire N__14466;
    wire N__14461;
    wire N__14460;
    wire N__14455;
    wire N__14452;
    wire N__14449;
    wire N__14446;
    wire N__14445;
    wire N__14442;
    wire N__14439;
    wire N__14434;
    wire N__14431;
    wire N__14428;
    wire N__14425;
    wire N__14422;
    wire N__14419;
    wire N__14416;
    wire VCCG0;
    wire GNDG0;
    wire \b2v_inst16.count_4_3 ;
    wire \b2v_inst16.count_4_5 ;
    wire bfn_1_2_0_;
    wire \b2v_inst16.un4_count_1_cry_1 ;
    wire \b2v_inst16.countZ0Z_3 ;
    wire \b2v_inst16.count_rst_8 ;
    wire \b2v_inst16.un4_count_1_cry_2_cZ0 ;
    wire \b2v_inst16.countZ0Z_4 ;
    wire \b2v_inst16.un4_count_1_cry_3 ;
    wire \b2v_inst16.countZ0Z_5 ;
    wire \b2v_inst16.count_rst_10 ;
    wire \b2v_inst16.un4_count_1_cry_4 ;
    wire \b2v_inst16.un4_count_1_cry_5 ;
    wire \b2v_inst16.countZ0Z_7 ;
    wire \b2v_inst16.un4_count_1_cry_6 ;
    wire \b2v_inst16.un4_count_1_cry_7 ;
    wire \b2v_inst16.un4_count_1_cry_8 ;
    wire bfn_1_3_0_;
    wire \b2v_inst16.un4_count_1_cry_9 ;
    wire \b2v_inst16.un4_count_1_cry_10_cZ0 ;
    wire \b2v_inst16.un4_count_1_cry_11 ;
    wire \b2v_inst16.un4_count_1_cry_12 ;
    wire \b2v_inst16.un4_count_1_cry_13 ;
    wire \b2v_inst16.un4_count_1_cry_14 ;
    wire \b2v_inst16.count_rst_7 ;
    wire \b2v_inst16.count_4_2 ;
    wire \b2v_inst16.count_rst_1 ;
    wire \b2v_inst16.count_4_12 ;
    wire \b2v_inst16.count_rst_0 ;
    wire \b2v_inst16.count_4_11 ;
    wire \b2v_inst16.count_rst_11 ;
    wire \b2v_inst16.count_4_6 ;
    wire \b2v_inst200.un25_clk_100khz_12_cascade_ ;
    wire \b2v_inst200.count_RNIC03N_3Z0Z_0_cascade_ ;
    wire \b2v_inst200.count_RNI_0_0_cascade_ ;
    wire \b2v_inst200.count_2_11 ;
    wire \b2v_inst200.count_2_10 ;
    wire \b2v_inst200.count_2_8 ;
    wire \b2v_inst200.count_2_0 ;
    wire \b2v_inst200.countZ0Z_0_cascade_ ;
    wire \b2v_inst200.un25_clk_100khz_13 ;
    wire \b2v_inst200.count_2_6 ;
    wire \b2v_inst200.count_2_14 ;
    wire \b2v_inst200.un25_clk_100khz_10 ;
    wire \b2v_inst200.count_2_3 ;
    wire \b2v_inst200.count_2_4 ;
    wire \b2v_inst200.count_2_5 ;
    wire \b2v_inst200.count_2_9 ;
    wire \b2v_inst200.countZ0Z_9_cascade_ ;
    wire \b2v_inst200.un25_clk_100khz_9 ;
    wire \b2v_inst200.count_2_12 ;
    wire \b2v_inst200.count_2_13 ;
    wire bfn_1_9_0_;
    wire \b2v_inst11.un1_count_clk_2_cry_1 ;
    wire \b2v_inst11.un1_count_clk_2_cry_2 ;
    wire \b2v_inst11.un1_count_clk_2_cry_3 ;
    wire \b2v_inst11.un1_count_clk_2_cry_4 ;
    wire \b2v_inst11.un1_count_clk_2_cry_5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_6 ;
    wire \b2v_inst11.un1_count_clk_2_cry_7_cZ0 ;
    wire \b2v_inst11.un1_count_clk_2_cry_8_cZ0 ;
    wire bfn_1_10_0_;
    wire \b2v_inst11.un1_count_clk_2_cry_9_cZ0 ;
    wire \b2v_inst11.un1_count_clk_2_cry_10_cZ0 ;
    wire \b2v_inst11.un1_count_clk_2_cry_11 ;
    wire \b2v_inst11.un1_count_clk_2_cry_12 ;
    wire \b2v_inst11.un1_count_clk_2_cry_13 ;
    wire \b2v_inst11.un1_count_clk_2_cry_14 ;
    wire \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5 ;
    wire \b2v_inst11.count_clk_0_5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0 ;
    wire \b2v_inst11.count_clk_0_15 ;
    wire \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ;
    wire \b2v_inst11.count_clk_0_6 ;
    wire \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5 ;
    wire \b2v_inst11.count_clk_0_8 ;
    wire \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5 ;
    wire \b2v_inst11.count_clk_0_7 ;
    wire \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5 ;
    wire \b2v_inst11.count_clk_0_9 ;
    wire \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5 ;
    wire \b2v_inst11.count_clk_0_4 ;
    wire \b2v_inst11.count_off_1_2 ;
    wire \b2v_inst11.count_offZ0Z_2 ;
    wire \b2v_inst11.count_off_1_2_cascade_ ;
    wire \b2v_inst11.un34_clk_100khz_1_cascade_ ;
    wire \b2v_inst11.un34_clk_100khz_0 ;
    wire \b2v_inst11.count_off_0_5 ;
    wire bfn_1_14_0_;
    wire \b2v_inst11.un3_count_off_1_axb_2 ;
    wire \b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152 ;
    wire \b2v_inst11.un3_count_off_1_cry_1 ;
    wire \b2v_inst11.un3_count_off_1_cry_2_cZ0 ;
    wire \b2v_inst11.un3_count_off_1_cry_3_cZ0 ;
    wire \b2v_inst11.count_offZ0Z_5 ;
    wire \b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882 ;
    wire \b2v_inst11.un3_count_off_1_cry_4_cZ0 ;
    wire \b2v_inst11.un3_count_off_1_axb_6 ;
    wire \b2v_inst11.un3_count_off_1_cry_5 ;
    wire \b2v_inst11.un3_count_off_1_cry_6 ;
    wire \b2v_inst11.un3_count_off_1_cry_7 ;
    wire \b2v_inst11.un3_count_off_1_cry_8 ;
    wire bfn_1_15_0_;
    wire \b2v_inst11.un3_count_off_1_cry_9 ;
    wire \b2v_inst11.un3_count_off_1_cry_10 ;
    wire \b2v_inst11.un3_count_off_1_cry_11 ;
    wire \b2v_inst11.un3_count_off_1_cry_12 ;
    wire \b2v_inst11.un3_count_off_1_cry_13 ;
    wire \b2v_inst11.un3_count_off_1_cry_14 ;
    wire \b2v_inst11.count_off_1_3_cascade_ ;
    wire \b2v_inst11.un3_count_off_1_axb_3 ;
    wire \b2v_inst11.count_offZ0Z_4 ;
    wire \b2v_inst11.count_off_1_3 ;
    wire \b2v_inst11.count_offZ0Z_4_cascade_ ;
    wire \b2v_inst11.un34_clk_100khz_2 ;
    wire \b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362 ;
    wire \b2v_inst11.count_offZ0Z_3 ;
    wire \b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672 ;
    wire \b2v_inst11.count_off_0_4 ;
    wire \b2v_inst11.count_off_0_14 ;
    wire \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5 ;
    wire \b2v_inst16.count_rst_12 ;
    wire \b2v_inst16.count_4_7 ;
    wire \b2v_inst16.count_rst_9 ;
    wire \b2v_inst16.count_4_4 ;
    wire \b2v_inst16.count_rst_6_cascade_ ;
    wire \b2v_inst16.count_rst_6 ;
    wire \b2v_inst16.countZ0Z_11 ;
    wire \b2v_inst16.countZ0Z_1_cascade_ ;
    wire \b2v_inst16.un4_count_1_axb_1 ;
    wire \b2v_inst16.count_4_1 ;
    wire \b2v_inst16.countZ0Z_2 ;
    wire \b2v_inst16.countZ0Z_6 ;
    wire \b2v_inst16.countZ0Z_12 ;
    wire \b2v_inst16.un13_clk_100khz_9 ;
    wire \b2v_inst16.un13_clk_100khz_8 ;
    wire \b2v_inst16.un13_clk_100khz_10_cascade_ ;
    wire \b2v_inst16.un13_clk_100khz_i_cascade_ ;
    wire \b2v_inst16.count_4_0 ;
    wire \b2v_inst16.count_rst_5_cascade_ ;
    wire \b2v_inst16.count_4_13 ;
    wire \b2v_inst16.count_rst_2 ;
    wire \b2v_inst16.countZ0Z_13 ;
    wire \b2v_inst16.countZ0Z_0 ;
    wire \b2v_inst16.countZ0Z_13_cascade_ ;
    wire \b2v_inst16.un13_clk_100khz_11 ;
    wire \b2v_inst16.countZ0Z_15 ;
    wire \b2v_inst16.count_rst_4 ;
    wire \b2v_inst16.count_4_15 ;
    wire \b2v_inst16.count_4_14 ;
    wire \b2v_inst16.count_rst_3 ;
    wire \b2v_inst16.countZ0Z_14 ;
    wire \b2v_inst200.count_2_15 ;
    wire \b2v_inst200.count_2_7 ;
    wire \b2v_inst200.un25_clk_100khz_11 ;
    wire \b2v_inst200.count_0_16 ;
    wire \b2v_inst200.count_0_17 ;
    wire \b2v_inst200.count_2_1 ;
    wire \b2v_inst200.count_2_2 ;
    wire \b2v_inst200.count_en_g ;
    wire \b2v_inst200.countZ0Z_0 ;
    wire \b2v_inst200.count_1_0 ;
    wire bfn_2_6_0_;
    wire \b2v_inst200.countZ0Z_1 ;
    wire \b2v_inst200.count_RNIC03N_5Z0Z_0 ;
    wire \b2v_inst200.un2_count_1_cry_1_cy ;
    wire \b2v_inst200.countZ0Z_2 ;
    wire \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ;
    wire \b2v_inst200.un2_count_1_cry_1 ;
    wire \b2v_inst200.countZ0Z_3 ;
    wire \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0 ;
    wire \b2v_inst200.un2_count_1_cry_2 ;
    wire \b2v_inst200.countZ0Z_4 ;
    wire \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ;
    wire \b2v_inst200.un2_count_1_cry_3 ;
    wire \b2v_inst200.countZ0Z_5 ;
    wire \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ;
    wire \b2v_inst200.un2_count_1_cry_4 ;
    wire \b2v_inst200.countZ0Z_6 ;
    wire \b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0 ;
    wire \b2v_inst200.un2_count_1_cry_5 ;
    wire \b2v_inst200.countZ0Z_7 ;
    wire \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ;
    wire \b2v_inst200.un2_count_1_cry_6 ;
    wire \b2v_inst200.un2_count_1_cry_7 ;
    wire \b2v_inst200.countZ0Z_8 ;
    wire \b2v_inst200.un2_count_1_cry_7_c_RNIP33EZ0 ;
    wire bfn_2_7_0_;
    wire \b2v_inst200.countZ0Z_9 ;
    wire \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0 ;
    wire \b2v_inst200.un2_count_1_cry_8 ;
    wire \b2v_inst200.countZ0Z_10 ;
    wire \b2v_inst200.un2_count_1_cry_9_c_RNIR75EZ0 ;
    wire \b2v_inst200.un2_count_1_cry_9 ;
    wire \b2v_inst200.countZ0Z_11 ;
    wire \b2v_inst200.un2_count_1_cry_10_c_RNI3AZ0Z29 ;
    wire \b2v_inst200.un2_count_1_cry_10 ;
    wire \b2v_inst200.countZ0Z_12 ;
    wire \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39 ;
    wire \b2v_inst200.un2_count_1_cry_11 ;
    wire \b2v_inst200.countZ0Z_13 ;
    wire \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49 ;
    wire \b2v_inst200.un2_count_1_cry_12 ;
    wire \b2v_inst200.countZ0Z_14 ;
    wire \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59 ;
    wire \b2v_inst200.un2_count_1_cry_13 ;
    wire \b2v_inst200.countZ0Z_15 ;
    wire \b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69 ;
    wire \b2v_inst200.un2_count_1_cry_14 ;
    wire \b2v_inst200.un2_count_1_cry_15 ;
    wire \b2v_inst200.countZ0Z_16 ;
    wire \b2v_inst200.count_1_16 ;
    wire bfn_2_8_0_;
    wire \b2v_inst200.countZ0Z_17 ;
    wire \b2v_inst200.un2_count_1_cry_16 ;
    wire \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ;
    wire \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AAZ0 ;
    wire \b2v_inst11.count_clk_0_11 ;
    wire \b2v_inst11.count_clkZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_clk_0_0 ;
    wire \b2v_inst11.count_clk_0_10 ;
    wire \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5 ;
    wire \b2v_inst11.count_clkZ0Z_10 ;
    wire \b2v_inst11.count_clkZ0Z_11 ;
    wire \b2v_inst11.count_clkZ0Z_10_cascade_ ;
    wire \b2v_inst11.count_clkZ0Z_15 ;
    wire \b2v_inst11.un2_count_clk_17_0_o2_1_4_cascade_ ;
    wire \b2v_inst11.count_clkZ0Z_14 ;
    wire \b2v_inst11.count_clk_0_13 ;
    wire \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CAZ0 ;
    wire \b2v_inst11.count_clkZ0Z_13 ;
    wire \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DAZ0 ;
    wire \b2v_inst11.count_clk_0_14 ;
    wire \b2v_inst11.count_clk_en_cascade_ ;
    wire \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5 ;
    wire \b2v_inst11.count_clk_0_2 ;
    wire \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_ ;
    wire \b2v_inst11.N_373 ;
    wire \b2v_inst11.N_373_cascade_ ;
    wire \b2v_inst11.count_clkZ0Z_8 ;
    wire \b2v_inst11.count_clkZ0Z_6 ;
    wire \b2v_inst11.count_clkZ0Z_4 ;
    wire \b2v_inst11.count_clkZ0Z_2 ;
    wire \b2v_inst11.count_clkZ0Z_3 ;
    wire \b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_ ;
    wire \b2v_inst11.count_clkZ0Z_7 ;
    wire \b2v_inst11.count_clk_RNIZ0Z_3_cascade_ ;
    wire \b2v_inst11.count_clk_en_0 ;
    wire \b2v_inst11.count_clkZ0Z_12 ;
    wire \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BAZ0 ;
    wire \b2v_inst11.count_clk_0_12 ;
    wire \b2v_inst11.count_clk_RNI_0Z0Z_0 ;
    wire \b2v_inst11.count_clkZ0Z_0 ;
    wire \b2v_inst11.count_clk_0_1 ;
    wire \b2v_inst11.count_clk_RNIZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_clkZ0Z_1_cascade_ ;
    wire \b2v_inst11.count_clkZ0Z_5 ;
    wire \b2v_inst11.N_187 ;
    wire \b2v_inst11.count_clkZ0Z_9 ;
    wire \b2v_inst11.count_clkZ0Z_1 ;
    wire \b2v_inst11.count_clk_RNIZ0Z_5 ;
    wire \b2v_inst11.N_172 ;
    wire \b2v_inst11.N_421 ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_i_1 ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_0_cascade_ ;
    wire \b2v_inst11.func_state_RNICC5V2_0_1 ;
    wire \b2v_inst11.count_off_1_11_cascade_ ;
    wire \b2v_inst11.un3_count_off_1_axb_11 ;
    wire \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5 ;
    wire \b2v_inst11.un34_clk_100khz_12 ;
    wire \b2v_inst11.un34_clk_100khz_4_cascade_ ;
    wire \b2v_inst11.count_off_0_12 ;
    wire \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5 ;
    wire \b2v_inst11.count_offZ0Z_12 ;
    wire \b2v_inst11.count_off_1_11 ;
    wire \b2v_inst11.count_offZ0Z_11 ;
    wire \b2v_inst11.count_offZ0Z_12_cascade_ ;
    wire \b2v_inst11.un34_clk_100khz_5 ;
    wire \b2v_inst11.count_offZ0Z_6 ;
    wire \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2 ;
    wire \b2v_inst11.count_off_1_9 ;
    wire \b2v_inst11.count_off_1_9_cascade_ ;
    wire \b2v_inst11.count_offZ0Z_9 ;
    wire \b2v_inst11.un3_count_off_1_axb_9 ;
    wire \b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92 ;
    wire \b2v_inst11.count_off_1_6 ;
    wire \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2 ;
    wire \b2v_inst11.count_off_0_15 ;
    wire \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5 ;
    wire \b2v_inst11.count_offZ0Z_15 ;
    wire \b2v_inst11.count_offZ0Z_13 ;
    wire \b2v_inst11.count_offZ0Z_14 ;
    wire \b2v_inst11.count_offZ0Z_15_cascade_ ;
    wire \b2v_inst11.un34_clk_100khz_11 ;
    wire \b2v_inst11.count_off_0_8 ;
    wire \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2 ;
    wire \b2v_inst11.count_offZ0Z_8 ;
    wire \b2v_inst11.count_offZ0Z_8_cascade_ ;
    wire \b2v_inst11.un34_clk_100khz_3 ;
    wire \b2v_inst11.count_offZ0Z_7 ;
    wire \b2v_inst11.count_off_1_7 ;
    wire \b2v_inst11.un3_count_off_1_axb_7 ;
    wire bfn_4_1_0_;
    wire \b2v_inst11.mult1_un96_sum_cry_2 ;
    wire \b2v_inst11.mult1_un96_sum_cry_3 ;
    wire \b2v_inst11.mult1_un96_sum_cry_4 ;
    wire \b2v_inst11.mult1_un96_sum_cry_5 ;
    wire \b2v_inst11.mult1_un96_sum_cry_6 ;
    wire \b2v_inst11.mult1_un96_sum_cry_7 ;
    wire \b2v_inst11.mult1_un96_sum_s_8_cascade_ ;
    wire bfn_4_2_0_;
    wire \b2v_inst11.mult1_un89_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un89_sum_cry_2 ;
    wire \b2v_inst11.mult1_un89_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un89_sum_cry_3 ;
    wire \b2v_inst11.mult1_un89_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un89_sum_cry_4 ;
    wire \b2v_inst11.mult1_un89_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un89_sum_cry_5 ;
    wire \b2v_inst11.mult1_un96_sum_axb_8 ;
    wire \b2v_inst11.mult1_un89_sum_cry_6 ;
    wire \b2v_inst11.mult1_un89_sum_cry_7 ;
    wire \b2v_inst11.mult1_un82_sum_i_0_8 ;
    wire bfn_4_3_0_;
    wire \b2v_inst11.mult1_un82_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_2 ;
    wire \b2v_inst11.mult1_un82_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_3 ;
    wire \b2v_inst11.mult1_un82_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_4 ;
    wire \b2v_inst11.mult1_un82_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_5 ;
    wire \b2v_inst11.mult1_un89_sum_axb_8 ;
    wire \b2v_inst11.mult1_un82_sum_cry_6 ;
    wire \b2v_inst11.mult1_un82_sum_cry_7 ;
    wire bfn_4_4_0_;
    wire \b2v_inst11.mult1_un75_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_2 ;
    wire \b2v_inst11.mult1_un75_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_3 ;
    wire \b2v_inst11.mult1_un75_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_4 ;
    wire \b2v_inst11.mult1_un75_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_5 ;
    wire \b2v_inst11.mult1_un82_sum_axb_8 ;
    wire \b2v_inst11.mult1_un75_sum_cry_6 ;
    wire \b2v_inst11.mult1_un75_sum_cry_7 ;
    wire \b2v_inst11.mult1_un75_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un75_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un40_sum_i_5_cascade_ ;
    wire \b2v_inst16.countZ0Z_10 ;
    wire \b2v_inst16.count_rst ;
    wire \b2v_inst16.count_4_10 ;
    wire bfn_4_6_0_;
    wire \b2v_inst11.mult1_un47_sum_cry_2 ;
    wire \b2v_inst11.mult1_un47_sum_cry_3 ;
    wire \b2v_inst11.mult1_un47_sum_cry_4 ;
    wire \b2v_inst11.mult1_un47_sum_cry_5 ;
    wire \b2v_inst200.count_enZ0 ;
    wire \b2v_inst11.un1_dutycycle_53_i_29 ;
    wire \b2v_inst11.mult1_un40_sum_i_l_ofx_4 ;
    wire \b2v_inst11.mult1_un47_sum_s_4_sf ;
    wire \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5 ;
    wire \b2v_inst11.count_clk_0_3 ;
    wire \b2v_inst11.count_clk_en ;
    wire \b2v_inst11.N_150_N ;
    wire \b2v_inst11.N_152_N_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_12_cascade_ ;
    wire \b2v_inst11.N_155_N_cascade_ ;
    wire \b2v_inst11.dutycycle_en_12 ;
    wire \b2v_inst11.dutycycle_en_12_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_15 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_12_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_10Z0Z_9_cascade_ ;
    wire \b2v_inst11.dutycycle_en_10 ;
    wire \b2v_inst11.dutycycleZ1Z_13 ;
    wire \b2v_inst11.dutycycleZ0Z_9_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_13_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_10_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIJU083Z0Z_8_cascade_ ;
    wire \b2v_inst11.N_108_f0_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIHTFQZ0Z_8 ;
    wire \b2v_inst11.dutycycle_RNI2NK31Z0Z_8_cascade_ ;
    wire \b2v_inst11.dutycycle_e_1_8 ;
    wire \b2v_inst11.dutycycleZ1Z_8 ;
    wire \b2v_inst11.N_108_f0 ;
    wire \b2v_inst11.dutycycle_e_1_8_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_1_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIJU083_0Z0Z_8 ;
    wire delayed_vccin_vccinaux_ok_RNIM6F44_0;
    wire \b2v_inst11.N_289_cascade_ ;
    wire \b2v_inst11.dutycycle_1_0_iv_i_0_2_cascade_ ;
    wire \b2v_inst11.N_302_cascade_ ;
    wire \b2v_inst11.N_301_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIGKEF3Z0Z_12 ;
    wire \b2v_inst11.dutycycleZ1Z_12 ;
    wire \b2v_inst11.dutycycle_RNIGKEF3Z0Z_12_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_10_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_56_a0_3_0_cascade_ ;
    wire \b2v_inst11.N_232_N ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_325_N_cascade_ ;
    wire \b2v_inst11.un1_func_state25_6_0_1_cascade_ ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_323_N ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_324_N ;
    wire \b2v_inst11.N_322 ;
    wire \b2v_inst11.count_offZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_offZ0Z_1 ;
    wire \b2v_inst11.count_off_RNIZ0Z_1 ;
    wire \b2v_inst11.count_off_RNIZ0Z_1_cascade_ ;
    wire \b2v_inst11.count_off_0_1 ;
    wire \b2v_inst11.count_offZ0Z_0 ;
    wire \b2v_inst11.count_off_0_0 ;
    wire \b2v_inst11.count_off_0_10 ;
    wire \b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2 ;
    wire \b2v_inst11.count_offZ0Z_10 ;
    wire \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5 ;
    wire \b2v_inst11.count_off_0_13 ;
    wire \b2v_inst11.count_off_enZ0 ;
    wire \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2 ;
    wire bfn_5_1_0_;
    wire \b2v_inst11.mult1_un110_sum_cry_2 ;
    wire \b2v_inst11.mult1_un110_sum_cry_3 ;
    wire \b2v_inst11.mult1_un110_sum_cry_4 ;
    wire \b2v_inst11.mult1_un110_sum_cry_5 ;
    wire \b2v_inst11.mult1_un110_sum_cry_6 ;
    wire \b2v_inst11.mult1_un110_sum_cry_7 ;
    wire \b2v_inst11.mult1_un89_sum_s_8 ;
    wire \b2v_inst11.mult1_un89_sum_i_0_8 ;
    wire bfn_5_2_0_;
    wire \b2v_inst11.mult1_un96_sum_i ;
    wire \b2v_inst11.mult1_un103_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_2 ;
    wire \b2v_inst11.mult1_un96_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_3 ;
    wire \b2v_inst11.mult1_un96_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_4 ;
    wire \b2v_inst11.mult1_un96_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_5 ;
    wire \b2v_inst11.mult1_un96_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un96_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un110_sum_axb_8 ;
    wire \b2v_inst11.mult1_un103_sum_cry_6 ;
    wire \b2v_inst11.mult1_un103_sum_axb_8 ;
    wire \b2v_inst11.mult1_un103_sum_cry_7 ;
    wire \b2v_inst11.mult1_un103_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un103_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un82_sum_i ;
    wire \b2v_inst11.mult1_un75_sum_i ;
    wire \b2v_inst11.mult1_un103_sum_i ;
    wire \b2v_inst11.mult1_un103_sum_s_8 ;
    wire bfn_5_4_0_;
    wire \b2v_inst11.mult1_un68_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_2_c ;
    wire \b2v_inst11.mult1_un68_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_3_c ;
    wire \b2v_inst11.mult1_un68_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_4_c ;
    wire \b2v_inst11.mult1_un68_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_5_c ;
    wire \b2v_inst11.mult1_un75_sum_axb_8 ;
    wire \b2v_inst11.mult1_un68_sum_cry_6_c ;
    wire \b2v_inst11.mult1_un68_sum_cry_7 ;
    wire \b2v_inst11.mult1_un68_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un68_sum_i_0_8 ;
    wire bfn_5_5_0_;
    wire \b2v_inst11.mult1_un61_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_2 ;
    wire \b2v_inst11.mult1_un61_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_3 ;
    wire \b2v_inst11.mult1_un61_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_4 ;
    wire \b2v_inst11.mult1_un61_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_5 ;
    wire \b2v_inst11.mult1_un68_sum_axb_8 ;
    wire \b2v_inst11.mult1_un61_sum_cry_6 ;
    wire \b2v_inst11.mult1_un61_sum_cry_7 ;
    wire bfn_5_6_0_;
    wire \b2v_inst11.mult1_un47_sum_i ;
    wire \b2v_inst11.mult1_un54_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un54_sum_cry_2 ;
    wire \b2v_inst11.mult1_un47_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un47_sum_l_fx_3 ;
    wire \b2v_inst11.mult1_un54_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un54_sum_cry_3 ;
    wire \b2v_inst11.mult1_un47_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un54_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un54_sum_cry_4 ;
    wire \b2v_inst11.mult1_un47_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un54_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un54_sum_cry_5 ;
    wire \b2v_inst11.mult1_un47_sum_l_fx_6 ;
    wire \b2v_inst11.mult1_un47_sum_s_6 ;
    wire \b2v_inst11.mult1_un61_sum_axb_8 ;
    wire \b2v_inst11.mult1_un54_sum_cry_6 ;
    wire \b2v_inst11.mult1_un40_sum_i_5 ;
    wire \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO ;
    wire \b2v_inst11.mult1_un54_sum_cry_7 ;
    wire \b2v_inst11.mult1_un54_sum_s_8 ;
    wire \b2v_inst11.mult1_un54_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un54_sum_i_8 ;
    wire \b2v_inst11.m15_e_2 ;
    wire bfn_5_7_0_;
    wire \b2v_inst11.un1_dutycycle_53_cry_0_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_1_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_2_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_3_cZ0 ;
    wire \b2v_inst11.mult1_un110_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_4_cZ0 ;
    wire \b2v_inst11.mult1_un103_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_5_cZ0 ;
    wire \b2v_inst11.mult1_un96_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_6_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_7_cZ0 ;
    wire bfn_5_8_0_;
    wire \b2v_inst11.mult1_un82_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_8_cZ0 ;
    wire \b2v_inst11.mult1_un75_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_9_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_10 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_11 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_13 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_12 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_13 ;
    wire \b2v_inst11.mult1_un47_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_13 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_14 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_15 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_14 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ;
    wire bfn_5_9_0_;
    wire \b2v_inst11.CO2 ;
    wire \b2v_inst11.CO2_THRU_CO ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_10 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_15 ;
    wire \b2v_inst11.un1_dutycycle_53_44_0_1_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_6Z0Z_9_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_11 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_15 ;
    wire \b2v_inst11.un1_m7_1_0_cascade_ ;
    wire \b2v_inst11.un1_i3_mux ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_11 ;
    wire \b2v_inst11.un1_dutycycle_53_44_0_2_tz ;
    wire \b2v_inst11.un1_dutycycle_53_39_0_0_1_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_39_0_0 ;
    wire \b2v_inst11.un1_dutycycle_53_39_1_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_41_0 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_13 ;
    wire \b2v_inst11.dutycycle_RNI_5Z0Z_9_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_10_1_0_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_7_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_12 ;
    wire \b2v_inst11.m18_i_1_0_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_11Z0Z_9 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_7 ;
    wire \b2v_inst11.dutycycle_RNI_5Z0Z_7 ;
    wire \b2v_inst11.dutycycle_RNI_5Z0Z_9 ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_7 ;
    wire \b2v_inst11.dutycycle_RNI_8Z0Z_9 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_7_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_11 ;
    wire \b2v_inst11.un1_dutycycle_53_13_1 ;
    wire \b2v_inst11.G_6_i_0_cascade_ ;
    wire \b2v_inst11.G_6_i_a4_1_1 ;
    wire \b2v_inst11.un1_dutycycle_53_7_1 ;
    wire \b2v_inst11.dutycycleZ0Z_11 ;
    wire \b2v_inst11.dutycycle_RNIGKEF3Z0Z_11 ;
    wire \b2v_inst11.dutycycleZ0Z_7_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_8_0 ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_11 ;
    wire \b2v_inst11.N_354 ;
    wire \b2v_inst11.N_354_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_11 ;
    wire \b2v_inst11.g2_1_1 ;
    wire \b2v_inst11.g3_0_1_cascade_ ;
    wire \b2v_inst11.N_14_0 ;
    wire \b2v_inst11.dutycycle_RNI_6Z0Z_5 ;
    wire \b2v_inst11.dutycycle_RNI_6Z0Z_5_cascade_ ;
    wire \b2v_inst11.count_clk_RNI_0Z0Z_1 ;
    wire \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_1_cascade_ ;
    wire \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_0_0 ;
    wire \b2v_inst11.N_122 ;
    wire \b2v_inst11.N_357 ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0 ;
    wire \b2v_inst11.un1_func_state25_6_0_a2_0 ;
    wire \b2v_inst11.N_327 ;
    wire \b2v_inst11.N_328 ;
    wire \b2v_inst11.func_state_1_m0_0_0_0_cascade_ ;
    wire bfn_6_1_0_;
    wire \b2v_inst11.mult1_un110_sum_i ;
    wire \b2v_inst11.mult1_un117_sum_cry_2 ;
    wire \b2v_inst11.mult1_un110_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un117_sum_cry_3 ;
    wire \b2v_inst11.mult1_un110_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un117_sum_cry_4 ;
    wire \b2v_inst11.mult1_un110_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un117_sum_cry_5 ;
    wire \b2v_inst11.mult1_un110_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un117_sum_cry_6 ;
    wire \b2v_inst11.mult1_un117_sum_axb_8 ;
    wire \b2v_inst11.mult1_un117_sum_cry_7 ;
    wire \b2v_inst11.mult1_un117_sum_s_8_cascade_ ;
    wire bfn_6_2_0_;
    wire \b2v_inst11.mult1_un124_sum_cry_2 ;
    wire \b2v_inst11.mult1_un117_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_3 ;
    wire \b2v_inst11.mult1_un117_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_4 ;
    wire \b2v_inst11.mult1_un117_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_5 ;
    wire \b2v_inst11.mult1_un117_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un117_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_6 ;
    wire \b2v_inst11.mult1_un124_sum_axb_8 ;
    wire \b2v_inst11.mult1_un124_sum_cry_7 ;
    wire \b2v_inst11.mult1_un110_sum_i_0_8 ;
    wire bfn_6_3_0_;
    wire \b2v_inst11.mult1_un124_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un131_sum_cry_2 ;
    wire \b2v_inst11.mult1_un131_sum_axb_4_l_fx ;
    wire \b2v_inst11.mult1_un124_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un131_sum_cry_3 ;
    wire \b2v_inst11.mult1_un124_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un131_sum_cry_4 ;
    wire \b2v_inst11.mult1_un124_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un131_sum_cry_5 ;
    wire \b2v_inst11.mult1_un131_sum_axb_7_l_fx ;
    wire \b2v_inst11.mult1_un124_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un131_sum_cry_6 ;
    wire \b2v_inst11.mult1_un131_sum_axb_8 ;
    wire \b2v_inst11.mult1_un131_sum_cry_7 ;
    wire \b2v_inst11.mult1_un131_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un68_sum ;
    wire \b2v_inst11.mult1_un68_sum_i ;
    wire \b2v_inst11.mult1_un117_sum_s_8 ;
    wire \b2v_inst11.mult1_un117_sum ;
    wire \b2v_inst11.mult1_un117_sum_i ;
    wire \b2v_inst11.mult1_un124_sum_s_8 ;
    wire \b2v_inst11.mult1_un124_sum ;
    wire \b2v_inst11.mult1_un124_sum_i ;
    wire \b2v_inst11.mult1_un89_sum ;
    wire \b2v_inst11.mult1_un89_sum_i ;
    wire \b2v_inst11.mult1_un61_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un110_sum_s_8 ;
    wire CONSTANT_ONE_NET;
    wire \b2v_inst11.mult1_un75_sum_s_8 ;
    wire \b2v_inst11.mult1_un61_sum_s_8 ;
    wire \b2v_inst11.mult1_un96_sum_s_8 ;
    wire \b2v_inst11.mult1_un54_sum ;
    wire \b2v_inst11.mult1_un54_sum_i ;
    wire \b2v_inst11.mult1_un61_sum ;
    wire \b2v_inst11.mult1_un61_sum_i ;
    wire \b2v_inst11.mult1_un68_sum_s_8 ;
    wire \b2v_inst16.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst16.curr_state_7_0_cascade_ ;
    wire \b2v_inst16.un13_clk_100khz_i ;
    wire \b2v_inst16.curr_state_0_1 ;
    wire \b2v_inst16.delayed_vddq_pwrgdZ0 ;
    wire b2v_inst16_un2_vpp_en_0_i;
    wire \b2v_inst16.curr_state_1_0 ;
    wire \b2v_inst16.curr_stateZ0Z_0 ;
    wire \b2v_inst16.curr_stateZ0Z_1 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_0 ;
    wire \b2v_inst200.count_RNIC03N_3Z0Z_0 ;
    wire V105A_EN_c;
    wire \b2v_inst11.dutycycle_RNIZ0Z_5 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_10 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_5 ;
    wire \b2v_inst11.dutycycleZ0Z_14 ;
    wire \b2v_inst11.dutycycle_en_11 ;
    wire \b2v_inst11.dutycycleZ0Z_13_cascade_ ;
    wire \b2v_inst11.un2_count_clk_17_0_a2_1_4 ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_4 ;
    wire \b2v_inst11.un1_dutycycle_53_50_a4_0_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_10 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_7 ;
    wire VCCST_OK_c;
    wire VDDQ_OK_c;
    wire VCCIO_EN_c;
    wire \b2v_inst11.dutycycle_RNIZ0Z_3 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_3_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_axb_7_1 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_9 ;
    wire \b2v_inst11.dutycycleZ0Z_8_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIAI7C4Z0Z_4_cascade_ ;
    wire \b2v_inst11.dutycycle_eena_2_0_1 ;
    wire \b2v_inst11.func_state_RNI3JFN6Z0Z_0_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI3JFN6Z0Z_4 ;
    wire \b2v_inst11.dutycycleZ1Z_4 ;
    wire \b2v_inst11.dutycycleZ1Z_9 ;
    wire \b2v_inst11.func_state_RNI3JFN6Z0Z_0 ;
    wire \b2v_inst11.dutycycle_RNI0KJ31Z0Z_7_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI74A23Z0Z_7_cascade_ ;
    wire \b2v_inst11.dutycycle_e_1_7 ;
    wire \b2v_inst11.dutycycle_RNI74A23Z0Z_7 ;
    wire \b2v_inst11.dutycycle_e_1_7_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI01TT1Z0Z_7 ;
    wire \b2v_inst11.dutycycle_RNI25OT3Z0Z_7_cascade_ ;
    wire \b2v_inst11.func_state_RNIGALV4Z0Z_0 ;
    wire \b2v_inst11.dutycycleZ1Z_7 ;
    wire \b2v_inst11.dutycycle_RNIGSFQZ0Z_7 ;
    wire bfn_6_13_0_;
    wire \b2v_inst11.un1_dutycycle_94_cry_0_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDUZ0Z8 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_1 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_2 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_3 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_4 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_5_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_6_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_7_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHPZ0Z49 ;
    wire bfn_6_14_0_;
    wire \b2v_inst11.dutycycleZ0Z_2 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_8_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_9_cZ0 ;
    wire \b2v_inst11.dutycycleZ0Z_7 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNPZ0Z5 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_10 ;
    wire \b2v_inst11.dutycycleZ0Z_10 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQZ0Z5 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_11 ;
    wire \b2v_inst11.dutycycleZ0Z_9 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_12 ;
    wire \b2v_inst11.dutycycleZ0Z_13 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_13 ;
    wire \b2v_inst11.dutycycleZ0Z_12 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_14 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5 ;
    wire \b2v_inst11.dutycycle_RNI_5Z0Z_5_cascade_ ;
    wire \b2v_inst11.N_156 ;
    wire \b2v_inst11.N_156_cascade_ ;
    wire \b2v_inst11.N_331 ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_307_N ;
    wire \b2v_inst11.dutycycle_RNI_5Z0Z_5 ;
    wire \b2v_inst11.N_4_cascade_ ;
    wire \b2v_inst11.func_state_RNI_0Z0Z_0_cascade_ ;
    wire \b2v_inst11.func_state_RNINJ641_0Z0Z_0 ;
    wire \b2v_inst11.func_state_RNINJ641_0Z0Z_0_cascade_ ;
    wire \b2v_inst11.count_off_RNIQCBN4Z0Z_9_cascade_ ;
    wire \b2v_inst11.N_333 ;
    wire \b2v_inst11.func_state_RNI_1Z0Z_1 ;
    wire \b2v_inst11.func_state_1_m2s2_i_1 ;
    wire \b2v_inst11.N_73 ;
    wire \b2v_inst11.func_state_1_m0_0 ;
    wire \b2v_inst11.N_73_cascade_ ;
    wire \b2v_inst11.count_off_RNIQCBN4Z0Z_9 ;
    wire \b2v_inst11.func_state_1_m0_1 ;
    wire bfn_7_2_0_;
    wire \b2v_inst11.mult1_un145_sum_cry_2 ;
    wire \b2v_inst11.mult1_un145_sum_cry_3 ;
    wire \b2v_inst11.mult1_un145_sum_cry_4 ;
    wire \b2v_inst11.mult1_un145_sum_cry_5 ;
    wire \b2v_inst11.mult1_un145_sum_cry_6 ;
    wire \b2v_inst11.mult1_un145_sum_cry_7 ;
    wire \b2v_inst11.mult1_un138_sum_i_0_8 ;
    wire bfn_7_3_0_;
    wire \b2v_inst11.mult1_un138_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_2 ;
    wire \b2v_inst11.mult1_un131_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_3 ;
    wire \b2v_inst11.mult1_un131_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_4 ;
    wire \b2v_inst11.mult1_un131_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_5 ;
    wire \b2v_inst11.mult1_un131_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un131_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un145_sum_axb_8 ;
    wire \b2v_inst11.mult1_un138_sum_cry_6 ;
    wire \b2v_inst11.mult1_un138_sum_axb_8 ;
    wire \b2v_inst11.mult1_un138_sum_cry_7 ;
    wire \b2v_inst11.mult1_un138_sum_s_8 ;
    wire \b2v_inst11.mult1_un138_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un82_sum_s_8 ;
    wire \b2v_inst11.mult1_un131_sum_s_8 ;
    wire \b2v_inst11.mult1_un138_sum ;
    wire \b2v_inst11.mult1_un138_sum_i ;
    wire \b2v_inst11.mult1_un131_sum ;
    wire \b2v_inst11.mult1_un131_sum_i ;
    wire \b2v_inst11.un1_count_cry_0_i ;
    wire bfn_7_5_0_;
    wire \b2v_inst11.un85_clk_100khz_1 ;
    wire \b2v_inst11.N_5647_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_0 ;
    wire \b2v_inst11.un85_clk_100khz_2 ;
    wire \b2v_inst11.N_5648_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_1 ;
    wire \b2v_inst11.un85_clk_100khz_3 ;
    wire \b2v_inst11.N_5649_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_2 ;
    wire \b2v_inst11.un85_clk_100khz_4 ;
    wire \b2v_inst11.N_5650_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_3 ;
    wire \b2v_inst11.un85_clk_100khz_5 ;
    wire \b2v_inst11.N_5651_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_4 ;
    wire \b2v_inst11.un85_clk_100khz_6 ;
    wire \b2v_inst11.N_5652_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_5 ;
    wire \b2v_inst11.un85_clk_100khz_7 ;
    wire \b2v_inst11.N_5653_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_6 ;
    wire \b2v_inst11.un85_clk_100khz_cry_7 ;
    wire \b2v_inst11.un85_clk_100khz_8 ;
    wire \b2v_inst11.N_5654_i ;
    wire bfn_7_6_0_;
    wire \b2v_inst11.un85_clk_100khz_9 ;
    wire \b2v_inst11.N_5655_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_8 ;
    wire \b2v_inst11.un85_clk_100khz_10 ;
    wire \b2v_inst11.N_5656_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_9 ;
    wire \b2v_inst11.un85_clk_100khz_11 ;
    wire \b2v_inst11.N_5657_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_10 ;
    wire \b2v_inst11.un85_clk_100khz_12 ;
    wire \b2v_inst11.N_5658_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_11 ;
    wire \b2v_inst11.un85_clk_100khz_13 ;
    wire \b2v_inst11.N_5659_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_12 ;
    wire \b2v_inst11.un85_clk_100khz_14 ;
    wire \b2v_inst11.N_5660_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_13 ;
    wire \b2v_inst11.mult1_un61_sum_i_8 ;
    wire \b2v_inst11.N_5661_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_14 ;
    wire \b2v_inst11.un85_clk_100khz_cry_15_cZ0 ;
    wire bfn_7_7_0_;
    wire \b2v_inst36.curr_state_RNI8TT2Z0Z_0 ;
    wire \b2v_inst11.pwm_out_en_cascade_ ;
    wire PWRBTN_LED_c;
    wire \b2v_inst11.pwm_out_1_sqmuxa_0 ;
    wire \b2v_inst11.curr_state_0_0 ;
    wire \b2v_inst11.curr_state_3_0 ;
    wire \b2v_inst11.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_0_sqmuxa_i_cascade_ ;
    wire \b2v_inst11.N_349 ;
    wire \b2v_inst11.un1_clk_100khz_32_and_i_o2_0_0_1 ;
    wire \b2v_inst11.dutycycle_RNIAI7C4Z0Z_10_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_5 ;
    wire \b2v_inst11.N_418 ;
    wire \b2v_inst11.func_state_RNIJU083Z0Z_0 ;
    wire \b2v_inst11.un1_clk_100khz_43_and_i_o2_0_0_1_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJTZ0Z69 ;
    wire \b2v_inst11.dutycycle_RNI4I3C2Z0Z_10 ;
    wire \b2v_inst11.dutycycle_RNI4I3C2Z0Z_10_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIAI7C4Z0Z_10 ;
    wire \b2v_inst11.dutycycleZ1Z_10 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_5 ;
    wire \b2v_inst11.d_i3_mux_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_5 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_3 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_3 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8 ;
    wire \b2v_inst11.dutycycle_e_1_3 ;
    wire \b2v_inst11.dutycycleZ1Z_3 ;
    wire \b2v_inst11.dutycycleZ0Z_6_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_1 ;
    wire \b2v_inst11.dutycycle_RNI_5Z0Z_3 ;
    wire \b2v_inst11.func_state_RNINJ641_0Z0Z_1_cascade_ ;
    wire \b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1_cascade_ ;
    wire \b2v_inst11.g0_2_3 ;
    wire \b2v_inst11.g0_2_2 ;
    wire \b2v_inst11.g0_1_1_0 ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3 ;
    wire \b2v_inst11.un1_clk_100khz_2_i_o3_out ;
    wire \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8 ;
    wire \b2v_inst11.dutycycle_1_0_1 ;
    wire \b2v_inst11.dutycycleZ1Z_1 ;
    wire \b2v_inst11.dutycycle_1_0_1_cascade_ ;
    wire \b2v_inst11.func_state_RNI_1Z0Z_0 ;
    wire \b2v_inst11.func_state_RNI_0Z0Z_1_cascade_ ;
    wire \b2v_inst11.un1_func_state25_4_i_a2_1_cascade_ ;
    wire \b2v_inst11.N_321 ;
    wire \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ;
    wire \b2v_inst11.dutycycle_1_0_0_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIZ0 ;
    wire \b2v_inst11.g1 ;
    wire \b2v_inst11.dutycycle_0_6 ;
    wire \b2v_inst11.g1_cascade_ ;
    wire \b2v_inst11.g1_0 ;
    wire \b2v_inst11.dutycycle_eena ;
    wire \b2v_inst11.dutycycle_1_0_0 ;
    wire \b2v_inst11.dutycycle_eena_cascade_ ;
    wire \b2v_inst11.dutycycleZ1Z_0 ;
    wire \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_sx ;
    wire \b2v_inst11.func_state_RNI_0Z0Z_1 ;
    wire \b2v_inst11.func_state_1_m0_0_0_1 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_0 ;
    wire \b2v_inst11.N_360 ;
    wire \b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_0_cascade_ ;
    wire \b2v_inst11.func_stateZ0Z_0 ;
    wire \b2v_inst11.func_stateZ0Z_0_cascade_ ;
    wire \b2v_inst11.N_3013_i_cascade_ ;
    wire \b2v_inst11.N_330 ;
    wire \b2v_inst11.func_state_RNI_0Z0Z_0 ;
    wire \b2v_inst11.g1_1 ;
    wire \b2v_inst11.func_state_RNI673P9Z0Z_0 ;
    wire \b2v_inst11.func_stateZ1Z_0 ;
    wire \b2v_inst11.count_off_RNIZ0Z_9 ;
    wire \b2v_inst11.N_335_cascade_ ;
    wire \b2v_inst11.count_off_RNIQ1RAS1Z0Z_9 ;
    wire \b2v_inst11.func_state_1_ss0_i_0_o2_0 ;
    wire \b2v_inst36.count_rst_11_cascade_ ;
    wire \b2v_inst36.countZ0Z_7_cascade_ ;
    wire \b2v_inst36.count_1_7 ;
    wire \b2v_inst36.count_rst_9_cascade_ ;
    wire \b2v_inst36.countZ0Z_5_cascade_ ;
    wire \b2v_inst36.count_1_5 ;
    wire \b2v_inst36.count_rst_7 ;
    wire \b2v_inst36.count_rst_6_cascade_ ;
    wire \b2v_inst36.countZ0Z_8_cascade_ ;
    wire \b2v_inst36.count_1_8 ;
    wire \b2v_inst36.count_rst_4_cascade_ ;
    wire \b2v_inst36.countZ0Z_10_cascade_ ;
    wire \b2v_inst36.count_1_10 ;
    wire bfn_8_3_0_;
    wire \b2v_inst11.mult1_un145_sum_i ;
    wire \b2v_inst11.mult1_un152_sum_cry_2 ;
    wire \b2v_inst11.mult1_un145_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_3 ;
    wire \b2v_inst11.mult1_un145_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_4 ;
    wire \b2v_inst11.mult1_un145_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_5 ;
    wire \b2v_inst11.mult1_un145_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un152_sum_cry_6 ;
    wire \b2v_inst11.mult1_un152_sum_axb_8 ;
    wire \b2v_inst11.mult1_un152_sum_cry_7 ;
    wire \b2v_inst11.mult1_un145_sum_s_8 ;
    wire \b2v_inst11.mult1_un145_sum_i_0_8 ;
    wire bfn_8_4_0_;
    wire \b2v_inst11.mult1_un159_sum_cry_1 ;
    wire \b2v_inst11.mult1_un152_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_2 ;
    wire \b2v_inst11.mult1_un152_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_3 ;
    wire \b2v_inst11.mult1_un152_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_4 ;
    wire \b2v_inst11.mult1_un152_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_5 ;
    wire \b2v_inst11.mult1_un159_sum_axb_7 ;
    wire \b2v_inst11.mult1_un159_sum_cry_6 ;
    wire \b2v_inst11.mult1_un152_sum_s_8 ;
    wire \b2v_inst11.mult1_un152_sum_i_0_8 ;
    wire \b2v_inst11.count_0_14 ;
    wire \b2v_inst11.count_0_6 ;
    wire \b2v_inst11.count_0_15 ;
    wire \b2v_inst11.count_0_7 ;
    wire bfn_8_6_0_;
    wire \b2v_inst11.un1_count_cry_1 ;
    wire \b2v_inst11.un1_count_cry_2 ;
    wire \b2v_inst11.un1_count_cry_3 ;
    wire \b2v_inst11.un1_count_cry_4 ;
    wire \b2v_inst11.un1_count_cry_5_c_RNIMQUDZ0 ;
    wire \b2v_inst11.un1_count_cry_5 ;
    wire \b2v_inst11.un1_count_cry_6_c_RNINSVDZ0 ;
    wire \b2v_inst11.un1_count_cry_6 ;
    wire \b2v_inst11.un1_count_cry_7 ;
    wire \b2v_inst11.un1_count_cry_8 ;
    wire bfn_8_7_0_;
    wire \b2v_inst11.un1_count_cry_9 ;
    wire \b2v_inst11.un1_count_cry_10 ;
    wire \b2v_inst11.un1_count_cry_11 ;
    wire \b2v_inst11.un1_count_cry_12 ;
    wire \b2v_inst11.un1_count_cry_13_c_RNI5AUZ0Z6 ;
    wire \b2v_inst11.un1_count_cry_13 ;
    wire \b2v_inst11.un1_count_cry_14 ;
    wire \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6 ;
    wire \b2v_inst11.un1_count_cry_9_c_RNIQ23EZ0 ;
    wire \b2v_inst11.count_0_10 ;
    wire \b2v_inst11.un1_count_cry_10_c_RNI24RZ0Z6 ;
    wire \b2v_inst11.count_0_11 ;
    wire \b2v_inst11.un1_count_cry_1_c_RNIIIQDZ0 ;
    wire \b2v_inst11.count_0_2 ;
    wire \b2v_inst11.un1_count_cry_11_c_RNI36SZ0Z6 ;
    wire \b2v_inst11.count_0_12 ;
    wire G_2727_cascade_;
    wire \b2v_inst5.curr_state_2_1 ;
    wire N_229_cascade_;
    wire \b2v_inst5.curr_stateZ0Z_1 ;
    wire \b2v_inst5.curr_stateZ0Z_1_cascade_ ;
    wire curr_state_RNI5VS71_0_1_cascade_;
    wire \b2v_inst11.mult1_un145_sum ;
    wire RSMRSTn_RNI8DFE_cascade_;
    wire \b2v_inst11.g0_1_1 ;
    wire \b2v_inst11.N_182 ;
    wire \b2v_inst11.func_state_RNIT4D71_0Z0Z_1 ;
    wire \b2v_inst11.dutycycle_0_5 ;
    wire \b2v_inst11.g1_4_0 ;
    wire \b2v_inst11.func_state_RNIT4D71_0Z0Z_1_cascade_ ;
    wire dutycycle_RNIIOE3D_0_5_cascade_;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_5_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_53_axb_3_1_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_2 ;
    wire \b2v_inst11.un1_i3_mux_1 ;
    wire \b2v_inst11.g0_6_2 ;
    wire \b2v_inst11.m15_e_3 ;
    wire \b2v_inst11.un1_dutycycle_inv_4_0 ;
    wire \b2v_inst11.g0_9_1 ;
    wire \b2v_inst11.g1_0_1_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_164_0 ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_5 ;
    wire \b2v_inst11.mult1_un152_sum_i ;
    wire \b2v_inst11.N_3013_i ;
    wire \b2v_inst11.N_221_iZ0 ;
    wire \b2v_inst11.func_state_cascade_ ;
    wire \b2v_inst11.N_303_cascade_ ;
    wire \b2v_inst11.dutycycle_eena_1 ;
    wire \b2v_inst11.N_70 ;
    wire \b2v_inst11.dutycycle_eena_1_cascade_ ;
    wire \b2v_inst11.dutycycleZ1Z_2 ;
    wire \b2v_inst11.dutycycle_eena_0 ;
    wire \b2v_inst11.N_169 ;
    wire \b2v_inst11.N_375 ;
    wire \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_sxZ0_cascade_ ;
    wire SYNTHESIZED_WIRE_47keep_fast;
    wire \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_1 ;
    wire \b2v_inst11.un1_clk_100khz_26_and_i_o2_1 ;
    wire \b2v_inst11.dutycycle_RNINJ641_0Z0Z_5 ;
    wire \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_cascade_ ;
    wire \b2v_inst11.N_183 ;
    wire \b2v_inst11.func_state_RNI_3Z0Z_1 ;
    wire \b2v_inst11.N_183_cascade_ ;
    wire \b2v_inst11.N_114_f0_1 ;
    wire \b2v_inst11.dutycycleZ0Z_6 ;
    wire \b2v_inst11.N_379 ;
    wire \b2v_inst6.curr_state_RNI8OKQ2Z0Z_0_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_52_and_i_a2Z0Z_1 ;
    wire \b2v_inst11.func_state_RNIDINH9Z0Z_0 ;
    wire \b2v_inst11.func_stateZ0Z_1 ;
    wire \b2v_inst6.curr_state_RNI8OKQ2Z0Z_0 ;
    wire \b2v_inst6.delayed_vccin_vccinaux_ok_0 ;
    wire SYNTHESIZED_WIRE_49_i_0_o3_0;
    wire VPP_OK_c;
    wire VDDQ_EN_c;
    wire VCCIO_OK_c;
    wire V5S_OK_c;
    wire \b2v_inst31.un8_outputZ0Z_0 ;
    wire V33S_OK_c;
    wire VCCIN_EN_c;
    wire bfn_9_1_0_;
    wire \b2v_inst36.un2_count_1_cry_1 ;
    wire \b2v_inst36.un2_count_1_cry_2 ;
    wire \b2v_inst36.un2_count_1_cry_3 ;
    wire \b2v_inst36.countZ0Z_5 ;
    wire \b2v_inst36.un2_count_1_cry_4_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_4 ;
    wire \b2v_inst36.un2_count_1_cry_5 ;
    wire \b2v_inst36.countZ0Z_7 ;
    wire \b2v_inst36.un2_count_1_cry_6_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_6 ;
    wire \b2v_inst36.un2_count_1_cry_7_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_7 ;
    wire \b2v_inst36.un2_count_1_cry_8 ;
    wire bfn_9_2_0_;
    wire \b2v_inst36.un2_count_1_cry_9_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_9 ;
    wire \b2v_inst36.un2_count_1_cry_10 ;
    wire \b2v_inst36.un2_count_1_cry_11 ;
    wire \b2v_inst36.un2_count_1_cry_12 ;
    wire \b2v_inst36.un2_count_1_cry_13 ;
    wire \b2v_inst36.un2_count_1_cry_14 ;
    wire \b2v_inst36.count_1_12 ;
    wire \b2v_inst36.count_en_cascade_ ;
    wire \b2v_inst36.count_rst_2 ;
    wire \b2v_inst36.count_rst_0 ;
    wire \b2v_inst36.count_1_14 ;
    wire \b2v_inst36.count_rst ;
    wire \b2v_inst36.count_1_15 ;
    wire \b2v_inst11.dutycycleZ0Z_0 ;
    wire bfn_9_4_0_;
    wire \b2v_inst11.mult1_un166_sum_cry_0 ;
    wire \b2v_inst11.mult1_un159_sum_cry_2_s ;
    wire \b2v_inst11.mult1_un166_sum_cry_1 ;
    wire \b2v_inst11.mult1_un159_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un166_sum_cry_2 ;
    wire \b2v_inst11.mult1_un159_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un159_sum_s_7 ;
    wire \b2v_inst11.mult1_un166_sum_cry_3 ;
    wire G_2890;
    wire \b2v_inst11.mult1_un159_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un166_sum_cry_4 ;
    wire \b2v_inst11.mult1_un166_sum_axb_6 ;
    wire \b2v_inst11.mult1_un166_sum_cry_5 ;
    wire \b2v_inst11.un85_clk_100khz_0 ;
    wire \b2v_inst11.dutycycle ;
    wire \b2v_inst11.mult1_un159_sum_i ;
    wire \b2v_inst11.countZ0Z_2 ;
    wire \b2v_inst11.countZ0Z_7 ;
    wire \b2v_inst11.countZ0Z_15 ;
    wire \b2v_inst11.countZ0Z_11 ;
    wire \b2v_inst11.countZ0Z_10 ;
    wire \b2v_inst11.countZ0Z_12 ;
    wire \b2v_inst11.un79_clk_100khzlt6 ;
    wire \b2v_inst11.countZ0Z_6 ;
    wire \b2v_inst11.un79_clk_100khzlto15_5_cascade_ ;
    wire \b2v_inst11.countZ0Z_14 ;
    wire \b2v_inst11.un79_clk_100khzlto15_7_cascade_ ;
    wire \b2v_inst11.un79_clk_100khzlto15_4 ;
    wire \b2v_inst11.count_RNIZ0Z_13 ;
    wire \b2v_inst11.curr_stateZ0Z_0 ;
    wire \b2v_inst11.count_RNIZ0Z_13_cascade_ ;
    wire \b2v_inst11.countZ0Z_3 ;
    wire \b2v_inst11.un1_count_cry_2_c_RNIJKRDZ0 ;
    wire \b2v_inst11.count_0_3 ;
    wire \b2v_inst11.countZ0Z_13 ;
    wire \b2v_inst11.un1_count_cry_12_c_RNI48TZ0Z6 ;
    wire \b2v_inst11.count_0_13 ;
    wire \b2v_inst11.countZ0Z_4 ;
    wire \b2v_inst11.un1_count_cry_3_c_RNIKMSDZ0 ;
    wire \b2v_inst11.count_0_4 ;
    wire \b2v_inst11.countZ0Z_5 ;
    wire \b2v_inst11.un1_count_cry_4_c_RNILOTDZ0 ;
    wire \b2v_inst11.count_0_5 ;
    wire \b2v_inst11.count_0_0 ;
    wire \b2v_inst11.count_RNI_2_0 ;
    wire \b2v_inst11.countZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_RNIZ0Z_1_cascade_ ;
    wire \b2v_inst11.countZ0Z_1 ;
    wire \b2v_inst11.countZ0Z_0 ;
    wire \b2v_inst11.countZ0Z_1_cascade_ ;
    wire \b2v_inst11.count_0_sqmuxa_i ;
    wire \b2v_inst11.count_0_1 ;
    wire \b2v_inst11.countZ0Z_8 ;
    wire \b2v_inst11.un1_count_cry_7_c_RNIOU0EZ0 ;
    wire \b2v_inst11.count_0_8 ;
    wire \b2v_inst11.countZ0Z_9 ;
    wire \b2v_inst11.un1_count_cry_8_c_RNIP02EZ0 ;
    wire \b2v_inst11.count_0_9 ;
    wire \b2v_inst5.curr_state_3_0 ;
    wire \b2v_inst5.curr_stateZ0Z_0 ;
    wire G_2727;
    wire \b2v_inst5.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst5.m4_0 ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1 ;
    wire \b2v_inst11.dutycycleZ0Z_4 ;
    wire \b2v_inst11.dutycycle_RNITBKN1Z0Z_7 ;
    wire N_229;
    wire \b2v_inst5.count_enZ0_cascade_ ;
    wire \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO ;
    wire \b2v_inst11.g0_2_1 ;
    wire \b2v_inst11.pwm_outZ0 ;
    wire \b2v_inst11.pwm_out_1_sqmuxa ;
    wire \b2v_inst20.un4_counter_0_and ;
    wire bfn_9_9_0_;
    wire \b2v_inst20.un4_counter_0 ;
    wire \b2v_inst20.un4_counter_1 ;
    wire \b2v_inst20.un4_counter_2 ;
    wire \b2v_inst20.un4_counter_3 ;
    wire \b2v_inst20.un4_counter_4 ;
    wire \b2v_inst20.un4_counter_5 ;
    wire \b2v_inst20.un4_counter_6 ;
    wire b2v_inst20_un4_counter_7;
    wire bfn_9_10_0_;
    wire \b2v_inst20.un4_counter_1_and ;
    wire curr_state_RNI5VS71_0_1;
    wire RSMRSTn_0;
    wire \b2v_inst11.N_234_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_52_and_i_0_0_cascade_ ;
    wire SYNTHESIZED_WIRE_47keep_rep1;
    wire b2v_inst20_un4_counter_7_THRU_CO;
    wire dutycycle_RNIIOE3D_0_5;
    wire b2v_inst11_count_off_1_sqmuxa_0_0_0;
    wire G_26_0_a5_1_0;
    wire G_26_0_a5_2_1_cascade_;
    wire G_26_0_0;
    wire \b2v_inst11.g2_0_1 ;
    wire \b2v_inst11.un1_dutycycle_172_m4 ;
    wire b2v_inst11_un1_dutycycle_172_m3_0_0_0_cascade_;
    wire \b2v_inst11.g2_1 ;
    wire \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z2 ;
    wire \b2v_inst11.g4_cascade_ ;
    wire b2v_inst16_delayed_vddq_pwrgd_en;
    wire \b2v_inst11.N_5 ;
    wire \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_xZ0 ;
    wire \b2v_inst11.dutycycleZ0Z_3 ;
    wire \b2v_inst11.N_12 ;
    wire \b2v_inst11.func_state_RNINJ641_0Z0Z_1 ;
    wire N_4;
    wire G_26_0_a5_2;
    wire \b2v_inst11.N_158 ;
    wire \b2v_inst11.N_3046_i ;
    wire \b2v_inst11.g3_0 ;
    wire \b2v_inst11.g2_0_cascade_ ;
    wire RSMRSTn_RNI8DFE;
    wire \b2v_inst11.N_228_N_0 ;
    wire \b2v_inst6.delayed_vccin_vccinaux_okZ0 ;
    wire \b2v_inst11.g1_4_2_0 ;
    wire \b2v_inst11.dutycycleZ0Z_8 ;
    wire N_19_i;
    wire \b2v_inst11.g0_8_0_0 ;
    wire SLP_S4n_c;
    wire GPIO_FPGA_PCH_5_c;
    wire \b2v_inst11.func_state ;
    wire SLP_S3n_c;
    wire \b2v_inst11.count_clk_RNIZ0Z_3 ;
    wire \b2v_inst11.g1_2_1_cascade_ ;
    wire \b2v_inst11.dutycycleZ1Z_6 ;
    wire \b2v_inst11.g1_2 ;
    wire \b2v_inst6.countZ0Z_11_cascade_ ;
    wire \b2v_inst6.count_3_11 ;
    wire \b2v_inst6.curr_state_RNIDMSJ1Z0Z_1 ;
    wire \b2v_inst6.count_rst_10 ;
    wire \b2v_inst6.count_rst_3_cascade_ ;
    wire \b2v_inst6.countZ0Z_4_cascade_ ;
    wire \b2v_inst6.count_3_4 ;
    wire G_2746_cascade_;
    wire \b2v_inst6.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst6.curr_state_2_0 ;
    wire VR_READY_VCCIN_c;
    wire VR_READY_VCCINAUX_c;
    wire SYNTHESIZED_WIRE_48_i_0_o3_2;
    wire \b2v_inst6.N_413_cascade_ ;
    wire \b2v_inst6.curr_state_7_1_cascade_ ;
    wire \b2v_inst6.curr_stateZ0Z_1 ;
    wire \b2v_inst6.curr_stateZ0Z_0 ;
    wire \b2v_inst6.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst6.N_413 ;
    wire \b2v_inst6.curr_state_1_1 ;
    wire \b2v_inst36.countZ0Z_1_cascade_ ;
    wire \b2v_inst36.count_rst_13 ;
    wire \b2v_inst36.countZ0Z_14 ;
    wire \b2v_inst36.countZ0Z_15 ;
    wire \b2v_inst36.count_1_1 ;
    wire \b2v_inst36.count_rst_12_cascade_ ;
    wire \b2v_inst36.countZ0Z_2 ;
    wire \b2v_inst36.countZ0Z_2_cascade_ ;
    wire \b2v_inst36.un2_count_1_cry_1_THRU_CO ;
    wire \b2v_inst36.count_1_2 ;
    wire \b2v_inst36.countZ0Z_3 ;
    wire \b2v_inst36.un2_count_1_cry_2_THRU_CO ;
    wire \b2v_inst36.count_1_3 ;
    wire \b2v_inst36.countZ0Z_8 ;
    wire \b2v_inst36.countZ0Z_10 ;
    wire \b2v_inst36.countZ0Z_1 ;
    wire \b2v_inst36.un12_clk_100khz_11 ;
    wire \b2v_inst36.un12_clk_100khz_10_cascade_ ;
    wire \b2v_inst36.un12_clk_100khz_8 ;
    wire \b2v_inst36.un2_count_1_axb_6 ;
    wire \b2v_inst36.count_rst_3 ;
    wire \b2v_inst36.countZ0Z_11 ;
    wire \b2v_inst36.un2_count_1_cry_10_THRU_CO ;
    wire \b2v_inst36.countZ0Z_11_cascade_ ;
    wire \b2v_inst36.count_1_11 ;
    wire \b2v_inst36.count_rst_8 ;
    wire \b2v_inst36.count_1_6 ;
    wire \b2v_inst36.countZ0Z_12 ;
    wire \b2v_inst36.countZ0Z_6_cascade_ ;
    wire \b2v_inst36.un12_clk_100khz_9 ;
    wire \b2v_inst36.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst36.curr_state_7_0_cascade_ ;
    wire \b2v_inst36.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst36.DSW_PWROK_0 ;
    wire \b2v_inst36.curr_state_3_1 ;
    wire \b2v_inst36.curr_state_7_1 ;
    wire \b2v_inst36.curr_stateZ0Z_0 ;
    wire \b2v_inst36.curr_state_4_0 ;
    wire \b2v_inst36.curr_stateZ0Z_1 ;
    wire V33DSW_OK_c;
    wire \b2v_inst36.N_2925_i ;
    wire \b2v_inst5.count_0_14 ;
    wire \b2v_inst5.count_0_7 ;
    wire \b2v_inst16.countZ0Z_8 ;
    wire \b2v_inst16.count_rst_13 ;
    wire \b2v_inst16.count_4_8 ;
    wire \b2v_inst16.countZ0Z_9 ;
    wire \b2v_inst16.count_rst_14 ;
    wire \b2v_inst16.count_4_9 ;
    wire \b2v_inst16.count_en ;
    wire \b2v_inst36.count_1_4 ;
    wire \b2v_inst36.count_rst_10 ;
    wire \b2v_inst36.countZ0Z_4 ;
    wire \b2v_inst5.N_2906_i_cascade_ ;
    wire \b2v_inst5.count_1_i_a2_1_0_cascade_ ;
    wire \b2v_inst5.count_0_12 ;
    wire \b2v_inst5.count_1_i_a2_0_0 ;
    wire \b2v_inst5.count_0_5 ;
    wire \b2v_inst5.count_0_6 ;
    wire \b2v_inst5.count_1_i_a2_2_0 ;
    wire bfn_11_7_0_;
    wire \b2v_inst5.un2_count_1_cry_1 ;
    wire \b2v_inst5.un2_count_1_cry_2 ;
    wire \b2v_inst5.un2_count_1_cry_3 ;
    wire \b2v_inst5.un2_count_1_axb_5 ;
    wire \b2v_inst5.count_rst_9 ;
    wire \b2v_inst5.un2_count_1_cry_4 ;
    wire \b2v_inst5.un2_count_1_axb_6 ;
    wire \b2v_inst5.count_rst_8 ;
    wire \b2v_inst5.un2_count_1_cry_5 ;
    wire \b2v_inst5.countZ0Z_7 ;
    wire \b2v_inst5.count_rst_7 ;
    wire \b2v_inst5.un2_count_1_cry_6 ;
    wire \b2v_inst5.un2_count_1_cry_7 ;
    wire \b2v_inst5.un2_count_1_cry_8 ;
    wire bfn_11_8_0_;
    wire \b2v_inst5.un2_count_1_cry_9 ;
    wire \b2v_inst5.un2_count_1_cry_10 ;
    wire \b2v_inst5.un2_count_1_axb_12 ;
    wire \b2v_inst5.count_rst_2 ;
    wire \b2v_inst5.un2_count_1_cry_11 ;
    wire \b2v_inst5.un2_count_1_cry_12 ;
    wire \b2v_inst5.countZ0Z_14 ;
    wire \b2v_inst5.count_rst_0 ;
    wire \b2v_inst5.un2_count_1_cry_13 ;
    wire \b2v_inst5.countZ0Z_15 ;
    wire \b2v_inst5.un2_count_1_cry_14 ;
    wire \b2v_inst5.count_rst ;
    wire \b2v_inst5.count_0_15 ;
    wire \b2v_inst20.counterZ0Z_1 ;
    wire \b2v_inst20.counterZ0Z_0 ;
    wire bfn_11_9_0_;
    wire \b2v_inst20.counterZ0Z_2 ;
    wire \b2v_inst20.counter_1_cry_1_THRU_CO ;
    wire \b2v_inst20.counter_1_cry_1 ;
    wire \b2v_inst20.counterZ0Z_3 ;
    wire \b2v_inst20.counter_1_cry_2_THRU_CO ;
    wire \b2v_inst20.counter_1_cry_2 ;
    wire \b2v_inst20.counterZ0Z_4 ;
    wire \b2v_inst20.counter_1_cry_3_THRU_CO ;
    wire \b2v_inst20.counter_1_cry_3 ;
    wire \b2v_inst20.counterZ0Z_5 ;
    wire \b2v_inst20.counter_1_cry_4_THRU_CO ;
    wire \b2v_inst20.counter_1_cry_4 ;
    wire \b2v_inst20.counterZ0Z_6 ;
    wire \b2v_inst20.counter_1_cry_5_THRU_CO ;
    wire \b2v_inst20.counter_1_cry_5 ;
    wire \b2v_inst20.counterZ0Z_7 ;
    wire \b2v_inst20.counter_1_cry_6 ;
    wire \b2v_inst20.counter_1_cry_7 ;
    wire \b2v_inst20.counter_1_cry_8 ;
    wire bfn_11_10_0_;
    wire \b2v_inst20.counter_1_cry_9 ;
    wire \b2v_inst20.counter_1_cry_10 ;
    wire \b2v_inst20.counter_1_cry_11 ;
    wire \b2v_inst20.counter_1_cry_12 ;
    wire \b2v_inst20.counter_1_cry_13 ;
    wire \b2v_inst20.counter_1_cry_14 ;
    wire \b2v_inst20.counter_1_cry_15 ;
    wire \b2v_inst20.counter_1_cry_16 ;
    wire bfn_11_11_0_;
    wire \b2v_inst20.counter_1_cry_17 ;
    wire \b2v_inst20.counter_1_cry_18 ;
    wire \b2v_inst20.counter_1_cry_19 ;
    wire \b2v_inst20.counter_1_cry_20 ;
    wire \b2v_inst20.counter_1_cry_21 ;
    wire \b2v_inst20.counter_1_cry_22 ;
    wire \b2v_inst20.counter_1_cry_23 ;
    wire \b2v_inst20.counter_1_cry_24 ;
    wire bfn_11_12_0_;
    wire \b2v_inst20.counter_1_cry_25 ;
    wire \b2v_inst20.counter_1_cry_26 ;
    wire \b2v_inst20.counter_1_cry_27 ;
    wire \b2v_inst20.counter_1_cry_28 ;
    wire \b2v_inst20.counter_1_cry_29 ;
    wire \b2v_inst20.counter_1_cry_30 ;
    wire bfn_11_13_0_;
    wire \b2v_inst6.un2_count_1_cry_1 ;
    wire \b2v_inst6.un2_count_1_cry_2 ;
    wire \b2v_inst6.un2_count_1_cry_3_THRU_CO ;
    wire \b2v_inst6.un2_count_1_cry_3 ;
    wire \b2v_inst6.un2_count_1_cry_4 ;
    wire \b2v_inst6.un2_count_1_cry_5 ;
    wire \b2v_inst6.un2_count_1_cry_6 ;
    wire \b2v_inst6.un2_count_1_cry_7 ;
    wire \b2v_inst6.un2_count_1_cry_8 ;
    wire bfn_11_14_0_;
    wire \b2v_inst6.un2_count_1_cry_9 ;
    wire \b2v_inst6.un2_count_1_cry_10_THRU_CO ;
    wire \b2v_inst6.un2_count_1_cry_10 ;
    wire \b2v_inst6.un2_count_1_cry_11 ;
    wire \b2v_inst6.un2_count_1_cry_12 ;
    wire \b2v_inst6.un2_count_1_cry_13 ;
    wire \b2v_inst6.un2_count_1_cry_14 ;
    wire \b2v_inst6.un2_count_1_cry_4_THRU_CO ;
    wire \b2v_inst6.count_rst_4_cascade_ ;
    wire \b2v_inst6.count_3_5 ;
    wire \b2v_inst6.count_rst_2_cascade_ ;
    wire \b2v_inst6.count_rst_8_cascade_ ;
    wire \b2v_inst6.count_rst_9 ;
    wire \b2v_inst6.count_3_10 ;
    wire \b2v_inst6.countZ0Z_11 ;
    wire \b2v_inst6.count_rst_6_cascade_ ;
    wire \b2v_inst6.countZ0Z_7 ;
    wire \b2v_inst6.un2_count_1_cry_6_THRU_CO ;
    wire \b2v_inst6.countZ0Z_7_cascade_ ;
    wire \b2v_inst6.count_3_7 ;
    wire \b2v_inst6.count_rst_7_cascade_ ;
    wire \b2v_inst6.countZ0Z_8 ;
    wire \b2v_inst6.countZ0Z_8_cascade_ ;
    wire \b2v_inst6.un2_count_1_cry_7_THRU_CO ;
    wire \b2v_inst6.count_3_8 ;
    wire \b2v_inst6.countZ0Z_9 ;
    wire \b2v_inst6.un2_count_1_cry_8_THRU_CO ;
    wire \b2v_inst6.count_3_9 ;
    wire \b2v_inst36.N_2928_i_cascade_ ;
    wire \b2v_inst36.count_1_13 ;
    wire \b2v_inst36.un2_count_1_cry_12_c_RNIS7LZ0Z1 ;
    wire \b2v_inst36.countZ0Z_13 ;
    wire \b2v_inst36.countZ0Z_9 ;
    wire \b2v_inst36.un2_count_1_cry_8_c_RNIH8IZ0Z8 ;
    wire \b2v_inst36.count_1_9 ;
    wire \b2v_inst36.count_rst_14 ;
    wire \b2v_inst36.countZ0Z_0 ;
    wire \b2v_inst36.N_2928_i ;
    wire \b2v_inst36.countZ0Z_0_cascade_ ;
    wire \b2v_inst36.N_1_i ;
    wire \b2v_inst36.count_1_0 ;
    wire \b2v_inst36.count_en ;
    wire \b2v_inst36.count_0_sqmuxa ;
    wire \b2v_inst5.count_rst_5 ;
    wire \b2v_inst5.count_rst_5_cascade_ ;
    wire \b2v_inst5.un2_count_1_axb_9 ;
    wire \b2v_inst5.un2_count_1_cry_8_THRU_CO ;
    wire \b2v_inst5.un2_count_1_axb_9_cascade_ ;
    wire \b2v_inst5.count_0_9 ;
    wire \b2v_inst5.count_rst_4_cascade_ ;
    wire \b2v_inst5.countZ0Z_10 ;
    wire \b2v_inst5.countZ0Z_10_cascade_ ;
    wire \b2v_inst5.un2_count_1_cry_9_THRU_CO ;
    wire \b2v_inst5.count_0_10 ;
    wire \b2v_inst5.count_RNIRHC7IZ0Z_2_cascade_ ;
    wire \b2v_inst5.countZ0Z_0 ;
    wire \b2v_inst5.countZ0Z_0_cascade_ ;
    wire \b2v_inst5.count_RNIZ0Z_0_cascade_ ;
    wire \b2v_inst5.count_RNIZ0Z_0 ;
    wire \b2v_inst5.count_0_1 ;
    wire \b2v_inst5.count_1_i_a2_11_0 ;
    wire \b2v_inst5.N_2906_i ;
    wire \b2v_inst5.count_0_0 ;
    wire \b2v_inst5.count_0_3 ;
    wire \b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9 ;
    wire \b2v_inst5.countZ0Z_3 ;
    wire \b2v_inst5.count_1_i_a2_6_0 ;
    wire \b2v_inst5.count_1_i_a2_4_0_cascade_ ;
    wire \b2v_inst5.count_1_i_a2_12_0 ;
    wire \b2v_inst5.count_0_2 ;
    wire \b2v_inst5.count_rst_12 ;
    wire \b2v_inst5.un2_count_1_axb_2 ;
    wire \b2v_inst5.countZ0Z_1 ;
    wire \b2v_inst5.count_1_i_a2_3_0 ;
    wire \b2v_inst5.count_0_11 ;
    wire \b2v_inst5.count_rst_3 ;
    wire \b2v_inst5.un2_count_1_axb_11 ;
    wire \b2v_inst5.count_1_i_a2_5_0 ;
    wire \b2v_inst5.count_rst_6_cascade_ ;
    wire \b2v_inst5.countZ0Z_8 ;
    wire \b2v_inst5.un2_count_1_cry_7_THRU_CO ;
    wire \b2v_inst5.countZ0Z_8_cascade_ ;
    wire \b2v_inst5.count_0_8 ;
    wire \b2v_inst5.count_rst_10 ;
    wire \b2v_inst5.count_rst_10_cascade_ ;
    wire \b2v_inst5.un2_count_1_axb_4 ;
    wire \b2v_inst5.un2_count_1_cry_3_THRU_CO ;
    wire \b2v_inst5.un2_count_1_axb_4_cascade_ ;
    wire \b2v_inst5.count_0_4 ;
    wire \b2v_inst5.N_390 ;
    wire \b2v_inst5.un2_count_1_cry_12_THRU_CO ;
    wire \b2v_inst5.count_0_sqmuxa ;
    wire \b2v_inst5.count_enZ0 ;
    wire \b2v_inst5.count_rst_1_cascade_ ;
    wire \b2v_inst5.count_0_13 ;
    wire \b2v_inst5.countZ0Z_13 ;
    wire \b2v_inst20.counterZ0Z_11 ;
    wire \b2v_inst20.counterZ0Z_8 ;
    wire \b2v_inst20.counterZ0Z_10 ;
    wire \b2v_inst20.counterZ0Z_9 ;
    wire \b2v_inst20.un4_counter_2_and ;
    wire \b2v_inst20.counterZ0Z_12 ;
    wire \b2v_inst20.counterZ0Z_14 ;
    wire \b2v_inst20.counterZ0Z_15 ;
    wire \b2v_inst20.counterZ0Z_13 ;
    wire \b2v_inst20.un4_counter_3_and ;
    wire \b2v_inst20.counterZ0Z_19 ;
    wire \b2v_inst20.counterZ0Z_16 ;
    wire \b2v_inst20.counterZ0Z_17 ;
    wire \b2v_inst20.counterZ0Z_18 ;
    wire \b2v_inst20.un4_counter_4_and ;
    wire \b2v_inst20.counterZ0Z_23 ;
    wire \b2v_inst20.counterZ0Z_22 ;
    wire \b2v_inst20.counterZ0Z_21 ;
    wire \b2v_inst20.counterZ0Z_20 ;
    wire \b2v_inst20.un4_counter_5_and ;
    wire \b2v_inst20.counterZ0Z_24 ;
    wire \b2v_inst20.counterZ0Z_27 ;
    wire \b2v_inst20.counterZ0Z_25 ;
    wire \b2v_inst20.counterZ0Z_26 ;
    wire \b2v_inst20.un4_counter_6_and ;
    wire \b2v_inst200.curr_stateZ0Z_1_cascade_ ;
    wire N_405;
    wire GPIO_FPGA_PCH_1_c;
    wire \b2v_inst200.count_RNI_0_0 ;
    wire N_405_cascade_;
    wire \b2v_inst200.m6_i_0_cascade_ ;
    wire \b2v_inst200.N_57_cascade_ ;
    wire \b2v_inst200.curr_stateZ0Z_0_cascade_ ;
    wire N_406_cascade_;
    wire \b2v_inst200.N_55 ;
    wire N_406;
    wire \b2v_inst200.curr_state_0_1 ;
    wire \b2v_inst200.N_202_cascade_ ;
    wire HDA_SDO_FPGA_c;
    wire \b2v_inst20.counterZ0Z_29 ;
    wire \b2v_inst20.counterZ0Z_28 ;
    wire \b2v_inst20.counterZ0Z_31 ;
    wire \b2v_inst20.counterZ0Z_30 ;
    wire \b2v_inst20.un4_counter_7_and ;
    wire \b2v_inst200.m11_0_a3_0 ;
    wire \b2v_inst200.N_202 ;
    wire G_2788;
    wire \b2v_inst200.curr_state_0_2 ;
    wire G_2788_cascade_;
    wire SYNTHESIZED_WIRE_47keep;
    wire \b2v_inst200.curr_stateZ0Z_2 ;
    wire \b2v_inst200.curr_stateZ0Z_2_cascade_ ;
    wire \b2v_inst200.HDA_SDO_FPGA_0 ;
    wire \b2v_inst200.curr_stateZ0Z_0 ;
    wire \b2v_inst200.curr_stateZ0Z_1 ;
    wire N_219;
    wire \b2v_inst200.m6_i_0 ;
    wire \b2v_inst200.curr_state_0_0 ;
    wire b2v_inst16_delayed_vddq_pwrgd_en_g;
    wire \b2v_inst6.count_rst_0_cascade_ ;
    wire \b2v_inst6.countZ0Z_1_cascade_ ;
    wire \b2v_inst6.count_3_1 ;
    wire \b2v_inst6.count_rst_1 ;
    wire \b2v_inst6.count_3_2 ;
    wire \b2v_inst6.count_3_6 ;
    wire \b2v_inst6.count_rst_5 ;
    wire \b2v_inst6.countZ0Z_6 ;
    wire \b2v_inst6.countZ0Z_10 ;
    wire \b2v_inst6.countZ0Z_2 ;
    wire \b2v_inst6.countZ0Z_6_cascade_ ;
    wire \b2v_inst6.countZ0Z_1 ;
    wire \b2v_inst6.countZ0Z_12 ;
    wire \b2v_inst6.count_rst_11 ;
    wire \b2v_inst6.count_3_12 ;
    wire \b2v_inst6.countZ0Z_13 ;
    wire \b2v_inst6.count_rst_12 ;
    wire \b2v_inst6.count_3_13 ;
    wire \b2v_inst6.countZ0Z_14 ;
    wire \b2v_inst6.count_rst_13 ;
    wire \b2v_inst6.count_3_14 ;
    wire \b2v_inst6.count_3_15 ;
    wire \b2v_inst6.count_rst_14 ;
    wire \b2v_inst6.countZ0Z_15 ;
    wire V5A_OK_c;
    wire V33A_OK_c;
    wire V1P8A_OK_c;
    wire V105A_OK_c;
    wire SYNTHESIZED_WIRE_26;
    wire \b2v_inst6.count_rst_cascade_ ;
    wire \b2v_inst6.countZ0Z_0_cascade_ ;
    wire \b2v_inst6.count_3_0 ;
    wire \b2v_inst6.un2_count_1_cry_2_THRU_CO ;
    wire \b2v_inst6.count_3_3 ;
    wire FPGA_OSC_0_c_g;
    wire \b2v_inst6.count_en ;
    wire \b2v_inst6.count_0_sqmuxa ;
    wire \b2v_inst6.countZ0Z_5 ;
    wire \b2v_inst6.countZ0Z_3 ;
    wire \b2v_inst6.countZ0Z_4 ;
    wire \b2v_inst6.countZ0Z_0 ;
    wire \b2v_inst6.un12_clk_100khz_10 ;
    wire \b2v_inst6.un12_clk_100khz_9 ;
    wire \b2v_inst6.un12_clk_100khz_11_cascade_ ;
    wire \b2v_inst6.un12_clk_100khz_8 ;
    wire \b2v_inst6.N_1_i ;
    wire \b2v_inst6.N_1_i_cascade_ ;
    wire \b2v_inst6.N_1_i_i ;
    wire _gnd_net_;

    PRE_IO_GBUF FPGA_OSC_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__35651),
            .GLOBALBUFFEROUTPUT(FPGA_OSC_0_c_g));
    IO_PAD FPGA_OSC_ibuf_gb_io_iopad (
            .OE(N__35653),
            .DIN(N__35652),
            .DOUT(N__35651),
            .PACKAGEPIN(FPGA_OSC));
    defparam FPGA_OSC_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam FPGA_OSC_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO FPGA_OSC_ibuf_gb_io_preio (
            .PADOEN(N__35653),
            .PADOUT(N__35652),
            .PADIN(N__35651),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V1P8A_OK_ibuf_iopad (
            .OE(N__35642),
            .DIN(N__35641),
            .DOUT(N__35640),
            .PACKAGEPIN(V1P8A_OK));
    defparam V1P8A_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V1P8A_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V1P8A_OK_ibuf_preio (
            .PADOEN(N__35642),
            .PADOUT(N__35641),
            .PADIN(N__35640),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V1P8A_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V5A_OK_ibuf_iopad (
            .OE(N__35633),
            .DIN(N__35632),
            .DOUT(N__35631),
            .PACKAGEPIN(V5A_OK));
    defparam V5A_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V5A_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V5A_OK_ibuf_preio (
            .PADOEN(N__35633),
            .PADOUT(N__35632),
            .PADIN(N__35631),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V5A_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PCH_PWROK_obuf_iopad (
            .OE(N__35624),
            .DIN(N__35623),
            .DOUT(N__35622),
            .PACKAGEPIN(PCH_PWROK));
    defparam PCH_PWROK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PCH_PWROK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PCH_PWROK_obuf_preio (
            .PADOEN(N__35624),
            .PADOUT(N__35623),
            .PADIN(N__35622),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17640),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCIN_EN_obuf_iopad (
            .OE(N__35615),
            .DIN(N__35614),
            .DOUT(N__35613),
            .PACKAGEPIN(VCCIN_EN));
    defparam VCCIN_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCIN_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCIN_EN_obuf_preio (
            .PADOEN(N__35615),
            .PADOUT(N__35614),
            .PADIN(N__35613),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24954),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33S_OK_ibuf_iopad (
            .OE(N__35606),
            .DIN(N__35605),
            .DOUT(N__35604),
            .PACKAGEPIN(V33S_OK));
    defparam V33S_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V33S_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V33S_OK_ibuf_preio (
            .PADOEN(N__35606),
            .PADOUT(N__35605),
            .PADIN(N__35604),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V33S_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V5S_ENn_obuf_iopad (
            .OE(N__35597),
            .DIN(N__35596),
            .DOUT(N__35595),
            .PACKAGEPIN(V5S_ENn));
    defparam V5S_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V5S_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V5S_ENn_obuf_preio (
            .PADOEN(N__35597),
            .PADOUT(N__35596),
            .PADIN(N__35595),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29685),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SLP_S4n_ibuf_iopad (
            .OE(N__35588),
            .DIN(N__35587),
            .DOUT(N__35586),
            .PACKAGEPIN(SLP_S4n));
    defparam SLP_S4n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SLP_S4n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SLP_S4n_ibuf_preio (
            .PADOEN(N__35588),
            .PADOUT(N__35587),
            .PADIN(N__35586),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SLP_S4n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD HDA_SDO_FPGA_obuf_iopad (
            .OE(N__35579),
            .DIN(N__35578),
            .DOUT(N__35577),
            .PACKAGEPIN(HDA_SDO_FPGA));
    defparam HDA_SDO_FPGA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HDA_SDO_FPGA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HDA_SDO_FPGA_obuf_preio (
            .PADOEN(N__35579),
            .PADOUT(N__35578),
            .PADIN(N__35577),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33505),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VR_READY_VCCINAUX_ibuf_iopad (
            .OE(N__35570),
            .DIN(N__35569),
            .DOUT(N__35568),
            .PACKAGEPIN(VR_READY_VCCINAUX));
    defparam VR_READY_VCCINAUX_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VR_READY_VCCINAUX_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VR_READY_VCCINAUX_ibuf_preio (
            .PADOEN(N__35570),
            .PADOUT(N__35569),
            .PADIN(N__35568),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VR_READY_VCCINAUX_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SLP_S3n_ibuf_iopad (
            .OE(N__35561),
            .DIN(N__35560),
            .DOUT(N__35559),
            .PACKAGEPIN(SLP_S3n));
    defparam SLP_S3n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SLP_S3n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SLP_S3n_ibuf_preio (
            .PADOEN(N__35561),
            .PADOUT(N__35560),
            .PADIN(N__35559),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SLP_S3n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCST_PWRGD_obuf_iopad (
            .OE(N__35552),
            .DIN(N__35551),
            .DOUT(N__35550),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam VCCST_PWRGD_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCST_PWRGD_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCST_PWRGD_obuf_preio (
            .PADOEN(N__35552),
            .PADOUT(N__35551),
            .PADIN(N__35550),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17625),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VPP_OK_ibuf_iopad (
            .OE(N__35543),
            .DIN(N__35542),
            .DOUT(N__35541),
            .PACKAGEPIN(VPP_OK));
    defparam VPP_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VPP_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VPP_OK_ibuf_preio (
            .PADOEN(N__35543),
            .PADOUT(N__35542),
            .PADIN(N__35541),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VPP_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33A_ENn_obuf_iopad (
            .OE(N__35534),
            .DIN(N__35533),
            .DOUT(N__35532),
            .PACKAGEPIN(V33A_ENn));
    defparam V33A_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V33A_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V33A_ENn_obuf_preio (
            .PADOEN(N__35534),
            .PADOUT(N__35533),
            .PADIN(N__35532),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V5S_OK_ibuf_iopad (
            .OE(N__35525),
            .DIN(N__35524),
            .DOUT(N__35523),
            .PACKAGEPIN(V5S_OK));
    defparam V5S_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V5S_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V5S_OK_ibuf_preio (
            .PADOEN(N__35525),
            .PADOUT(N__35524),
            .PADIN(N__35523),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V5S_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33A_OK_ibuf_iopad (
            .OE(N__35516),
            .DIN(N__35515),
            .DOUT(N__35514),
            .PACKAGEPIN(V33A_OK));
    defparam V33A_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V33A_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V33A_OK_ibuf_preio (
            .PADOEN(N__35516),
            .PADOUT(N__35515),
            .PADIN(N__35514),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V33A_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VPP_EN_obuf_iopad (
            .OE(N__35507),
            .DIN(N__35506),
            .DOUT(N__35505),
            .PACKAGEPIN(VPP_EN));
    defparam VPP_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VPP_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VPP_EN_obuf_preio (
            .PADOEN(N__35507),
            .PADOUT(N__35506),
            .PADIN(N__35505),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20290),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PWRBTN_LED_obuf_iopad (
            .OE(N__35498),
            .DIN(N__35497),
            .DOUT(N__35496),
            .PACKAGEPIN(PWRBTN_LED));
    defparam PWRBTN_LED_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PWRBTN_LED_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PWRBTN_LED_obuf_preio (
            .PADOEN(N__35498),
            .PADOUT(N__35497),
            .PADIN(N__35496),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22144),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCIO_OK_ibuf_iopad (
            .OE(N__35489),
            .DIN(N__35488),
            .DOUT(N__35487),
            .PACKAGEPIN(VCCIO_OK));
    defparam VCCIO_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCIO_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VCCIO_OK_ibuf_preio (
            .PADOEN(N__35489),
            .PADOUT(N__35488),
            .PADIN(N__35487),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VCCIO_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33S_ENn_obuf_iopad (
            .OE(N__35480),
            .DIN(N__35479),
            .DOUT(N__35478),
            .PACKAGEPIN(V33S_ENn));
    defparam V33S_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V33S_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V33S_ENn_obuf_preio (
            .PADOEN(N__35480),
            .PADOUT(N__35479),
            .PADIN(N__35478),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29686),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RSMRSTn_obuf_iopad (
            .OE(N__35471),
            .DIN(N__35470),
            .DOUT(N__35469),
            .PACKAGEPIN(RSMRSTn));
    defparam RSMRSTn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RSMRSTn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RSMRSTn_obuf_preio (
            .PADOEN(N__35471),
            .PADOUT(N__35470),
            .PADIN(N__35469),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29119),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V105A_EN_obuf_iopad (
            .OE(N__35462),
            .DIN(N__35461),
            .DOUT(N__35460),
            .PACKAGEPIN(V105A_EN));
    defparam V105A_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V105A_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V105A_EN_obuf_preio (
            .PADOEN(N__35462),
            .PADOUT(N__35461),
            .PADIN(N__35460),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20494),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V1P8A_EN_obuf_iopad (
            .OE(N__35453),
            .DIN(N__35452),
            .DOUT(N__35451),
            .PACKAGEPIN(V1P8A_EN));
    defparam V1P8A_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V1P8A_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V1P8A_EN_obuf_preio (
            .PADOEN(N__35453),
            .PADOUT(N__35452),
            .PADIN(N__35451),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VDDQ_OK_ibuf_iopad (
            .OE(N__35444),
            .DIN(N__35443),
            .DOUT(N__35442),
            .PACKAGEPIN(VDDQ_OK));
    defparam VDDQ_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VDDQ_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VDDQ_OK_ibuf_preio (
            .PADOEN(N__35444),
            .PADOUT(N__35443),
            .PADIN(N__35442),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VDDQ_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCST_ENn_obuf_iopad (
            .OE(N__35435),
            .DIN(N__35434),
            .DOUT(N__35433),
            .PACKAGEPIN(VCCST_ENn));
    defparam VCCST_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCST_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCST_ENn_obuf_preio (
            .PADOEN(N__35435),
            .PADOUT(N__35434),
            .PADIN(N__35433),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25096),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCST_OK_ibuf_iopad (
            .OE(N__35426),
            .DIN(N__35425),
            .DOUT(N__35424),
            .PACKAGEPIN(VCCST_OK));
    defparam VCCST_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCST_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VCCST_OK_ibuf_preio (
            .PADOEN(N__35426),
            .PADOUT(N__35425),
            .PADIN(N__35424),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VCCST_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DSW_PWROK_obuf_iopad (
            .OE(N__35417),
            .DIN(N__35416),
            .DOUT(N__35415),
            .PACKAGEPIN(DSW_PWROK));
    defparam DSW_PWROK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DSW_PWROK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DSW_PWROK_obuf_preio (
            .PADOEN(N__35417),
            .PADOUT(N__35416),
            .PADIN(N__35415),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20493),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SYS_PWROK_obuf_iopad (
            .OE(N__35408),
            .DIN(N__35407),
            .DOUT(N__35406),
            .PACKAGEPIN(SYS_PWROK));
    defparam SYS_PWROK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SYS_PWROK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SYS_PWROK_obuf_preio (
            .PADOEN(N__35408),
            .PADOUT(N__35407),
            .PADIN(N__35406),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17641),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO_FPGA_PCH_5_ibuf_iopad (
            .OE(N__35399),
            .DIN(N__35398),
            .DOUT(N__35397),
            .PACKAGEPIN(GPIO_FPGA_PCH_5));
    defparam GPIO_FPGA_PCH_5_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO_FPGA_PCH_5_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO GPIO_FPGA_PCH_5_ibuf_preio (
            .PADOEN(N__35399),
            .PADOUT(N__35398),
            .PADIN(N__35397),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(GPIO_FPGA_PCH_5_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33DSW_OK_ibuf_iopad (
            .OE(N__35390),
            .DIN(N__35389),
            .DOUT(N__35388),
            .PACKAGEPIN(V33DSW_OK));
    defparam V33DSW_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V33DSW_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V33DSW_OK_ibuf_preio (
            .PADOEN(N__35390),
            .PADOUT(N__35389),
            .PADIN(N__35388),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V33DSW_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V105A_OK_ibuf_iopad (
            .OE(N__35381),
            .DIN(N__35380),
            .DOUT(N__35379),
            .PACKAGEPIN(V105A_OK));
    defparam V105A_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V105A_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V105A_OK_ibuf_preio (
            .PADOEN(N__35381),
            .PADOUT(N__35380),
            .PADIN(N__35379),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V105A_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VR_READY_VCCIN_ibuf_iopad (
            .OE(N__35372),
            .DIN(N__35371),
            .DOUT(N__35370),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam VR_READY_VCCIN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VR_READY_VCCIN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VR_READY_VCCIN_ibuf_preio (
            .PADOEN(N__35372),
            .PADOUT(N__35371),
            .PADIN(N__35370),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VR_READY_VCCIN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VDDQ_EN_obuf_iopad (
            .OE(N__35363),
            .DIN(N__35362),
            .DOUT(N__35361),
            .PACKAGEPIN(VDDQ_EN));
    defparam VDDQ_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VDDQ_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VDDQ_EN_obuf_preio (
            .PADOEN(N__35363),
            .PADOUT(N__35362),
            .PADIN(N__35361),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24994),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO_FPGA_PCH_1_ibuf_iopad (
            .OE(N__35354),
            .DIN(N__35353),
            .DOUT(N__35352),
            .PACKAGEPIN(GPIO_FPGA_PCH_1));
    defparam GPIO_FPGA_PCH_1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO_FPGA_PCH_1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO GPIO_FPGA_PCH_1_ibuf_preio (
            .PADOEN(N__35354),
            .PADOUT(N__35353),
            .PADIN(N__35352),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(GPIO_FPGA_PCH_1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V5A_EN_obuf_iopad (
            .OE(N__35345),
            .DIN(N__35344),
            .DOUT(N__35343),
            .PACKAGEPIN(V5A_EN));
    defparam V5A_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V5A_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V5A_EN_obuf_preio (
            .PADOEN(N__35345),
            .PADOUT(N__35344),
            .PADIN(N__35343),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20125),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCINAUX_EN_obuf_iopad (
            .OE(N__35336),
            .DIN(N__35335),
            .DOUT(N__35334),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam VCCINAUX_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCINAUX_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCINAUX_EN_obuf_preio (
            .PADOEN(N__35336),
            .PADOUT(N__35335),
            .PADIN(N__35334),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24955),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCIO_EN_obuf_iopad (
            .OE(N__35327),
            .DIN(N__35326),
            .DOUT(N__35325),
            .PACKAGEPIN(VCCIO_EN));
    defparam VCCIO_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCIO_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCIO_EN_obuf_preio (
            .PADOEN(N__35327),
            .PADOUT(N__35326),
            .PADIN(N__35325),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20605),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    SRMux I__8172 (
            .O(N__35308),
            .I(N__35304));
    SRMux I__8171 (
            .O(N__35307),
            .I(N__35301));
    LocalMux I__8170 (
            .O(N__35304),
            .I(N__35298));
    LocalMux I__8169 (
            .O(N__35301),
            .I(N__35285));
    IoSpan4Mux I__8168 (
            .O(N__35298),
            .I(N__35285));
    SRMux I__8167 (
            .O(N__35297),
            .I(N__35280));
    InMux I__8166 (
            .O(N__35296),
            .I(N__35280));
    SRMux I__8165 (
            .O(N__35295),
            .I(N__35267));
    SRMux I__8164 (
            .O(N__35294),
            .I(N__35264));
    InMux I__8163 (
            .O(N__35293),
            .I(N__35255));
    InMux I__8162 (
            .O(N__35292),
            .I(N__35255));
    InMux I__8161 (
            .O(N__35291),
            .I(N__35255));
    InMux I__8160 (
            .O(N__35290),
            .I(N__35255));
    Span4Mux_s1_v I__8159 (
            .O(N__35285),
            .I(N__35250));
    LocalMux I__8158 (
            .O(N__35280),
            .I(N__35250));
    InMux I__8157 (
            .O(N__35279),
            .I(N__35239));
    InMux I__8156 (
            .O(N__35278),
            .I(N__35239));
    InMux I__8155 (
            .O(N__35277),
            .I(N__35239));
    InMux I__8154 (
            .O(N__35276),
            .I(N__35239));
    InMux I__8153 (
            .O(N__35275),
            .I(N__35239));
    InMux I__8152 (
            .O(N__35274),
            .I(N__35234));
    InMux I__8151 (
            .O(N__35273),
            .I(N__35234));
    InMux I__8150 (
            .O(N__35272),
            .I(N__35229));
    InMux I__8149 (
            .O(N__35271),
            .I(N__35229));
    SRMux I__8148 (
            .O(N__35270),
            .I(N__35219));
    LocalMux I__8147 (
            .O(N__35267),
            .I(N__35214));
    LocalMux I__8146 (
            .O(N__35264),
            .I(N__35214));
    LocalMux I__8145 (
            .O(N__35255),
            .I(N__35211));
    Span4Mux_v I__8144 (
            .O(N__35250),
            .I(N__35206));
    LocalMux I__8143 (
            .O(N__35239),
            .I(N__35206));
    LocalMux I__8142 (
            .O(N__35234),
            .I(N__35196));
    LocalMux I__8141 (
            .O(N__35229),
            .I(N__35196));
    SRMux I__8140 (
            .O(N__35228),
            .I(N__35193));
    InMux I__8139 (
            .O(N__35227),
            .I(N__35186));
    InMux I__8138 (
            .O(N__35226),
            .I(N__35186));
    InMux I__8137 (
            .O(N__35225),
            .I(N__35186));
    InMux I__8136 (
            .O(N__35224),
            .I(N__35179));
    InMux I__8135 (
            .O(N__35223),
            .I(N__35179));
    InMux I__8134 (
            .O(N__35222),
            .I(N__35179));
    LocalMux I__8133 (
            .O(N__35219),
            .I(N__35175));
    Span4Mux_v I__8132 (
            .O(N__35214),
            .I(N__35168));
    Span4Mux_v I__8131 (
            .O(N__35211),
            .I(N__35168));
    Span4Mux_s1_v I__8130 (
            .O(N__35206),
            .I(N__35168));
    InMux I__8129 (
            .O(N__35205),
            .I(N__35157));
    InMux I__8128 (
            .O(N__35204),
            .I(N__35157));
    InMux I__8127 (
            .O(N__35203),
            .I(N__35157));
    InMux I__8126 (
            .O(N__35202),
            .I(N__35157));
    InMux I__8125 (
            .O(N__35201),
            .I(N__35157));
    Span4Mux_s2_h I__8124 (
            .O(N__35196),
            .I(N__35154));
    LocalMux I__8123 (
            .O(N__35193),
            .I(N__35147));
    LocalMux I__8122 (
            .O(N__35186),
            .I(N__35147));
    LocalMux I__8121 (
            .O(N__35179),
            .I(N__35147));
    InMux I__8120 (
            .O(N__35178),
            .I(N__35144));
    Odrv4 I__8119 (
            .O(N__35175),
            .I(\b2v_inst6.count_0_sqmuxa ));
    Odrv4 I__8118 (
            .O(N__35168),
            .I(\b2v_inst6.count_0_sqmuxa ));
    LocalMux I__8117 (
            .O(N__35157),
            .I(\b2v_inst6.count_0_sqmuxa ));
    Odrv4 I__8116 (
            .O(N__35154),
            .I(\b2v_inst6.count_0_sqmuxa ));
    Odrv4 I__8115 (
            .O(N__35147),
            .I(\b2v_inst6.count_0_sqmuxa ));
    LocalMux I__8114 (
            .O(N__35144),
            .I(\b2v_inst6.count_0_sqmuxa ));
    InMux I__8113 (
            .O(N__35131),
            .I(N__35127));
    CascadeMux I__8112 (
            .O(N__35130),
            .I(N__35122));
    LocalMux I__8111 (
            .O(N__35127),
            .I(N__35119));
    InMux I__8110 (
            .O(N__35126),
            .I(N__35116));
    InMux I__8109 (
            .O(N__35125),
            .I(N__35113));
    InMux I__8108 (
            .O(N__35122),
            .I(N__35110));
    Span4Mux_v I__8107 (
            .O(N__35119),
            .I(N__35107));
    LocalMux I__8106 (
            .O(N__35116),
            .I(N__35104));
    LocalMux I__8105 (
            .O(N__35113),
            .I(\b2v_inst6.countZ0Z_5 ));
    LocalMux I__8104 (
            .O(N__35110),
            .I(\b2v_inst6.countZ0Z_5 ));
    Odrv4 I__8103 (
            .O(N__35107),
            .I(\b2v_inst6.countZ0Z_5 ));
    Odrv4 I__8102 (
            .O(N__35104),
            .I(\b2v_inst6.countZ0Z_5 ));
    CascadeMux I__8101 (
            .O(N__35095),
            .I(N__35089));
    CascadeMux I__8100 (
            .O(N__35094),
            .I(N__35086));
    InMux I__8099 (
            .O(N__35093),
            .I(N__35083));
    InMux I__8098 (
            .O(N__35092),
            .I(N__35080));
    InMux I__8097 (
            .O(N__35089),
            .I(N__35077));
    InMux I__8096 (
            .O(N__35086),
            .I(N__35074));
    LocalMux I__8095 (
            .O(N__35083),
            .I(N__35071));
    LocalMux I__8094 (
            .O(N__35080),
            .I(\b2v_inst6.countZ0Z_3 ));
    LocalMux I__8093 (
            .O(N__35077),
            .I(\b2v_inst6.countZ0Z_3 ));
    LocalMux I__8092 (
            .O(N__35074),
            .I(\b2v_inst6.countZ0Z_3 ));
    Odrv4 I__8091 (
            .O(N__35071),
            .I(\b2v_inst6.countZ0Z_3 ));
    CascadeMux I__8090 (
            .O(N__35062),
            .I(N__35059));
    InMux I__8089 (
            .O(N__35059),
            .I(N__35055));
    InMux I__8088 (
            .O(N__35058),
            .I(N__35051));
    LocalMux I__8087 (
            .O(N__35055),
            .I(N__35048));
    CascadeMux I__8086 (
            .O(N__35054),
            .I(N__35045));
    LocalMux I__8085 (
            .O(N__35051),
            .I(N__35042));
    Span4Mux_s3_h I__8084 (
            .O(N__35048),
            .I(N__35039));
    InMux I__8083 (
            .O(N__35045),
            .I(N__35036));
    Span4Mux_s2_h I__8082 (
            .O(N__35042),
            .I(N__35033));
    Odrv4 I__8081 (
            .O(N__35039),
            .I(\b2v_inst6.countZ0Z_4 ));
    LocalMux I__8080 (
            .O(N__35036),
            .I(\b2v_inst6.countZ0Z_4 ));
    Odrv4 I__8079 (
            .O(N__35033),
            .I(\b2v_inst6.countZ0Z_4 ));
    CascadeMux I__8078 (
            .O(N__35026),
            .I(N__35022));
    InMux I__8077 (
            .O(N__35025),
            .I(N__35017));
    InMux I__8076 (
            .O(N__35022),
            .I(N__35013));
    InMux I__8075 (
            .O(N__35021),
            .I(N__35008));
    InMux I__8074 (
            .O(N__35020),
            .I(N__35008));
    LocalMux I__8073 (
            .O(N__35017),
            .I(N__35005));
    InMux I__8072 (
            .O(N__35016),
            .I(N__35002));
    LocalMux I__8071 (
            .O(N__35013),
            .I(N__34999));
    LocalMux I__8070 (
            .O(N__35008),
            .I(N__34996));
    Odrv4 I__8069 (
            .O(N__35005),
            .I(\b2v_inst6.countZ0Z_0 ));
    LocalMux I__8068 (
            .O(N__35002),
            .I(\b2v_inst6.countZ0Z_0 ));
    Odrv4 I__8067 (
            .O(N__34999),
            .I(\b2v_inst6.countZ0Z_0 ));
    Odrv12 I__8066 (
            .O(N__34996),
            .I(\b2v_inst6.countZ0Z_0 ));
    InMux I__8065 (
            .O(N__34987),
            .I(N__34984));
    LocalMux I__8064 (
            .O(N__34984),
            .I(\b2v_inst6.un12_clk_100khz_10 ));
    InMux I__8063 (
            .O(N__34981),
            .I(N__34978));
    LocalMux I__8062 (
            .O(N__34978),
            .I(N__34975));
    Odrv4 I__8061 (
            .O(N__34975),
            .I(\b2v_inst6.un12_clk_100khz_9 ));
    CascadeMux I__8060 (
            .O(N__34972),
            .I(\b2v_inst6.un12_clk_100khz_11_cascade_ ));
    InMux I__8059 (
            .O(N__34969),
            .I(N__34966));
    LocalMux I__8058 (
            .O(N__34966),
            .I(N__34963));
    Odrv4 I__8057 (
            .O(N__34963),
            .I(\b2v_inst6.un12_clk_100khz_8 ));
    InMux I__8056 (
            .O(N__34960),
            .I(N__34954));
    InMux I__8055 (
            .O(N__34959),
            .I(N__34954));
    LocalMux I__8054 (
            .O(N__34954),
            .I(N__34951));
    Span4Mux_h I__8053 (
            .O(N__34951),
            .I(N__34948));
    Odrv4 I__8052 (
            .O(N__34948),
            .I(\b2v_inst6.N_1_i ));
    CascadeMux I__8051 (
            .O(N__34945),
            .I(\b2v_inst6.N_1_i_cascade_ ));
    InMux I__8050 (
            .O(N__34942),
            .I(N__34930));
    InMux I__8049 (
            .O(N__34941),
            .I(N__34930));
    InMux I__8048 (
            .O(N__34940),
            .I(N__34917));
    InMux I__8047 (
            .O(N__34939),
            .I(N__34917));
    InMux I__8046 (
            .O(N__34938),
            .I(N__34917));
    InMux I__8045 (
            .O(N__34937),
            .I(N__34917));
    InMux I__8044 (
            .O(N__34936),
            .I(N__34917));
    InMux I__8043 (
            .O(N__34935),
            .I(N__34911));
    LocalMux I__8042 (
            .O(N__34930),
            .I(N__34908));
    CascadeMux I__8041 (
            .O(N__34929),
            .I(N__34905));
    CascadeMux I__8040 (
            .O(N__34928),
            .I(N__34900));
    LocalMux I__8039 (
            .O(N__34917),
            .I(N__34897));
    InMux I__8038 (
            .O(N__34916),
            .I(N__34891));
    InMux I__8037 (
            .O(N__34915),
            .I(N__34886));
    InMux I__8036 (
            .O(N__34914),
            .I(N__34886));
    LocalMux I__8035 (
            .O(N__34911),
            .I(N__34881));
    Span4Mux_v I__8034 (
            .O(N__34908),
            .I(N__34881));
    InMux I__8033 (
            .O(N__34905),
            .I(N__34872));
    InMux I__8032 (
            .O(N__34904),
            .I(N__34872));
    InMux I__8031 (
            .O(N__34903),
            .I(N__34872));
    InMux I__8030 (
            .O(N__34900),
            .I(N__34872));
    Span4Mux_h I__8029 (
            .O(N__34897),
            .I(N__34869));
    InMux I__8028 (
            .O(N__34896),
            .I(N__34862));
    InMux I__8027 (
            .O(N__34895),
            .I(N__34862));
    InMux I__8026 (
            .O(N__34894),
            .I(N__34862));
    LocalMux I__8025 (
            .O(N__34891),
            .I(\b2v_inst6.N_1_i_i ));
    LocalMux I__8024 (
            .O(N__34886),
            .I(\b2v_inst6.N_1_i_i ));
    Odrv4 I__8023 (
            .O(N__34881),
            .I(\b2v_inst6.N_1_i_i ));
    LocalMux I__8022 (
            .O(N__34872),
            .I(\b2v_inst6.N_1_i_i ));
    Odrv4 I__8021 (
            .O(N__34869),
            .I(\b2v_inst6.N_1_i_i ));
    LocalMux I__8020 (
            .O(N__34862),
            .I(\b2v_inst6.N_1_i_i ));
    InMux I__8019 (
            .O(N__34849),
            .I(N__34845));
    InMux I__8018 (
            .O(N__34848),
            .I(N__34842));
    LocalMux I__8017 (
            .O(N__34845),
            .I(\b2v_inst6.countZ0Z_14 ));
    LocalMux I__8016 (
            .O(N__34842),
            .I(\b2v_inst6.countZ0Z_14 ));
    InMux I__8015 (
            .O(N__34837),
            .I(N__34831));
    InMux I__8014 (
            .O(N__34836),
            .I(N__34831));
    LocalMux I__8013 (
            .O(N__34831),
            .I(\b2v_inst6.count_rst_13 ));
    InMux I__8012 (
            .O(N__34828),
            .I(N__34825));
    LocalMux I__8011 (
            .O(N__34825),
            .I(\b2v_inst6.count_3_14 ));
    InMux I__8010 (
            .O(N__34822),
            .I(N__34819));
    LocalMux I__8009 (
            .O(N__34819),
            .I(\b2v_inst6.count_3_15 ));
    InMux I__8008 (
            .O(N__34816),
            .I(N__34812));
    InMux I__8007 (
            .O(N__34815),
            .I(N__34809));
    LocalMux I__8006 (
            .O(N__34812),
            .I(\b2v_inst6.count_rst_14 ));
    LocalMux I__8005 (
            .O(N__34809),
            .I(\b2v_inst6.count_rst_14 ));
    CascadeMux I__8004 (
            .O(N__34804),
            .I(N__34800));
    InMux I__8003 (
            .O(N__34803),
            .I(N__34797));
    InMux I__8002 (
            .O(N__34800),
            .I(N__34794));
    LocalMux I__8001 (
            .O(N__34797),
            .I(\b2v_inst6.countZ0Z_15 ));
    LocalMux I__8000 (
            .O(N__34794),
            .I(\b2v_inst6.countZ0Z_15 ));
    InMux I__7999 (
            .O(N__34789),
            .I(N__34786));
    LocalMux I__7998 (
            .O(N__34786),
            .I(V5A_OK_c));
    InMux I__7997 (
            .O(N__34783),
            .I(N__34780));
    LocalMux I__7996 (
            .O(N__34780),
            .I(V33A_OK_c));
    CascadeMux I__7995 (
            .O(N__34777),
            .I(N__34774));
    InMux I__7994 (
            .O(N__34774),
            .I(N__34771));
    LocalMux I__7993 (
            .O(N__34771),
            .I(V1P8A_OK_c));
    InMux I__7992 (
            .O(N__34768),
            .I(N__34765));
    LocalMux I__7991 (
            .O(N__34765),
            .I(N__34762));
    IoSpan4Mux I__7990 (
            .O(N__34762),
            .I(N__34759));
    Odrv4 I__7989 (
            .O(N__34759),
            .I(V105A_OK_c));
    InMux I__7988 (
            .O(N__34756),
            .I(N__34744));
    InMux I__7987 (
            .O(N__34755),
            .I(N__34744));
    InMux I__7986 (
            .O(N__34754),
            .I(N__34744));
    InMux I__7985 (
            .O(N__34753),
            .I(N__34744));
    LocalMux I__7984 (
            .O(N__34744),
            .I(N__34740));
    InMux I__7983 (
            .O(N__34743),
            .I(N__34737));
    Span12Mux_v I__7982 (
            .O(N__34740),
            .I(N__34732));
    LocalMux I__7981 (
            .O(N__34737),
            .I(N__34732));
    Odrv12 I__7980 (
            .O(N__34732),
            .I(SYNTHESIZED_WIRE_26));
    CascadeMux I__7979 (
            .O(N__34729),
            .I(\b2v_inst6.count_rst_cascade_ ));
    CascadeMux I__7978 (
            .O(N__34726),
            .I(\b2v_inst6.countZ0Z_0_cascade_ ));
    InMux I__7977 (
            .O(N__34723),
            .I(N__34720));
    LocalMux I__7976 (
            .O(N__34720),
            .I(\b2v_inst6.count_3_0 ));
    InMux I__7975 (
            .O(N__34717),
            .I(N__34713));
    InMux I__7974 (
            .O(N__34716),
            .I(N__34710));
    LocalMux I__7973 (
            .O(N__34713),
            .I(N__34707));
    LocalMux I__7972 (
            .O(N__34710),
            .I(N__34704));
    Odrv4 I__7971 (
            .O(N__34707),
            .I(\b2v_inst6.un2_count_1_cry_2_THRU_CO ));
    Odrv4 I__7970 (
            .O(N__34704),
            .I(\b2v_inst6.un2_count_1_cry_2_THRU_CO ));
    InMux I__7969 (
            .O(N__34699),
            .I(N__34696));
    LocalMux I__7968 (
            .O(N__34696),
            .I(N__34693));
    Odrv4 I__7967 (
            .O(N__34693),
            .I(\b2v_inst6.count_3_3 ));
    ClkMux I__7966 (
            .O(N__34690),
            .I(N__34441));
    ClkMux I__7965 (
            .O(N__34689),
            .I(N__34441));
    ClkMux I__7964 (
            .O(N__34688),
            .I(N__34441));
    ClkMux I__7963 (
            .O(N__34687),
            .I(N__34441));
    ClkMux I__7962 (
            .O(N__34686),
            .I(N__34441));
    ClkMux I__7961 (
            .O(N__34685),
            .I(N__34441));
    ClkMux I__7960 (
            .O(N__34684),
            .I(N__34441));
    ClkMux I__7959 (
            .O(N__34683),
            .I(N__34441));
    ClkMux I__7958 (
            .O(N__34682),
            .I(N__34441));
    ClkMux I__7957 (
            .O(N__34681),
            .I(N__34441));
    ClkMux I__7956 (
            .O(N__34680),
            .I(N__34441));
    ClkMux I__7955 (
            .O(N__34679),
            .I(N__34441));
    ClkMux I__7954 (
            .O(N__34678),
            .I(N__34441));
    ClkMux I__7953 (
            .O(N__34677),
            .I(N__34441));
    ClkMux I__7952 (
            .O(N__34676),
            .I(N__34441));
    ClkMux I__7951 (
            .O(N__34675),
            .I(N__34441));
    ClkMux I__7950 (
            .O(N__34674),
            .I(N__34441));
    ClkMux I__7949 (
            .O(N__34673),
            .I(N__34441));
    ClkMux I__7948 (
            .O(N__34672),
            .I(N__34441));
    ClkMux I__7947 (
            .O(N__34671),
            .I(N__34441));
    ClkMux I__7946 (
            .O(N__34670),
            .I(N__34441));
    ClkMux I__7945 (
            .O(N__34669),
            .I(N__34441));
    ClkMux I__7944 (
            .O(N__34668),
            .I(N__34441));
    ClkMux I__7943 (
            .O(N__34667),
            .I(N__34441));
    ClkMux I__7942 (
            .O(N__34666),
            .I(N__34441));
    ClkMux I__7941 (
            .O(N__34665),
            .I(N__34441));
    ClkMux I__7940 (
            .O(N__34664),
            .I(N__34441));
    ClkMux I__7939 (
            .O(N__34663),
            .I(N__34441));
    ClkMux I__7938 (
            .O(N__34662),
            .I(N__34441));
    ClkMux I__7937 (
            .O(N__34661),
            .I(N__34441));
    ClkMux I__7936 (
            .O(N__34660),
            .I(N__34441));
    ClkMux I__7935 (
            .O(N__34659),
            .I(N__34441));
    ClkMux I__7934 (
            .O(N__34658),
            .I(N__34441));
    ClkMux I__7933 (
            .O(N__34657),
            .I(N__34441));
    ClkMux I__7932 (
            .O(N__34656),
            .I(N__34441));
    ClkMux I__7931 (
            .O(N__34655),
            .I(N__34441));
    ClkMux I__7930 (
            .O(N__34654),
            .I(N__34441));
    ClkMux I__7929 (
            .O(N__34653),
            .I(N__34441));
    ClkMux I__7928 (
            .O(N__34652),
            .I(N__34441));
    ClkMux I__7927 (
            .O(N__34651),
            .I(N__34441));
    ClkMux I__7926 (
            .O(N__34650),
            .I(N__34441));
    ClkMux I__7925 (
            .O(N__34649),
            .I(N__34441));
    ClkMux I__7924 (
            .O(N__34648),
            .I(N__34441));
    ClkMux I__7923 (
            .O(N__34647),
            .I(N__34441));
    ClkMux I__7922 (
            .O(N__34646),
            .I(N__34441));
    ClkMux I__7921 (
            .O(N__34645),
            .I(N__34441));
    ClkMux I__7920 (
            .O(N__34644),
            .I(N__34441));
    ClkMux I__7919 (
            .O(N__34643),
            .I(N__34441));
    ClkMux I__7918 (
            .O(N__34642),
            .I(N__34441));
    ClkMux I__7917 (
            .O(N__34641),
            .I(N__34441));
    ClkMux I__7916 (
            .O(N__34640),
            .I(N__34441));
    ClkMux I__7915 (
            .O(N__34639),
            .I(N__34441));
    ClkMux I__7914 (
            .O(N__34638),
            .I(N__34441));
    ClkMux I__7913 (
            .O(N__34637),
            .I(N__34441));
    ClkMux I__7912 (
            .O(N__34636),
            .I(N__34441));
    ClkMux I__7911 (
            .O(N__34635),
            .I(N__34441));
    ClkMux I__7910 (
            .O(N__34634),
            .I(N__34441));
    ClkMux I__7909 (
            .O(N__34633),
            .I(N__34441));
    ClkMux I__7908 (
            .O(N__34632),
            .I(N__34441));
    ClkMux I__7907 (
            .O(N__34631),
            .I(N__34441));
    ClkMux I__7906 (
            .O(N__34630),
            .I(N__34441));
    ClkMux I__7905 (
            .O(N__34629),
            .I(N__34441));
    ClkMux I__7904 (
            .O(N__34628),
            .I(N__34441));
    ClkMux I__7903 (
            .O(N__34627),
            .I(N__34441));
    ClkMux I__7902 (
            .O(N__34626),
            .I(N__34441));
    ClkMux I__7901 (
            .O(N__34625),
            .I(N__34441));
    ClkMux I__7900 (
            .O(N__34624),
            .I(N__34441));
    ClkMux I__7899 (
            .O(N__34623),
            .I(N__34441));
    ClkMux I__7898 (
            .O(N__34622),
            .I(N__34441));
    ClkMux I__7897 (
            .O(N__34621),
            .I(N__34441));
    ClkMux I__7896 (
            .O(N__34620),
            .I(N__34441));
    ClkMux I__7895 (
            .O(N__34619),
            .I(N__34441));
    ClkMux I__7894 (
            .O(N__34618),
            .I(N__34441));
    ClkMux I__7893 (
            .O(N__34617),
            .I(N__34441));
    ClkMux I__7892 (
            .O(N__34616),
            .I(N__34441));
    ClkMux I__7891 (
            .O(N__34615),
            .I(N__34441));
    ClkMux I__7890 (
            .O(N__34614),
            .I(N__34441));
    ClkMux I__7889 (
            .O(N__34613),
            .I(N__34441));
    ClkMux I__7888 (
            .O(N__34612),
            .I(N__34441));
    ClkMux I__7887 (
            .O(N__34611),
            .I(N__34441));
    ClkMux I__7886 (
            .O(N__34610),
            .I(N__34441));
    ClkMux I__7885 (
            .O(N__34609),
            .I(N__34441));
    ClkMux I__7884 (
            .O(N__34608),
            .I(N__34441));
    GlobalMux I__7883 (
            .O(N__34441),
            .I(N__34438));
    gio2CtrlBuf I__7882 (
            .O(N__34438),
            .I(FPGA_OSC_0_c_g));
    CEMux I__7881 (
            .O(N__34435),
            .I(N__34431));
    CEMux I__7880 (
            .O(N__34434),
            .I(N__34422));
    LocalMux I__7879 (
            .O(N__34431),
            .I(N__34411));
    CEMux I__7878 (
            .O(N__34430),
            .I(N__34408));
    CEMux I__7877 (
            .O(N__34429),
            .I(N__34405));
    InMux I__7876 (
            .O(N__34428),
            .I(N__34396));
    InMux I__7875 (
            .O(N__34427),
            .I(N__34396));
    InMux I__7874 (
            .O(N__34426),
            .I(N__34396));
    InMux I__7873 (
            .O(N__34425),
            .I(N__34396));
    LocalMux I__7872 (
            .O(N__34422),
            .I(N__34393));
    CEMux I__7871 (
            .O(N__34421),
            .I(N__34390));
    CEMux I__7870 (
            .O(N__34420),
            .I(N__34387));
    InMux I__7869 (
            .O(N__34419),
            .I(N__34382));
    InMux I__7868 (
            .O(N__34418),
            .I(N__34382));
    CEMux I__7867 (
            .O(N__34417),
            .I(N__34373));
    InMux I__7866 (
            .O(N__34416),
            .I(N__34373));
    InMux I__7865 (
            .O(N__34415),
            .I(N__34373));
    InMux I__7864 (
            .O(N__34414),
            .I(N__34373));
    Span4Mux_s3_h I__7863 (
            .O(N__34411),
            .I(N__34365));
    LocalMux I__7862 (
            .O(N__34408),
            .I(N__34358));
    LocalMux I__7861 (
            .O(N__34405),
            .I(N__34358));
    LocalMux I__7860 (
            .O(N__34396),
            .I(N__34358));
    Span4Mux_s1_v I__7859 (
            .O(N__34393),
            .I(N__34353));
    LocalMux I__7858 (
            .O(N__34390),
            .I(N__34353));
    LocalMux I__7857 (
            .O(N__34387),
            .I(N__34350));
    LocalMux I__7856 (
            .O(N__34382),
            .I(N__34347));
    LocalMux I__7855 (
            .O(N__34373),
            .I(N__34342));
    InMux I__7854 (
            .O(N__34372),
            .I(N__34333));
    InMux I__7853 (
            .O(N__34371),
            .I(N__34333));
    InMux I__7852 (
            .O(N__34370),
            .I(N__34333));
    InMux I__7851 (
            .O(N__34369),
            .I(N__34333));
    InMux I__7850 (
            .O(N__34368),
            .I(N__34330));
    Span4Mux_h I__7849 (
            .O(N__34365),
            .I(N__34325));
    Span4Mux_s3_h I__7848 (
            .O(N__34358),
            .I(N__34325));
    Span4Mux_s1_h I__7847 (
            .O(N__34353),
            .I(N__34318));
    Span4Mux_s1_h I__7846 (
            .O(N__34350),
            .I(N__34318));
    Span4Mux_s1_v I__7845 (
            .O(N__34347),
            .I(N__34318));
    InMux I__7844 (
            .O(N__34346),
            .I(N__34313));
    InMux I__7843 (
            .O(N__34345),
            .I(N__34313));
    Span4Mux_s3_h I__7842 (
            .O(N__34342),
            .I(N__34310));
    LocalMux I__7841 (
            .O(N__34333),
            .I(N__34305));
    LocalMux I__7840 (
            .O(N__34330),
            .I(N__34305));
    Odrv4 I__7839 (
            .O(N__34325),
            .I(\b2v_inst6.count_en ));
    Odrv4 I__7838 (
            .O(N__34318),
            .I(\b2v_inst6.count_en ));
    LocalMux I__7837 (
            .O(N__34313),
            .I(\b2v_inst6.count_en ));
    Odrv4 I__7836 (
            .O(N__34310),
            .I(\b2v_inst6.count_en ));
    Odrv12 I__7835 (
            .O(N__34305),
            .I(\b2v_inst6.count_en ));
    CascadeMux I__7834 (
            .O(N__34294),
            .I(\b2v_inst6.countZ0Z_1_cascade_ ));
    InMux I__7833 (
            .O(N__34291),
            .I(N__34288));
    LocalMux I__7832 (
            .O(N__34288),
            .I(\b2v_inst6.count_3_1 ));
    InMux I__7831 (
            .O(N__34285),
            .I(N__34279));
    InMux I__7830 (
            .O(N__34284),
            .I(N__34279));
    LocalMux I__7829 (
            .O(N__34279),
            .I(\b2v_inst6.count_rst_1 ));
    InMux I__7828 (
            .O(N__34276),
            .I(N__34273));
    LocalMux I__7827 (
            .O(N__34273),
            .I(\b2v_inst6.count_3_2 ));
    InMux I__7826 (
            .O(N__34270),
            .I(N__34267));
    LocalMux I__7825 (
            .O(N__34267),
            .I(\b2v_inst6.count_3_6 ));
    InMux I__7824 (
            .O(N__34264),
            .I(N__34258));
    InMux I__7823 (
            .O(N__34263),
            .I(N__34258));
    LocalMux I__7822 (
            .O(N__34258),
            .I(\b2v_inst6.count_rst_5 ));
    InMux I__7821 (
            .O(N__34255),
            .I(N__34252));
    LocalMux I__7820 (
            .O(N__34252),
            .I(\b2v_inst6.countZ0Z_6 ));
    InMux I__7819 (
            .O(N__34249),
            .I(N__34246));
    LocalMux I__7818 (
            .O(N__34246),
            .I(N__34243));
    Span4Mux_s0_h I__7817 (
            .O(N__34243),
            .I(N__34239));
    InMux I__7816 (
            .O(N__34242),
            .I(N__34236));
    Odrv4 I__7815 (
            .O(N__34239),
            .I(\b2v_inst6.countZ0Z_10 ));
    LocalMux I__7814 (
            .O(N__34236),
            .I(\b2v_inst6.countZ0Z_10 ));
    InMux I__7813 (
            .O(N__34231),
            .I(N__34227));
    InMux I__7812 (
            .O(N__34230),
            .I(N__34224));
    LocalMux I__7811 (
            .O(N__34227),
            .I(\b2v_inst6.countZ0Z_2 ));
    LocalMux I__7810 (
            .O(N__34224),
            .I(\b2v_inst6.countZ0Z_2 ));
    CascadeMux I__7809 (
            .O(N__34219),
            .I(\b2v_inst6.countZ0Z_6_cascade_ ));
    InMux I__7808 (
            .O(N__34216),
            .I(N__34209));
    InMux I__7807 (
            .O(N__34215),
            .I(N__34209));
    InMux I__7806 (
            .O(N__34214),
            .I(N__34206));
    LocalMux I__7805 (
            .O(N__34209),
            .I(\b2v_inst6.countZ0Z_1 ));
    LocalMux I__7804 (
            .O(N__34206),
            .I(\b2v_inst6.countZ0Z_1 ));
    InMux I__7803 (
            .O(N__34201),
            .I(N__34197));
    InMux I__7802 (
            .O(N__34200),
            .I(N__34194));
    LocalMux I__7801 (
            .O(N__34197),
            .I(\b2v_inst6.countZ0Z_12 ));
    LocalMux I__7800 (
            .O(N__34194),
            .I(\b2v_inst6.countZ0Z_12 ));
    InMux I__7799 (
            .O(N__34189),
            .I(N__34183));
    InMux I__7798 (
            .O(N__34188),
            .I(N__34183));
    LocalMux I__7797 (
            .O(N__34183),
            .I(\b2v_inst6.count_rst_11 ));
    InMux I__7796 (
            .O(N__34180),
            .I(N__34177));
    LocalMux I__7795 (
            .O(N__34177),
            .I(\b2v_inst6.count_3_12 ));
    InMux I__7794 (
            .O(N__34174),
            .I(N__34170));
    InMux I__7793 (
            .O(N__34173),
            .I(N__34167));
    LocalMux I__7792 (
            .O(N__34170),
            .I(\b2v_inst6.countZ0Z_13 ));
    LocalMux I__7791 (
            .O(N__34167),
            .I(\b2v_inst6.countZ0Z_13 ));
    InMux I__7790 (
            .O(N__34162),
            .I(N__34156));
    InMux I__7789 (
            .O(N__34161),
            .I(N__34156));
    LocalMux I__7788 (
            .O(N__34156),
            .I(\b2v_inst6.count_rst_12 ));
    InMux I__7787 (
            .O(N__34153),
            .I(N__34150));
    LocalMux I__7786 (
            .O(N__34150),
            .I(\b2v_inst6.count_3_13 ));
    InMux I__7785 (
            .O(N__34147),
            .I(N__34142));
    InMux I__7784 (
            .O(N__34146),
            .I(N__34139));
    InMux I__7783 (
            .O(N__34145),
            .I(N__34136));
    LocalMux I__7782 (
            .O(N__34142),
            .I(N__34129));
    LocalMux I__7781 (
            .O(N__34139),
            .I(N__34129));
    LocalMux I__7780 (
            .O(N__34136),
            .I(N__34129));
    Span12Mux_s9_v I__7779 (
            .O(N__34129),
            .I(N__34126));
    Odrv12 I__7778 (
            .O(N__34126),
            .I(\b2v_inst200.m11_0_a3_0 ));
    CascadeMux I__7777 (
            .O(N__34123),
            .I(N__34120));
    InMux I__7776 (
            .O(N__34120),
            .I(N__34117));
    LocalMux I__7775 (
            .O(N__34117),
            .I(\b2v_inst200.N_202 ));
    InMux I__7774 (
            .O(N__34114),
            .I(N__34111));
    LocalMux I__7773 (
            .O(N__34111),
            .I(N__34108));
    Odrv4 I__7772 (
            .O(N__34108),
            .I(G_2788));
    InMux I__7771 (
            .O(N__34105),
            .I(N__34102));
    LocalMux I__7770 (
            .O(N__34102),
            .I(N__34099));
    Odrv4 I__7769 (
            .O(N__34099),
            .I(\b2v_inst200.curr_state_0_2 ));
    CascadeMux I__7768 (
            .O(N__34096),
            .I(G_2788_cascade_));
    InMux I__7767 (
            .O(N__34093),
            .I(N__34080));
    InMux I__7766 (
            .O(N__34092),
            .I(N__34080));
    CascadeMux I__7765 (
            .O(N__34091),
            .I(N__34066));
    InMux I__7764 (
            .O(N__34090),
            .I(N__34061));
    InMux I__7763 (
            .O(N__34089),
            .I(N__34041));
    InMux I__7762 (
            .O(N__34088),
            .I(N__34041));
    InMux I__7761 (
            .O(N__34087),
            .I(N__34041));
    InMux I__7760 (
            .O(N__34086),
            .I(N__34041));
    CascadeMux I__7759 (
            .O(N__34085),
            .I(N__34038));
    LocalMux I__7758 (
            .O(N__34080),
            .I(N__34033));
    InMux I__7757 (
            .O(N__34079),
            .I(N__34024));
    InMux I__7756 (
            .O(N__34078),
            .I(N__34024));
    InMux I__7755 (
            .O(N__34077),
            .I(N__34024));
    InMux I__7754 (
            .O(N__34076),
            .I(N__34024));
    InMux I__7753 (
            .O(N__34075),
            .I(N__34017));
    InMux I__7752 (
            .O(N__34074),
            .I(N__34017));
    InMux I__7751 (
            .O(N__34073),
            .I(N__34017));
    InMux I__7750 (
            .O(N__34072),
            .I(N__34012));
    InMux I__7749 (
            .O(N__34071),
            .I(N__34012));
    InMux I__7748 (
            .O(N__34070),
            .I(N__34007));
    InMux I__7747 (
            .O(N__34069),
            .I(N__34007));
    InMux I__7746 (
            .O(N__34066),
            .I(N__34003));
    InMux I__7745 (
            .O(N__34065),
            .I(N__33998));
    InMux I__7744 (
            .O(N__34064),
            .I(N__33998));
    LocalMux I__7743 (
            .O(N__34061),
            .I(N__33995));
    InMux I__7742 (
            .O(N__34060),
            .I(N__33991));
    InMux I__7741 (
            .O(N__34059),
            .I(N__33986));
    InMux I__7740 (
            .O(N__34058),
            .I(N__33986));
    InMux I__7739 (
            .O(N__34057),
            .I(N__33983));
    InMux I__7738 (
            .O(N__34056),
            .I(N__33974));
    InMux I__7737 (
            .O(N__34055),
            .I(N__33974));
    InMux I__7736 (
            .O(N__34054),
            .I(N__33974));
    InMux I__7735 (
            .O(N__34053),
            .I(N__33974));
    InMux I__7734 (
            .O(N__34052),
            .I(N__33967));
    InMux I__7733 (
            .O(N__34051),
            .I(N__33967));
    InMux I__7732 (
            .O(N__34050),
            .I(N__33967));
    LocalMux I__7731 (
            .O(N__34041),
            .I(N__33964));
    InMux I__7730 (
            .O(N__34038),
            .I(N__33957));
    InMux I__7729 (
            .O(N__34037),
            .I(N__33957));
    InMux I__7728 (
            .O(N__34036),
            .I(N__33957));
    Span4Mux_h I__7727 (
            .O(N__34033),
            .I(N__33952));
    LocalMux I__7726 (
            .O(N__34024),
            .I(N__33952));
    LocalMux I__7725 (
            .O(N__34017),
            .I(N__33949));
    LocalMux I__7724 (
            .O(N__34012),
            .I(N__33946));
    LocalMux I__7723 (
            .O(N__34007),
            .I(N__33943));
    InMux I__7722 (
            .O(N__34006),
            .I(N__33940));
    LocalMux I__7721 (
            .O(N__34003),
            .I(N__33933));
    LocalMux I__7720 (
            .O(N__33998),
            .I(N__33933));
    Span4Mux_h I__7719 (
            .O(N__33995),
            .I(N__33933));
    InMux I__7718 (
            .O(N__33994),
            .I(N__33930));
    LocalMux I__7717 (
            .O(N__33991),
            .I(N__33924));
    LocalMux I__7716 (
            .O(N__33986),
            .I(N__33924));
    LocalMux I__7715 (
            .O(N__33983),
            .I(N__33919));
    LocalMux I__7714 (
            .O(N__33974),
            .I(N__33919));
    LocalMux I__7713 (
            .O(N__33967),
            .I(N__33912));
    Span4Mux_h I__7712 (
            .O(N__33964),
            .I(N__33912));
    LocalMux I__7711 (
            .O(N__33957),
            .I(N__33912));
    Sp12to4 I__7710 (
            .O(N__33952),
            .I(N__33907));
    Span12Mux_s2_h I__7709 (
            .O(N__33949),
            .I(N__33907));
    Span4Mux_s0_h I__7708 (
            .O(N__33946),
            .I(N__33899));
    Span4Mux_v I__7707 (
            .O(N__33943),
            .I(N__33899));
    LocalMux I__7706 (
            .O(N__33940),
            .I(N__33896));
    Span4Mux_v I__7705 (
            .O(N__33933),
            .I(N__33891));
    LocalMux I__7704 (
            .O(N__33930),
            .I(N__33891));
    InMux I__7703 (
            .O(N__33929),
            .I(N__33888));
    Span12Mux_v I__7702 (
            .O(N__33924),
            .I(N__33885));
    Span12Mux_s8_v I__7701 (
            .O(N__33919),
            .I(N__33880));
    Sp12to4 I__7700 (
            .O(N__33912),
            .I(N__33880));
    Span12Mux_v I__7699 (
            .O(N__33907),
            .I(N__33877));
    InMux I__7698 (
            .O(N__33906),
            .I(N__33870));
    InMux I__7697 (
            .O(N__33905),
            .I(N__33870));
    InMux I__7696 (
            .O(N__33904),
            .I(N__33870));
    Span4Mux_h I__7695 (
            .O(N__33899),
            .I(N__33863));
    Span4Mux_h I__7694 (
            .O(N__33896),
            .I(N__33863));
    Span4Mux_h I__7693 (
            .O(N__33891),
            .I(N__33863));
    LocalMux I__7692 (
            .O(N__33888),
            .I(SYNTHESIZED_WIRE_47keep));
    Odrv12 I__7691 (
            .O(N__33885),
            .I(SYNTHESIZED_WIRE_47keep));
    Odrv12 I__7690 (
            .O(N__33880),
            .I(SYNTHESIZED_WIRE_47keep));
    Odrv12 I__7689 (
            .O(N__33877),
            .I(SYNTHESIZED_WIRE_47keep));
    LocalMux I__7688 (
            .O(N__33870),
            .I(SYNTHESIZED_WIRE_47keep));
    Odrv4 I__7687 (
            .O(N__33863),
            .I(SYNTHESIZED_WIRE_47keep));
    InMux I__7686 (
            .O(N__33850),
            .I(N__33844));
    InMux I__7685 (
            .O(N__33849),
            .I(N__33844));
    LocalMux I__7684 (
            .O(N__33844),
            .I(\b2v_inst200.curr_stateZ0Z_2 ));
    CascadeMux I__7683 (
            .O(N__33841),
            .I(\b2v_inst200.curr_stateZ0Z_2_cascade_ ));
    InMux I__7682 (
            .O(N__33838),
            .I(N__33835));
    LocalMux I__7681 (
            .O(N__33835),
            .I(\b2v_inst200.HDA_SDO_FPGA_0 ));
    InMux I__7680 (
            .O(N__33832),
            .I(N__33823));
    InMux I__7679 (
            .O(N__33831),
            .I(N__33823));
    InMux I__7678 (
            .O(N__33830),
            .I(N__33823));
    LocalMux I__7677 (
            .O(N__33823),
            .I(N__33818));
    InMux I__7676 (
            .O(N__33822),
            .I(N__33813));
    InMux I__7675 (
            .O(N__33821),
            .I(N__33813));
    Odrv4 I__7674 (
            .O(N__33818),
            .I(\b2v_inst200.curr_stateZ0Z_0 ));
    LocalMux I__7673 (
            .O(N__33813),
            .I(\b2v_inst200.curr_stateZ0Z_0 ));
    InMux I__7672 (
            .O(N__33808),
            .I(N__33797));
    InMux I__7671 (
            .O(N__33807),
            .I(N__33797));
    InMux I__7670 (
            .O(N__33806),
            .I(N__33794));
    InMux I__7669 (
            .O(N__33805),
            .I(N__33785));
    InMux I__7668 (
            .O(N__33804),
            .I(N__33785));
    InMux I__7667 (
            .O(N__33803),
            .I(N__33785));
    InMux I__7666 (
            .O(N__33802),
            .I(N__33785));
    LocalMux I__7665 (
            .O(N__33797),
            .I(\b2v_inst200.curr_stateZ0Z_1 ));
    LocalMux I__7664 (
            .O(N__33794),
            .I(\b2v_inst200.curr_stateZ0Z_1 ));
    LocalMux I__7663 (
            .O(N__33785),
            .I(\b2v_inst200.curr_stateZ0Z_1 ));
    InMux I__7662 (
            .O(N__33778),
            .I(N__33774));
    CascadeMux I__7661 (
            .O(N__33777),
            .I(N__33771));
    LocalMux I__7660 (
            .O(N__33774),
            .I(N__33764));
    InMux I__7659 (
            .O(N__33771),
            .I(N__33759));
    InMux I__7658 (
            .O(N__33770),
            .I(N__33759));
    InMux I__7657 (
            .O(N__33769),
            .I(N__33752));
    InMux I__7656 (
            .O(N__33768),
            .I(N__33752));
    InMux I__7655 (
            .O(N__33767),
            .I(N__33752));
    Span4Mux_h I__7654 (
            .O(N__33764),
            .I(N__33749));
    LocalMux I__7653 (
            .O(N__33759),
            .I(N__33746));
    LocalMux I__7652 (
            .O(N__33752),
            .I(N__33743));
    Span4Mux_h I__7651 (
            .O(N__33749),
            .I(N__33738));
    Span4Mux_s2_h I__7650 (
            .O(N__33746),
            .I(N__33738));
    Span4Mux_s2_h I__7649 (
            .O(N__33743),
            .I(N__33735));
    Odrv4 I__7648 (
            .O(N__33738),
            .I(N_219));
    Odrv4 I__7647 (
            .O(N__33735),
            .I(N_219));
    InMux I__7646 (
            .O(N__33730),
            .I(N__33727));
    LocalMux I__7645 (
            .O(N__33727),
            .I(\b2v_inst200.m6_i_0 ));
    InMux I__7644 (
            .O(N__33724),
            .I(N__33721));
    LocalMux I__7643 (
            .O(N__33721),
            .I(\b2v_inst200.curr_state_0_0 ));
    InMux I__7642 (
            .O(N__33718),
            .I(N__33709));
    InMux I__7641 (
            .O(N__33717),
            .I(N__33706));
    InMux I__7640 (
            .O(N__33716),
            .I(N__33703));
    InMux I__7639 (
            .O(N__33715),
            .I(N__33698));
    InMux I__7638 (
            .O(N__33714),
            .I(N__33698));
    InMux I__7637 (
            .O(N__33713),
            .I(N__33693));
    InMux I__7636 (
            .O(N__33712),
            .I(N__33693));
    LocalMux I__7635 (
            .O(N__33709),
            .I(N__33690));
    LocalMux I__7634 (
            .O(N__33706),
            .I(N__33675));
    LocalMux I__7633 (
            .O(N__33703),
            .I(N__33672));
    LocalMux I__7632 (
            .O(N__33698),
            .I(N__33669));
    LocalMux I__7631 (
            .O(N__33693),
            .I(N__33666));
    Glb2LocalMux I__7630 (
            .O(N__33690),
            .I(N__33631));
    CEMux I__7629 (
            .O(N__33689),
            .I(N__33631));
    CEMux I__7628 (
            .O(N__33688),
            .I(N__33631));
    CEMux I__7627 (
            .O(N__33687),
            .I(N__33631));
    CEMux I__7626 (
            .O(N__33686),
            .I(N__33631));
    CEMux I__7625 (
            .O(N__33685),
            .I(N__33631));
    CEMux I__7624 (
            .O(N__33684),
            .I(N__33631));
    CEMux I__7623 (
            .O(N__33683),
            .I(N__33631));
    CEMux I__7622 (
            .O(N__33682),
            .I(N__33631));
    CEMux I__7621 (
            .O(N__33681),
            .I(N__33631));
    CEMux I__7620 (
            .O(N__33680),
            .I(N__33631));
    CEMux I__7619 (
            .O(N__33679),
            .I(N__33631));
    CEMux I__7618 (
            .O(N__33678),
            .I(N__33631));
    Glb2LocalMux I__7617 (
            .O(N__33675),
            .I(N__33631));
    Glb2LocalMux I__7616 (
            .O(N__33672),
            .I(N__33631));
    Glb2LocalMux I__7615 (
            .O(N__33669),
            .I(N__33631));
    Glb2LocalMux I__7614 (
            .O(N__33666),
            .I(N__33631));
    GlobalMux I__7613 (
            .O(N__33631),
            .I(N__33628));
    gio2CtrlBuf I__7612 (
            .O(N__33628),
            .I(b2v_inst16_delayed_vddq_pwrgd_en_g));
    CascadeMux I__7611 (
            .O(N__33625),
            .I(\b2v_inst6.count_rst_0_cascade_ ));
    InMux I__7610 (
            .O(N__33622),
            .I(N__33619));
    LocalMux I__7609 (
            .O(N__33619),
            .I(GPIO_FPGA_PCH_1_c));
    InMux I__7608 (
            .O(N__33616),
            .I(N__33613));
    LocalMux I__7607 (
            .O(N__33613),
            .I(N__33610));
    Span4Mux_v I__7606 (
            .O(N__33610),
            .I(N__33605));
    InMux I__7605 (
            .O(N__33609),
            .I(N__33599));
    InMux I__7604 (
            .O(N__33608),
            .I(N__33599));
    Sp12to4 I__7603 (
            .O(N__33605),
            .I(N__33596));
    CascadeMux I__7602 (
            .O(N__33604),
            .I(N__33587));
    LocalMux I__7601 (
            .O(N__33599),
            .I(N__33582));
    Span12Mux_s11_h I__7600 (
            .O(N__33596),
            .I(N__33579));
    InMux I__7599 (
            .O(N__33595),
            .I(N__33570));
    InMux I__7598 (
            .O(N__33594),
            .I(N__33570));
    InMux I__7597 (
            .O(N__33593),
            .I(N__33570));
    InMux I__7596 (
            .O(N__33592),
            .I(N__33570));
    InMux I__7595 (
            .O(N__33591),
            .I(N__33561));
    InMux I__7594 (
            .O(N__33590),
            .I(N__33561));
    InMux I__7593 (
            .O(N__33587),
            .I(N__33561));
    InMux I__7592 (
            .O(N__33586),
            .I(N__33561));
    InMux I__7591 (
            .O(N__33585),
            .I(N__33558));
    Odrv4 I__7590 (
            .O(N__33582),
            .I(\b2v_inst200.count_RNI_0_0 ));
    Odrv12 I__7589 (
            .O(N__33579),
            .I(\b2v_inst200.count_RNI_0_0 ));
    LocalMux I__7588 (
            .O(N__33570),
            .I(\b2v_inst200.count_RNI_0_0 ));
    LocalMux I__7587 (
            .O(N__33561),
            .I(\b2v_inst200.count_RNI_0_0 ));
    LocalMux I__7586 (
            .O(N__33558),
            .I(\b2v_inst200.count_RNI_0_0 ));
    CascadeMux I__7585 (
            .O(N__33547),
            .I(N_405_cascade_));
    CascadeMux I__7584 (
            .O(N__33544),
            .I(\b2v_inst200.m6_i_0_cascade_ ));
    CascadeMux I__7583 (
            .O(N__33541),
            .I(\b2v_inst200.N_57_cascade_ ));
    CascadeMux I__7582 (
            .O(N__33538),
            .I(\b2v_inst200.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__7581 (
            .O(N__33535),
            .I(N_406_cascade_));
    InMux I__7580 (
            .O(N__33532),
            .I(N__33529));
    LocalMux I__7579 (
            .O(N__33529),
            .I(\b2v_inst200.N_55 ));
    CascadeMux I__7578 (
            .O(N__33526),
            .I(N__33523));
    InMux I__7577 (
            .O(N__33523),
            .I(N__33517));
    InMux I__7576 (
            .O(N__33522),
            .I(N__33517));
    LocalMux I__7575 (
            .O(N__33517),
            .I(N_406));
    InMux I__7574 (
            .O(N__33514),
            .I(N__33511));
    LocalMux I__7573 (
            .O(N__33511),
            .I(\b2v_inst200.curr_state_0_1 ));
    CascadeMux I__7572 (
            .O(N__33508),
            .I(\b2v_inst200.N_202_cascade_ ));
    IoInMux I__7571 (
            .O(N__33505),
            .I(N__33502));
    LocalMux I__7570 (
            .O(N__33502),
            .I(N__33499));
    IoSpan4Mux I__7569 (
            .O(N__33499),
            .I(N__33496));
    Span4Mux_s3_h I__7568 (
            .O(N__33496),
            .I(N__33493));
    Span4Mux_h I__7567 (
            .O(N__33493),
            .I(N__33490));
    Span4Mux_h I__7566 (
            .O(N__33490),
            .I(N__33487));
    Odrv4 I__7565 (
            .O(N__33487),
            .I(HDA_SDO_FPGA_c));
    InMux I__7564 (
            .O(N__33484),
            .I(N__33480));
    InMux I__7563 (
            .O(N__33483),
            .I(N__33477));
    LocalMux I__7562 (
            .O(N__33480),
            .I(\b2v_inst20.counterZ0Z_29 ));
    LocalMux I__7561 (
            .O(N__33477),
            .I(\b2v_inst20.counterZ0Z_29 ));
    InMux I__7560 (
            .O(N__33472),
            .I(N__33468));
    InMux I__7559 (
            .O(N__33471),
            .I(N__33465));
    LocalMux I__7558 (
            .O(N__33468),
            .I(\b2v_inst20.counterZ0Z_28 ));
    LocalMux I__7557 (
            .O(N__33465),
            .I(\b2v_inst20.counterZ0Z_28 ));
    CascadeMux I__7556 (
            .O(N__33460),
            .I(N__33456));
    InMux I__7555 (
            .O(N__33459),
            .I(N__33453));
    InMux I__7554 (
            .O(N__33456),
            .I(N__33450));
    LocalMux I__7553 (
            .O(N__33453),
            .I(\b2v_inst20.counterZ0Z_31 ));
    LocalMux I__7552 (
            .O(N__33450),
            .I(\b2v_inst20.counterZ0Z_31 ));
    InMux I__7551 (
            .O(N__33445),
            .I(N__33441));
    InMux I__7550 (
            .O(N__33444),
            .I(N__33438));
    LocalMux I__7549 (
            .O(N__33441),
            .I(\b2v_inst20.counterZ0Z_30 ));
    LocalMux I__7548 (
            .O(N__33438),
            .I(\b2v_inst20.counterZ0Z_30 ));
    InMux I__7547 (
            .O(N__33433),
            .I(N__33430));
    LocalMux I__7546 (
            .O(N__33430),
            .I(N__33427));
    Span4Mux_h I__7545 (
            .O(N__33427),
            .I(N__33424));
    Odrv4 I__7544 (
            .O(N__33424),
            .I(\b2v_inst20.un4_counter_7_and ));
    InMux I__7543 (
            .O(N__33421),
            .I(N__33417));
    InMux I__7542 (
            .O(N__33420),
            .I(N__33414));
    LocalMux I__7541 (
            .O(N__33417),
            .I(\b2v_inst20.counterZ0Z_11 ));
    LocalMux I__7540 (
            .O(N__33414),
            .I(\b2v_inst20.counterZ0Z_11 ));
    InMux I__7539 (
            .O(N__33409),
            .I(N__33405));
    InMux I__7538 (
            .O(N__33408),
            .I(N__33402));
    LocalMux I__7537 (
            .O(N__33405),
            .I(\b2v_inst20.counterZ0Z_8 ));
    LocalMux I__7536 (
            .O(N__33402),
            .I(\b2v_inst20.counterZ0Z_8 ));
    CascadeMux I__7535 (
            .O(N__33397),
            .I(N__33393));
    InMux I__7534 (
            .O(N__33396),
            .I(N__33390));
    InMux I__7533 (
            .O(N__33393),
            .I(N__33387));
    LocalMux I__7532 (
            .O(N__33390),
            .I(\b2v_inst20.counterZ0Z_10 ));
    LocalMux I__7531 (
            .O(N__33387),
            .I(\b2v_inst20.counterZ0Z_10 ));
    InMux I__7530 (
            .O(N__33382),
            .I(N__33378));
    InMux I__7529 (
            .O(N__33381),
            .I(N__33375));
    LocalMux I__7528 (
            .O(N__33378),
            .I(\b2v_inst20.counterZ0Z_9 ));
    LocalMux I__7527 (
            .O(N__33375),
            .I(\b2v_inst20.counterZ0Z_9 ));
    CascadeMux I__7526 (
            .O(N__33370),
            .I(N__33367));
    InMux I__7525 (
            .O(N__33367),
            .I(N__33364));
    LocalMux I__7524 (
            .O(N__33364),
            .I(N__33361));
    Span4Mux_v I__7523 (
            .O(N__33361),
            .I(N__33358));
    Odrv4 I__7522 (
            .O(N__33358),
            .I(\b2v_inst20.un4_counter_2_and ));
    InMux I__7521 (
            .O(N__33355),
            .I(N__33351));
    InMux I__7520 (
            .O(N__33354),
            .I(N__33348));
    LocalMux I__7519 (
            .O(N__33351),
            .I(\b2v_inst20.counterZ0Z_12 ));
    LocalMux I__7518 (
            .O(N__33348),
            .I(\b2v_inst20.counterZ0Z_12 ));
    InMux I__7517 (
            .O(N__33343),
            .I(N__33339));
    InMux I__7516 (
            .O(N__33342),
            .I(N__33336));
    LocalMux I__7515 (
            .O(N__33339),
            .I(\b2v_inst20.counterZ0Z_14 ));
    LocalMux I__7514 (
            .O(N__33336),
            .I(\b2v_inst20.counterZ0Z_14 ));
    CascadeMux I__7513 (
            .O(N__33331),
            .I(N__33327));
    InMux I__7512 (
            .O(N__33330),
            .I(N__33324));
    InMux I__7511 (
            .O(N__33327),
            .I(N__33321));
    LocalMux I__7510 (
            .O(N__33324),
            .I(\b2v_inst20.counterZ0Z_15 ));
    LocalMux I__7509 (
            .O(N__33321),
            .I(\b2v_inst20.counterZ0Z_15 ));
    InMux I__7508 (
            .O(N__33316),
            .I(N__33312));
    InMux I__7507 (
            .O(N__33315),
            .I(N__33309));
    LocalMux I__7506 (
            .O(N__33312),
            .I(\b2v_inst20.counterZ0Z_13 ));
    LocalMux I__7505 (
            .O(N__33309),
            .I(\b2v_inst20.counterZ0Z_13 ));
    InMux I__7504 (
            .O(N__33304),
            .I(N__33301));
    LocalMux I__7503 (
            .O(N__33301),
            .I(N__33298));
    Span4Mux_v I__7502 (
            .O(N__33298),
            .I(N__33295));
    Odrv4 I__7501 (
            .O(N__33295),
            .I(\b2v_inst20.un4_counter_3_and ));
    InMux I__7500 (
            .O(N__33292),
            .I(N__33288));
    InMux I__7499 (
            .O(N__33291),
            .I(N__33285));
    LocalMux I__7498 (
            .O(N__33288),
            .I(\b2v_inst20.counterZ0Z_19 ));
    LocalMux I__7497 (
            .O(N__33285),
            .I(\b2v_inst20.counterZ0Z_19 ));
    InMux I__7496 (
            .O(N__33280),
            .I(N__33276));
    InMux I__7495 (
            .O(N__33279),
            .I(N__33273));
    LocalMux I__7494 (
            .O(N__33276),
            .I(\b2v_inst20.counterZ0Z_16 ));
    LocalMux I__7493 (
            .O(N__33273),
            .I(\b2v_inst20.counterZ0Z_16 ));
    CascadeMux I__7492 (
            .O(N__33268),
            .I(N__33264));
    InMux I__7491 (
            .O(N__33267),
            .I(N__33261));
    InMux I__7490 (
            .O(N__33264),
            .I(N__33258));
    LocalMux I__7489 (
            .O(N__33261),
            .I(\b2v_inst20.counterZ0Z_17 ));
    LocalMux I__7488 (
            .O(N__33258),
            .I(\b2v_inst20.counterZ0Z_17 ));
    InMux I__7487 (
            .O(N__33253),
            .I(N__33249));
    InMux I__7486 (
            .O(N__33252),
            .I(N__33246));
    LocalMux I__7485 (
            .O(N__33249),
            .I(\b2v_inst20.counterZ0Z_18 ));
    LocalMux I__7484 (
            .O(N__33246),
            .I(\b2v_inst20.counterZ0Z_18 ));
    CascadeMux I__7483 (
            .O(N__33241),
            .I(N__33238));
    InMux I__7482 (
            .O(N__33238),
            .I(N__33235));
    LocalMux I__7481 (
            .O(N__33235),
            .I(N__33232));
    Span4Mux_h I__7480 (
            .O(N__33232),
            .I(N__33229));
    Odrv4 I__7479 (
            .O(N__33229),
            .I(\b2v_inst20.un4_counter_4_and ));
    InMux I__7478 (
            .O(N__33226),
            .I(N__33222));
    InMux I__7477 (
            .O(N__33225),
            .I(N__33219));
    LocalMux I__7476 (
            .O(N__33222),
            .I(\b2v_inst20.counterZ0Z_23 ));
    LocalMux I__7475 (
            .O(N__33219),
            .I(\b2v_inst20.counterZ0Z_23 ));
    InMux I__7474 (
            .O(N__33214),
            .I(N__33210));
    InMux I__7473 (
            .O(N__33213),
            .I(N__33207));
    LocalMux I__7472 (
            .O(N__33210),
            .I(\b2v_inst20.counterZ0Z_22 ));
    LocalMux I__7471 (
            .O(N__33207),
            .I(\b2v_inst20.counterZ0Z_22 ));
    CascadeMux I__7470 (
            .O(N__33202),
            .I(N__33198));
    InMux I__7469 (
            .O(N__33201),
            .I(N__33195));
    InMux I__7468 (
            .O(N__33198),
            .I(N__33192));
    LocalMux I__7467 (
            .O(N__33195),
            .I(\b2v_inst20.counterZ0Z_21 ));
    LocalMux I__7466 (
            .O(N__33192),
            .I(\b2v_inst20.counterZ0Z_21 ));
    InMux I__7465 (
            .O(N__33187),
            .I(N__33183));
    InMux I__7464 (
            .O(N__33186),
            .I(N__33180));
    LocalMux I__7463 (
            .O(N__33183),
            .I(\b2v_inst20.counterZ0Z_20 ));
    LocalMux I__7462 (
            .O(N__33180),
            .I(\b2v_inst20.counterZ0Z_20 ));
    CascadeMux I__7461 (
            .O(N__33175),
            .I(N__33172));
    InMux I__7460 (
            .O(N__33172),
            .I(N__33169));
    LocalMux I__7459 (
            .O(N__33169),
            .I(N__33166));
    Span4Mux_h I__7458 (
            .O(N__33166),
            .I(N__33163));
    Odrv4 I__7457 (
            .O(N__33163),
            .I(\b2v_inst20.un4_counter_5_and ));
    InMux I__7456 (
            .O(N__33160),
            .I(N__33156));
    InMux I__7455 (
            .O(N__33159),
            .I(N__33153));
    LocalMux I__7454 (
            .O(N__33156),
            .I(\b2v_inst20.counterZ0Z_24 ));
    LocalMux I__7453 (
            .O(N__33153),
            .I(\b2v_inst20.counterZ0Z_24 ));
    InMux I__7452 (
            .O(N__33148),
            .I(N__33144));
    InMux I__7451 (
            .O(N__33147),
            .I(N__33141));
    LocalMux I__7450 (
            .O(N__33144),
            .I(N__33138));
    LocalMux I__7449 (
            .O(N__33141),
            .I(\b2v_inst20.counterZ0Z_27 ));
    Odrv4 I__7448 (
            .O(N__33138),
            .I(\b2v_inst20.counterZ0Z_27 ));
    CascadeMux I__7447 (
            .O(N__33133),
            .I(N__33130));
    InMux I__7446 (
            .O(N__33130),
            .I(N__33126));
    InMux I__7445 (
            .O(N__33129),
            .I(N__33123));
    LocalMux I__7444 (
            .O(N__33126),
            .I(N__33120));
    LocalMux I__7443 (
            .O(N__33123),
            .I(\b2v_inst20.counterZ0Z_25 ));
    Odrv4 I__7442 (
            .O(N__33120),
            .I(\b2v_inst20.counterZ0Z_25 ));
    InMux I__7441 (
            .O(N__33115),
            .I(N__33111));
    InMux I__7440 (
            .O(N__33114),
            .I(N__33108));
    LocalMux I__7439 (
            .O(N__33111),
            .I(N__33105));
    LocalMux I__7438 (
            .O(N__33108),
            .I(\b2v_inst20.counterZ0Z_26 ));
    Odrv4 I__7437 (
            .O(N__33105),
            .I(\b2v_inst20.counterZ0Z_26 ));
    CascadeMux I__7436 (
            .O(N__33100),
            .I(N__33097));
    InMux I__7435 (
            .O(N__33097),
            .I(N__33094));
    LocalMux I__7434 (
            .O(N__33094),
            .I(N__33091));
    Span4Mux_h I__7433 (
            .O(N__33091),
            .I(N__33088));
    Odrv4 I__7432 (
            .O(N__33088),
            .I(\b2v_inst20.un4_counter_6_and ));
    CascadeMux I__7431 (
            .O(N__33085),
            .I(\b2v_inst200.curr_stateZ0Z_1_cascade_ ));
    InMux I__7430 (
            .O(N__33082),
            .I(N__33078));
    InMux I__7429 (
            .O(N__33081),
            .I(N__33075));
    LocalMux I__7428 (
            .O(N__33078),
            .I(N__33072));
    LocalMux I__7427 (
            .O(N__33075),
            .I(N__33069));
    Span4Mux_v I__7426 (
            .O(N__33072),
            .I(N__33066));
    Span4Mux_h I__7425 (
            .O(N__33069),
            .I(N__33063));
    Span4Mux_h I__7424 (
            .O(N__33066),
            .I(N__33060));
    Span4Mux_h I__7423 (
            .O(N__33063),
            .I(N__33057));
    Span4Mux_h I__7422 (
            .O(N__33060),
            .I(N__33054));
    Odrv4 I__7421 (
            .O(N__33057),
            .I(N_405));
    Odrv4 I__7420 (
            .O(N__33054),
            .I(N_405));
    CascadeMux I__7419 (
            .O(N__33049),
            .I(\b2v_inst5.count_rst_6_cascade_ ));
    InMux I__7418 (
            .O(N__33046),
            .I(N__33041));
    InMux I__7417 (
            .O(N__33045),
            .I(N__33038));
    InMux I__7416 (
            .O(N__33044),
            .I(N__33035));
    LocalMux I__7415 (
            .O(N__33041),
            .I(\b2v_inst5.countZ0Z_8 ));
    LocalMux I__7414 (
            .O(N__33038),
            .I(\b2v_inst5.countZ0Z_8 ));
    LocalMux I__7413 (
            .O(N__33035),
            .I(\b2v_inst5.countZ0Z_8 ));
    InMux I__7412 (
            .O(N__33028),
            .I(N__33022));
    InMux I__7411 (
            .O(N__33027),
            .I(N__33022));
    LocalMux I__7410 (
            .O(N__33022),
            .I(\b2v_inst5.un2_count_1_cry_7_THRU_CO ));
    CascadeMux I__7409 (
            .O(N__33019),
            .I(\b2v_inst5.countZ0Z_8_cascade_ ));
    InMux I__7408 (
            .O(N__33016),
            .I(N__33013));
    LocalMux I__7407 (
            .O(N__33013),
            .I(\b2v_inst5.count_0_8 ));
    InMux I__7406 (
            .O(N__33010),
            .I(N__33007));
    LocalMux I__7405 (
            .O(N__33007),
            .I(\b2v_inst5.count_rst_10 ));
    CascadeMux I__7404 (
            .O(N__33004),
            .I(\b2v_inst5.count_rst_10_cascade_ ));
    CascadeMux I__7403 (
            .O(N__33001),
            .I(N__32998));
    InMux I__7402 (
            .O(N__32998),
            .I(N__32994));
    InMux I__7401 (
            .O(N__32997),
            .I(N__32991));
    LocalMux I__7400 (
            .O(N__32994),
            .I(\b2v_inst5.un2_count_1_axb_4 ));
    LocalMux I__7399 (
            .O(N__32991),
            .I(\b2v_inst5.un2_count_1_axb_4 ));
    InMux I__7398 (
            .O(N__32986),
            .I(N__32980));
    InMux I__7397 (
            .O(N__32985),
            .I(N__32980));
    LocalMux I__7396 (
            .O(N__32980),
            .I(\b2v_inst5.un2_count_1_cry_3_THRU_CO ));
    CascadeMux I__7395 (
            .O(N__32977),
            .I(\b2v_inst5.un2_count_1_axb_4_cascade_ ));
    CascadeMux I__7394 (
            .O(N__32974),
            .I(N__32971));
    InMux I__7393 (
            .O(N__32971),
            .I(N__32967));
    InMux I__7392 (
            .O(N__32970),
            .I(N__32964));
    LocalMux I__7391 (
            .O(N__32967),
            .I(\b2v_inst5.count_0_4 ));
    LocalMux I__7390 (
            .O(N__32964),
            .I(\b2v_inst5.count_0_4 ));
    InMux I__7389 (
            .O(N__32959),
            .I(N__32956));
    LocalMux I__7388 (
            .O(N__32956),
            .I(N__32943));
    InMux I__7387 (
            .O(N__32955),
            .I(N__32932));
    InMux I__7386 (
            .O(N__32954),
            .I(N__32932));
    InMux I__7385 (
            .O(N__32953),
            .I(N__32932));
    InMux I__7384 (
            .O(N__32952),
            .I(N__32932));
    InMux I__7383 (
            .O(N__32951),
            .I(N__32932));
    InMux I__7382 (
            .O(N__32950),
            .I(N__32921));
    InMux I__7381 (
            .O(N__32949),
            .I(N__32921));
    InMux I__7380 (
            .O(N__32948),
            .I(N__32921));
    InMux I__7379 (
            .O(N__32947),
            .I(N__32921));
    InMux I__7378 (
            .O(N__32946),
            .I(N__32921));
    Span4Mux_v I__7377 (
            .O(N__32943),
            .I(N__32918));
    LocalMux I__7376 (
            .O(N__32932),
            .I(N__32915));
    LocalMux I__7375 (
            .O(N__32921),
            .I(\b2v_inst5.N_390 ));
    Odrv4 I__7374 (
            .O(N__32918),
            .I(\b2v_inst5.N_390 ));
    Odrv4 I__7373 (
            .O(N__32915),
            .I(\b2v_inst5.N_390 ));
    InMux I__7372 (
            .O(N__32908),
            .I(N__32905));
    LocalMux I__7371 (
            .O(N__32905),
            .I(N__32901));
    InMux I__7370 (
            .O(N__32904),
            .I(N__32898));
    Odrv4 I__7369 (
            .O(N__32901),
            .I(\b2v_inst5.un2_count_1_cry_12_THRU_CO ));
    LocalMux I__7368 (
            .O(N__32898),
            .I(\b2v_inst5.un2_count_1_cry_12_THRU_CO ));
    SRMux I__7367 (
            .O(N__32893),
            .I(N__32889));
    SRMux I__7366 (
            .O(N__32892),
            .I(N__32886));
    LocalMux I__7365 (
            .O(N__32889),
            .I(N__32877));
    LocalMux I__7364 (
            .O(N__32886),
            .I(N__32874));
    SRMux I__7363 (
            .O(N__32885),
            .I(N__32871));
    CascadeMux I__7362 (
            .O(N__32884),
            .I(N__32862));
    CascadeMux I__7361 (
            .O(N__32883),
            .I(N__32858));
    SRMux I__7360 (
            .O(N__32882),
            .I(N__32855));
    SRMux I__7359 (
            .O(N__32881),
            .I(N__32852));
    SRMux I__7358 (
            .O(N__32880),
            .I(N__32849));
    Span4Mux_h I__7357 (
            .O(N__32877),
            .I(N__32842));
    Span4Mux_v I__7356 (
            .O(N__32874),
            .I(N__32842));
    LocalMux I__7355 (
            .O(N__32871),
            .I(N__32842));
    CascadeMux I__7354 (
            .O(N__32870),
            .I(N__32836));
    CascadeMux I__7353 (
            .O(N__32869),
            .I(N__32829));
    CascadeMux I__7352 (
            .O(N__32868),
            .I(N__32825));
    SRMux I__7351 (
            .O(N__32867),
            .I(N__32822));
    InMux I__7350 (
            .O(N__32866),
            .I(N__32819));
    InMux I__7349 (
            .O(N__32865),
            .I(N__32810));
    InMux I__7348 (
            .O(N__32862),
            .I(N__32810));
    InMux I__7347 (
            .O(N__32861),
            .I(N__32810));
    InMux I__7346 (
            .O(N__32858),
            .I(N__32810));
    LocalMux I__7345 (
            .O(N__32855),
            .I(N__32799));
    LocalMux I__7344 (
            .O(N__32852),
            .I(N__32794));
    LocalMux I__7343 (
            .O(N__32849),
            .I(N__32794));
    Span4Mux_v I__7342 (
            .O(N__32842),
            .I(N__32791));
    InMux I__7341 (
            .O(N__32841),
            .I(N__32786));
    InMux I__7340 (
            .O(N__32840),
            .I(N__32786));
    InMux I__7339 (
            .O(N__32839),
            .I(N__32779));
    InMux I__7338 (
            .O(N__32836),
            .I(N__32779));
    InMux I__7337 (
            .O(N__32835),
            .I(N__32779));
    InMux I__7336 (
            .O(N__32834),
            .I(N__32772));
    InMux I__7335 (
            .O(N__32833),
            .I(N__32772));
    InMux I__7334 (
            .O(N__32832),
            .I(N__32772));
    InMux I__7333 (
            .O(N__32829),
            .I(N__32765));
    InMux I__7332 (
            .O(N__32828),
            .I(N__32765));
    InMux I__7331 (
            .O(N__32825),
            .I(N__32765));
    LocalMux I__7330 (
            .O(N__32822),
            .I(N__32762));
    LocalMux I__7329 (
            .O(N__32819),
            .I(N__32757));
    LocalMux I__7328 (
            .O(N__32810),
            .I(N__32757));
    InMux I__7327 (
            .O(N__32809),
            .I(N__32752));
    InMux I__7326 (
            .O(N__32808),
            .I(N__32752));
    InMux I__7325 (
            .O(N__32807),
            .I(N__32747));
    InMux I__7324 (
            .O(N__32806),
            .I(N__32747));
    InMux I__7323 (
            .O(N__32805),
            .I(N__32742));
    InMux I__7322 (
            .O(N__32804),
            .I(N__32742));
    InMux I__7321 (
            .O(N__32803),
            .I(N__32737));
    InMux I__7320 (
            .O(N__32802),
            .I(N__32737));
    Span4Mux_v I__7319 (
            .O(N__32799),
            .I(N__32730));
    Span4Mux_v I__7318 (
            .O(N__32794),
            .I(N__32730));
    Span4Mux_s0_h I__7317 (
            .O(N__32791),
            .I(N__32730));
    LocalMux I__7316 (
            .O(N__32786),
            .I(N__32725));
    LocalMux I__7315 (
            .O(N__32779),
            .I(N__32725));
    LocalMux I__7314 (
            .O(N__32772),
            .I(N__32720));
    LocalMux I__7313 (
            .O(N__32765),
            .I(N__32720));
    Span4Mux_v I__7312 (
            .O(N__32762),
            .I(N__32707));
    Span4Mux_s1_h I__7311 (
            .O(N__32757),
            .I(N__32707));
    LocalMux I__7310 (
            .O(N__32752),
            .I(N__32707));
    LocalMux I__7309 (
            .O(N__32747),
            .I(N__32707));
    LocalMux I__7308 (
            .O(N__32742),
            .I(N__32707));
    LocalMux I__7307 (
            .O(N__32737),
            .I(N__32707));
    Span4Mux_h I__7306 (
            .O(N__32730),
            .I(N__32704));
    Span4Mux_s3_h I__7305 (
            .O(N__32725),
            .I(N__32701));
    Span4Mux_s3_h I__7304 (
            .O(N__32720),
            .I(N__32698));
    Span4Mux_v I__7303 (
            .O(N__32707),
            .I(N__32695));
    Odrv4 I__7302 (
            .O(N__32704),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv4 I__7301 (
            .O(N__32701),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv4 I__7300 (
            .O(N__32698),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv4 I__7299 (
            .O(N__32695),
            .I(\b2v_inst5.count_0_sqmuxa ));
    CEMux I__7298 (
            .O(N__32686),
            .I(N__32683));
    LocalMux I__7297 (
            .O(N__32683),
            .I(N__32675));
    InMux I__7296 (
            .O(N__32682),
            .I(N__32668));
    InMux I__7295 (
            .O(N__32681),
            .I(N__32668));
    CEMux I__7294 (
            .O(N__32680),
            .I(N__32668));
    CEMux I__7293 (
            .O(N__32679),
            .I(N__32665));
    CascadeMux I__7292 (
            .O(N__32678),
            .I(N__32661));
    Span4Mux_s3_v I__7291 (
            .O(N__32675),
            .I(N__32652));
    LocalMux I__7290 (
            .O(N__32668),
            .I(N__32652));
    LocalMux I__7289 (
            .O(N__32665),
            .I(N__32652));
    CascadeMux I__7288 (
            .O(N__32664),
            .I(N__32638));
    InMux I__7287 (
            .O(N__32661),
            .I(N__32626));
    CEMux I__7286 (
            .O(N__32660),
            .I(N__32626));
    CEMux I__7285 (
            .O(N__32659),
            .I(N__32623));
    Span4Mux_v I__7284 (
            .O(N__32652),
            .I(N__32620));
    InMux I__7283 (
            .O(N__32651),
            .I(N__32615));
    InMux I__7282 (
            .O(N__32650),
            .I(N__32615));
    InMux I__7281 (
            .O(N__32649),
            .I(N__32608));
    InMux I__7280 (
            .O(N__32648),
            .I(N__32608));
    InMux I__7279 (
            .O(N__32647),
            .I(N__32608));
    CEMux I__7278 (
            .O(N__32646),
            .I(N__32599));
    InMux I__7277 (
            .O(N__32645),
            .I(N__32599));
    InMux I__7276 (
            .O(N__32644),
            .I(N__32599));
    InMux I__7275 (
            .O(N__32643),
            .I(N__32599));
    InMux I__7274 (
            .O(N__32642),
            .I(N__32596));
    InMux I__7273 (
            .O(N__32641),
            .I(N__32589));
    InMux I__7272 (
            .O(N__32638),
            .I(N__32589));
    InMux I__7271 (
            .O(N__32637),
            .I(N__32589));
    InMux I__7270 (
            .O(N__32636),
            .I(N__32584));
    CEMux I__7269 (
            .O(N__32635),
            .I(N__32584));
    InMux I__7268 (
            .O(N__32634),
            .I(N__32581));
    InMux I__7267 (
            .O(N__32633),
            .I(N__32574));
    InMux I__7266 (
            .O(N__32632),
            .I(N__32574));
    InMux I__7265 (
            .O(N__32631),
            .I(N__32574));
    LocalMux I__7264 (
            .O(N__32626),
            .I(N__32571));
    LocalMux I__7263 (
            .O(N__32623),
            .I(N__32556));
    Span4Mux_s0_h I__7262 (
            .O(N__32620),
            .I(N__32556));
    LocalMux I__7261 (
            .O(N__32615),
            .I(N__32556));
    LocalMux I__7260 (
            .O(N__32608),
            .I(N__32556));
    LocalMux I__7259 (
            .O(N__32599),
            .I(N__32556));
    LocalMux I__7258 (
            .O(N__32596),
            .I(N__32556));
    LocalMux I__7257 (
            .O(N__32589),
            .I(N__32556));
    LocalMux I__7256 (
            .O(N__32584),
            .I(N__32553));
    LocalMux I__7255 (
            .O(N__32581),
            .I(N__32548));
    LocalMux I__7254 (
            .O(N__32574),
            .I(N__32548));
    Span4Mux_s2_h I__7253 (
            .O(N__32571),
            .I(N__32543));
    Span4Mux_v I__7252 (
            .O(N__32556),
            .I(N__32540));
    Span4Mux_s2_h I__7251 (
            .O(N__32553),
            .I(N__32535));
    Span4Mux_s2_h I__7250 (
            .O(N__32548),
            .I(N__32535));
    InMux I__7249 (
            .O(N__32547),
            .I(N__32530));
    InMux I__7248 (
            .O(N__32546),
            .I(N__32530));
    Odrv4 I__7247 (
            .O(N__32543),
            .I(\b2v_inst5.count_enZ0 ));
    Odrv4 I__7246 (
            .O(N__32540),
            .I(\b2v_inst5.count_enZ0 ));
    Odrv4 I__7245 (
            .O(N__32535),
            .I(\b2v_inst5.count_enZ0 ));
    LocalMux I__7244 (
            .O(N__32530),
            .I(\b2v_inst5.count_enZ0 ));
    CascadeMux I__7243 (
            .O(N__32521),
            .I(\b2v_inst5.count_rst_1_cascade_ ));
    InMux I__7242 (
            .O(N__32518),
            .I(N__32515));
    LocalMux I__7241 (
            .O(N__32515),
            .I(N__32512));
    Odrv12 I__7240 (
            .O(N__32512),
            .I(\b2v_inst5.count_0_13 ));
    InMux I__7239 (
            .O(N__32509),
            .I(N__32506));
    LocalMux I__7238 (
            .O(N__32506),
            .I(N__32501));
    CascadeMux I__7237 (
            .O(N__32505),
            .I(N__32497));
    InMux I__7236 (
            .O(N__32504),
            .I(N__32494));
    Span4Mux_v I__7235 (
            .O(N__32501),
            .I(N__32491));
    InMux I__7234 (
            .O(N__32500),
            .I(N__32488));
    InMux I__7233 (
            .O(N__32497),
            .I(N__32485));
    LocalMux I__7232 (
            .O(N__32494),
            .I(N__32482));
    Odrv4 I__7231 (
            .O(N__32491),
            .I(\b2v_inst5.countZ0Z_13 ));
    LocalMux I__7230 (
            .O(N__32488),
            .I(\b2v_inst5.countZ0Z_13 ));
    LocalMux I__7229 (
            .O(N__32485),
            .I(\b2v_inst5.countZ0Z_13 ));
    Odrv12 I__7228 (
            .O(N__32482),
            .I(\b2v_inst5.countZ0Z_13 ));
    CascadeMux I__7227 (
            .O(N__32473),
            .I(N__32470));
    InMux I__7226 (
            .O(N__32470),
            .I(N__32466));
    InMux I__7225 (
            .O(N__32469),
            .I(N__32463));
    LocalMux I__7224 (
            .O(N__32466),
            .I(N__32460));
    LocalMux I__7223 (
            .O(N__32463),
            .I(\b2v_inst5.countZ0Z_3 ));
    Odrv4 I__7222 (
            .O(N__32460),
            .I(\b2v_inst5.countZ0Z_3 ));
    InMux I__7221 (
            .O(N__32455),
            .I(N__32452));
    LocalMux I__7220 (
            .O(N__32452),
            .I(N__32449));
    Odrv12 I__7219 (
            .O(N__32449),
            .I(\b2v_inst5.count_1_i_a2_6_0 ));
    CascadeMux I__7218 (
            .O(N__32446),
            .I(\b2v_inst5.count_1_i_a2_4_0_cascade_ ));
    InMux I__7217 (
            .O(N__32443),
            .I(N__32438));
    InMux I__7216 (
            .O(N__32442),
            .I(N__32433));
    InMux I__7215 (
            .O(N__32441),
            .I(N__32433));
    LocalMux I__7214 (
            .O(N__32438),
            .I(N__32430));
    LocalMux I__7213 (
            .O(N__32433),
            .I(\b2v_inst5.count_1_i_a2_12_0 ));
    Odrv4 I__7212 (
            .O(N__32430),
            .I(\b2v_inst5.count_1_i_a2_12_0 ));
    InMux I__7211 (
            .O(N__32425),
            .I(N__32419));
    InMux I__7210 (
            .O(N__32424),
            .I(N__32419));
    LocalMux I__7209 (
            .O(N__32419),
            .I(\b2v_inst5.count_0_2 ));
    InMux I__7208 (
            .O(N__32416),
            .I(N__32407));
    InMux I__7207 (
            .O(N__32415),
            .I(N__32407));
    InMux I__7206 (
            .O(N__32414),
            .I(N__32407));
    LocalMux I__7205 (
            .O(N__32407),
            .I(\b2v_inst5.count_rst_12 ));
    InMux I__7204 (
            .O(N__32404),
            .I(N__32401));
    LocalMux I__7203 (
            .O(N__32401),
            .I(\b2v_inst5.un2_count_1_axb_2 ));
    CascadeMux I__7202 (
            .O(N__32398),
            .I(N__32393));
    InMux I__7201 (
            .O(N__32397),
            .I(N__32390));
    InMux I__7200 (
            .O(N__32396),
            .I(N__32387));
    InMux I__7199 (
            .O(N__32393),
            .I(N__32384));
    LocalMux I__7198 (
            .O(N__32390),
            .I(\b2v_inst5.countZ0Z_1 ));
    LocalMux I__7197 (
            .O(N__32387),
            .I(\b2v_inst5.countZ0Z_1 ));
    LocalMux I__7196 (
            .O(N__32384),
            .I(\b2v_inst5.countZ0Z_1 ));
    InMux I__7195 (
            .O(N__32377),
            .I(N__32374));
    LocalMux I__7194 (
            .O(N__32374),
            .I(\b2v_inst5.count_1_i_a2_3_0 ));
    CascadeMux I__7193 (
            .O(N__32371),
            .I(N__32368));
    InMux I__7192 (
            .O(N__32368),
            .I(N__32362));
    InMux I__7191 (
            .O(N__32367),
            .I(N__32362));
    LocalMux I__7190 (
            .O(N__32362),
            .I(\b2v_inst5.count_0_11 ));
    InMux I__7189 (
            .O(N__32359),
            .I(N__32350));
    InMux I__7188 (
            .O(N__32358),
            .I(N__32350));
    InMux I__7187 (
            .O(N__32357),
            .I(N__32350));
    LocalMux I__7186 (
            .O(N__32350),
            .I(\b2v_inst5.count_rst_3 ));
    InMux I__7185 (
            .O(N__32347),
            .I(N__32344));
    LocalMux I__7184 (
            .O(N__32344),
            .I(\b2v_inst5.un2_count_1_axb_11 ));
    InMux I__7183 (
            .O(N__32341),
            .I(N__32338));
    LocalMux I__7182 (
            .O(N__32338),
            .I(\b2v_inst5.count_1_i_a2_5_0 ));
    CascadeMux I__7181 (
            .O(N__32335),
            .I(\b2v_inst5.count_RNIRHC7IZ0Z_2_cascade_ ));
    InMux I__7180 (
            .O(N__32332),
            .I(N__32328));
    InMux I__7179 (
            .O(N__32331),
            .I(N__32325));
    LocalMux I__7178 (
            .O(N__32328),
            .I(\b2v_inst5.countZ0Z_0 ));
    LocalMux I__7177 (
            .O(N__32325),
            .I(\b2v_inst5.countZ0Z_0 ));
    CascadeMux I__7176 (
            .O(N__32320),
            .I(\b2v_inst5.countZ0Z_0_cascade_ ));
    CascadeMux I__7175 (
            .O(N__32317),
            .I(\b2v_inst5.count_RNIZ0Z_0_cascade_ ));
    InMux I__7174 (
            .O(N__32314),
            .I(N__32311));
    LocalMux I__7173 (
            .O(N__32311),
            .I(\b2v_inst5.count_RNIZ0Z_0 ));
    InMux I__7172 (
            .O(N__32308),
            .I(N__32305));
    LocalMux I__7171 (
            .O(N__32305),
            .I(\b2v_inst5.count_0_1 ));
    InMux I__7170 (
            .O(N__32302),
            .I(N__32299));
    LocalMux I__7169 (
            .O(N__32299),
            .I(N__32294));
    InMux I__7168 (
            .O(N__32298),
            .I(N__32289));
    InMux I__7167 (
            .O(N__32297),
            .I(N__32289));
    Odrv4 I__7166 (
            .O(N__32294),
            .I(\b2v_inst5.count_1_i_a2_11_0 ));
    LocalMux I__7165 (
            .O(N__32289),
            .I(\b2v_inst5.count_1_i_a2_11_0 ));
    InMux I__7164 (
            .O(N__32284),
            .I(N__32278));
    InMux I__7163 (
            .O(N__32283),
            .I(N__32278));
    LocalMux I__7162 (
            .O(N__32278),
            .I(\b2v_inst5.N_2906_i ));
    InMux I__7161 (
            .O(N__32275),
            .I(N__32272));
    LocalMux I__7160 (
            .O(N__32272),
            .I(\b2v_inst5.count_0_0 ));
    CascadeMux I__7159 (
            .O(N__32269),
            .I(N__32266));
    InMux I__7158 (
            .O(N__32266),
            .I(N__32263));
    LocalMux I__7157 (
            .O(N__32263),
            .I(\b2v_inst5.count_0_3 ));
    InMux I__7156 (
            .O(N__32260),
            .I(N__32254));
    InMux I__7155 (
            .O(N__32259),
            .I(N__32254));
    LocalMux I__7154 (
            .O(N__32254),
            .I(\b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9 ));
    InMux I__7153 (
            .O(N__32251),
            .I(N__32248));
    LocalMux I__7152 (
            .O(N__32248),
            .I(\b2v_inst36.count_rst_14 ));
    InMux I__7151 (
            .O(N__32245),
            .I(N__32242));
    LocalMux I__7150 (
            .O(N__32242),
            .I(N__32238));
    InMux I__7149 (
            .O(N__32241),
            .I(N__32232));
    Span4Mux_s1_v I__7148 (
            .O(N__32238),
            .I(N__32229));
    InMux I__7147 (
            .O(N__32237),
            .I(N__32222));
    InMux I__7146 (
            .O(N__32236),
            .I(N__32222));
    InMux I__7145 (
            .O(N__32235),
            .I(N__32222));
    LocalMux I__7144 (
            .O(N__32232),
            .I(\b2v_inst36.countZ0Z_0 ));
    Odrv4 I__7143 (
            .O(N__32229),
            .I(\b2v_inst36.countZ0Z_0 ));
    LocalMux I__7142 (
            .O(N__32222),
            .I(\b2v_inst36.countZ0Z_0 ));
    InMux I__7141 (
            .O(N__32215),
            .I(N__32209));
    InMux I__7140 (
            .O(N__32214),
            .I(N__32209));
    LocalMux I__7139 (
            .O(N__32209),
            .I(N__32202));
    InMux I__7138 (
            .O(N__32208),
            .I(N__32190));
    InMux I__7137 (
            .O(N__32207),
            .I(N__32183));
    InMux I__7136 (
            .O(N__32206),
            .I(N__32183));
    InMux I__7135 (
            .O(N__32205),
            .I(N__32183));
    Span4Mux_s1_v I__7134 (
            .O(N__32202),
            .I(N__32174));
    InMux I__7133 (
            .O(N__32201),
            .I(N__32167));
    InMux I__7132 (
            .O(N__32200),
            .I(N__32167));
    InMux I__7131 (
            .O(N__32199),
            .I(N__32167));
    InMux I__7130 (
            .O(N__32198),
            .I(N__32160));
    InMux I__7129 (
            .O(N__32197),
            .I(N__32160));
    InMux I__7128 (
            .O(N__32196),
            .I(N__32160));
    InMux I__7127 (
            .O(N__32195),
            .I(N__32153));
    InMux I__7126 (
            .O(N__32194),
            .I(N__32153));
    InMux I__7125 (
            .O(N__32193),
            .I(N__32153));
    LocalMux I__7124 (
            .O(N__32190),
            .I(N__32148));
    LocalMux I__7123 (
            .O(N__32183),
            .I(N__32148));
    InMux I__7122 (
            .O(N__32182),
            .I(N__32140));
    InMux I__7121 (
            .O(N__32181),
            .I(N__32137));
    InMux I__7120 (
            .O(N__32180),
            .I(N__32128));
    InMux I__7119 (
            .O(N__32179),
            .I(N__32128));
    InMux I__7118 (
            .O(N__32178),
            .I(N__32128));
    InMux I__7117 (
            .O(N__32177),
            .I(N__32128));
    Span4Mux_h I__7116 (
            .O(N__32174),
            .I(N__32125));
    LocalMux I__7115 (
            .O(N__32167),
            .I(N__32116));
    LocalMux I__7114 (
            .O(N__32160),
            .I(N__32116));
    LocalMux I__7113 (
            .O(N__32153),
            .I(N__32116));
    Span12Mux_s1_v I__7112 (
            .O(N__32148),
            .I(N__32116));
    InMux I__7111 (
            .O(N__32147),
            .I(N__32105));
    InMux I__7110 (
            .O(N__32146),
            .I(N__32105));
    InMux I__7109 (
            .O(N__32145),
            .I(N__32105));
    InMux I__7108 (
            .O(N__32144),
            .I(N__32105));
    InMux I__7107 (
            .O(N__32143),
            .I(N__32105));
    LocalMux I__7106 (
            .O(N__32140),
            .I(\b2v_inst36.N_2928_i ));
    LocalMux I__7105 (
            .O(N__32137),
            .I(\b2v_inst36.N_2928_i ));
    LocalMux I__7104 (
            .O(N__32128),
            .I(\b2v_inst36.N_2928_i ));
    Odrv4 I__7103 (
            .O(N__32125),
            .I(\b2v_inst36.N_2928_i ));
    Odrv12 I__7102 (
            .O(N__32116),
            .I(\b2v_inst36.N_2928_i ));
    LocalMux I__7101 (
            .O(N__32105),
            .I(\b2v_inst36.N_2928_i ));
    CascadeMux I__7100 (
            .O(N__32092),
            .I(\b2v_inst36.countZ0Z_0_cascade_ ));
    CascadeMux I__7099 (
            .O(N__32089),
            .I(N__32077));
    InMux I__7098 (
            .O(N__32088),
            .I(N__32066));
    InMux I__7097 (
            .O(N__32087),
            .I(N__32066));
    InMux I__7096 (
            .O(N__32086),
            .I(N__32066));
    InMux I__7095 (
            .O(N__32085),
            .I(N__32066));
    InMux I__7094 (
            .O(N__32084),
            .I(N__32066));
    InMux I__7093 (
            .O(N__32083),
            .I(N__32057));
    InMux I__7092 (
            .O(N__32082),
            .I(N__32057));
    InMux I__7091 (
            .O(N__32081),
            .I(N__32057));
    InMux I__7090 (
            .O(N__32080),
            .I(N__32057));
    InMux I__7089 (
            .O(N__32077),
            .I(N__32048));
    LocalMux I__7088 (
            .O(N__32066),
            .I(N__32043));
    LocalMux I__7087 (
            .O(N__32057),
            .I(N__32043));
    CascadeMux I__7086 (
            .O(N__32056),
            .I(N__32039));
    CascadeMux I__7085 (
            .O(N__32055),
            .I(N__32035));
    InMux I__7084 (
            .O(N__32054),
            .I(N__32030));
    InMux I__7083 (
            .O(N__32053),
            .I(N__32027));
    InMux I__7082 (
            .O(N__32052),
            .I(N__32024));
    InMux I__7081 (
            .O(N__32051),
            .I(N__32021));
    LocalMux I__7080 (
            .O(N__32048),
            .I(N__32018));
    Span4Mux_s1_v I__7079 (
            .O(N__32043),
            .I(N__32015));
    InMux I__7078 (
            .O(N__32042),
            .I(N__32008));
    InMux I__7077 (
            .O(N__32039),
            .I(N__32008));
    InMux I__7076 (
            .O(N__32038),
            .I(N__32008));
    InMux I__7075 (
            .O(N__32035),
            .I(N__32001));
    InMux I__7074 (
            .O(N__32034),
            .I(N__32001));
    InMux I__7073 (
            .O(N__32033),
            .I(N__32001));
    LocalMux I__7072 (
            .O(N__32030),
            .I(\b2v_inst36.N_1_i ));
    LocalMux I__7071 (
            .O(N__32027),
            .I(\b2v_inst36.N_1_i ));
    LocalMux I__7070 (
            .O(N__32024),
            .I(\b2v_inst36.N_1_i ));
    LocalMux I__7069 (
            .O(N__32021),
            .I(\b2v_inst36.N_1_i ));
    Odrv12 I__7068 (
            .O(N__32018),
            .I(\b2v_inst36.N_1_i ));
    Odrv4 I__7067 (
            .O(N__32015),
            .I(\b2v_inst36.N_1_i ));
    LocalMux I__7066 (
            .O(N__32008),
            .I(\b2v_inst36.N_1_i ));
    LocalMux I__7065 (
            .O(N__32001),
            .I(\b2v_inst36.N_1_i ));
    InMux I__7064 (
            .O(N__31984),
            .I(N__31981));
    LocalMux I__7063 (
            .O(N__31981),
            .I(\b2v_inst36.count_1_0 ));
    CascadeMux I__7062 (
            .O(N__31978),
            .I(N__31971));
    CEMux I__7061 (
            .O(N__31977),
            .I(N__31967));
    CEMux I__7060 (
            .O(N__31976),
            .I(N__31955));
    CEMux I__7059 (
            .O(N__31975),
            .I(N__31946));
    InMux I__7058 (
            .O(N__31974),
            .I(N__31946));
    InMux I__7057 (
            .O(N__31971),
            .I(N__31946));
    InMux I__7056 (
            .O(N__31970),
            .I(N__31946));
    LocalMux I__7055 (
            .O(N__31967),
            .I(N__31943));
    InMux I__7054 (
            .O(N__31966),
            .I(N__31936));
    InMux I__7053 (
            .O(N__31965),
            .I(N__31936));
    InMux I__7052 (
            .O(N__31964),
            .I(N__31936));
    InMux I__7051 (
            .O(N__31963),
            .I(N__31929));
    CEMux I__7050 (
            .O(N__31962),
            .I(N__31926));
    InMux I__7049 (
            .O(N__31961),
            .I(N__31921));
    InMux I__7048 (
            .O(N__31960),
            .I(N__31921));
    InMux I__7047 (
            .O(N__31959),
            .I(N__31916));
    CEMux I__7046 (
            .O(N__31958),
            .I(N__31916));
    LocalMux I__7045 (
            .O(N__31955),
            .I(N__31912));
    LocalMux I__7044 (
            .O(N__31946),
            .I(N__31909));
    Span4Mux_s2_v I__7043 (
            .O(N__31943),
            .I(N__31904));
    LocalMux I__7042 (
            .O(N__31936),
            .I(N__31901));
    CEMux I__7041 (
            .O(N__31935),
            .I(N__31892));
    InMux I__7040 (
            .O(N__31934),
            .I(N__31892));
    InMux I__7039 (
            .O(N__31933),
            .I(N__31892));
    InMux I__7038 (
            .O(N__31932),
            .I(N__31892));
    LocalMux I__7037 (
            .O(N__31929),
            .I(N__31889));
    LocalMux I__7036 (
            .O(N__31926),
            .I(N__31884));
    LocalMux I__7035 (
            .O(N__31921),
            .I(N__31884));
    LocalMux I__7034 (
            .O(N__31916),
            .I(N__31881));
    InMux I__7033 (
            .O(N__31915),
            .I(N__31878));
    Span4Mux_s2_v I__7032 (
            .O(N__31912),
            .I(N__31873));
    Span4Mux_s2_v I__7031 (
            .O(N__31909),
            .I(N__31873));
    InMux I__7030 (
            .O(N__31908),
            .I(N__31868));
    InMux I__7029 (
            .O(N__31907),
            .I(N__31868));
    Span4Mux_s1_h I__7028 (
            .O(N__31904),
            .I(N__31863));
    Span4Mux_s2_v I__7027 (
            .O(N__31901),
            .I(N__31863));
    LocalMux I__7026 (
            .O(N__31892),
            .I(N__31860));
    Span4Mux_s3_h I__7025 (
            .O(N__31889),
            .I(N__31855));
    Span4Mux_s3_h I__7024 (
            .O(N__31884),
            .I(N__31855));
    Odrv4 I__7023 (
            .O(N__31881),
            .I(\b2v_inst36.count_en ));
    LocalMux I__7022 (
            .O(N__31878),
            .I(\b2v_inst36.count_en ));
    Odrv4 I__7021 (
            .O(N__31873),
            .I(\b2v_inst36.count_en ));
    LocalMux I__7020 (
            .O(N__31868),
            .I(\b2v_inst36.count_en ));
    Odrv4 I__7019 (
            .O(N__31863),
            .I(\b2v_inst36.count_en ));
    Odrv4 I__7018 (
            .O(N__31860),
            .I(\b2v_inst36.count_en ));
    Odrv4 I__7017 (
            .O(N__31855),
            .I(\b2v_inst36.count_en ));
    SRMux I__7016 (
            .O(N__31840),
            .I(N__31837));
    LocalMux I__7015 (
            .O(N__31837),
            .I(N__31832));
    SRMux I__7014 (
            .O(N__31836),
            .I(N__31829));
    SRMux I__7013 (
            .O(N__31835),
            .I(N__31824));
    Span4Mux_h I__7012 (
            .O(N__31832),
            .I(N__31819));
    LocalMux I__7011 (
            .O(N__31829),
            .I(N__31819));
    SRMux I__7010 (
            .O(N__31828),
            .I(N__31816));
    SRMux I__7009 (
            .O(N__31827),
            .I(N__31812));
    LocalMux I__7008 (
            .O(N__31824),
            .I(N__31809));
    Span4Mux_s1_h I__7007 (
            .O(N__31819),
            .I(N__31804));
    LocalMux I__7006 (
            .O(N__31816),
            .I(N__31804));
    SRMux I__7005 (
            .O(N__31815),
            .I(N__31801));
    LocalMux I__7004 (
            .O(N__31812),
            .I(N__31797));
    Span4Mux_h I__7003 (
            .O(N__31809),
            .I(N__31794));
    Span4Mux_s1_v I__7002 (
            .O(N__31804),
            .I(N__31789));
    LocalMux I__7001 (
            .O(N__31801),
            .I(N__31789));
    InMux I__7000 (
            .O(N__31800),
            .I(N__31786));
    Span4Mux_s2_v I__6999 (
            .O(N__31797),
            .I(N__31782));
    Span4Mux_s2_v I__6998 (
            .O(N__31794),
            .I(N__31779));
    Span4Mux_s1_h I__6997 (
            .O(N__31789),
            .I(N__31776));
    LocalMux I__6996 (
            .O(N__31786),
            .I(N__31773));
    InMux I__6995 (
            .O(N__31785),
            .I(N__31770));
    Odrv4 I__6994 (
            .O(N__31782),
            .I(\b2v_inst36.count_0_sqmuxa ));
    Odrv4 I__6993 (
            .O(N__31779),
            .I(\b2v_inst36.count_0_sqmuxa ));
    Odrv4 I__6992 (
            .O(N__31776),
            .I(\b2v_inst36.count_0_sqmuxa ));
    Odrv4 I__6991 (
            .O(N__31773),
            .I(\b2v_inst36.count_0_sqmuxa ));
    LocalMux I__6990 (
            .O(N__31770),
            .I(\b2v_inst36.count_0_sqmuxa ));
    InMux I__6989 (
            .O(N__31759),
            .I(N__31756));
    LocalMux I__6988 (
            .O(N__31756),
            .I(\b2v_inst5.count_rst_5 ));
    CascadeMux I__6987 (
            .O(N__31753),
            .I(\b2v_inst5.count_rst_5_cascade_ ));
    InMux I__6986 (
            .O(N__31750),
            .I(N__31747));
    LocalMux I__6985 (
            .O(N__31747),
            .I(N__31744));
    Span4Mux_v I__6984 (
            .O(N__31744),
            .I(N__31740));
    InMux I__6983 (
            .O(N__31743),
            .I(N__31737));
    Odrv4 I__6982 (
            .O(N__31740),
            .I(\b2v_inst5.un2_count_1_axb_9 ));
    LocalMux I__6981 (
            .O(N__31737),
            .I(\b2v_inst5.un2_count_1_axb_9 ));
    InMux I__6980 (
            .O(N__31732),
            .I(N__31726));
    InMux I__6979 (
            .O(N__31731),
            .I(N__31726));
    LocalMux I__6978 (
            .O(N__31726),
            .I(N__31723));
    Odrv4 I__6977 (
            .O(N__31723),
            .I(\b2v_inst5.un2_count_1_cry_8_THRU_CO ));
    CascadeMux I__6976 (
            .O(N__31720),
            .I(\b2v_inst5.un2_count_1_axb_9_cascade_ ));
    InMux I__6975 (
            .O(N__31717),
            .I(N__31711));
    InMux I__6974 (
            .O(N__31716),
            .I(N__31711));
    LocalMux I__6973 (
            .O(N__31711),
            .I(\b2v_inst5.count_0_9 ));
    CascadeMux I__6972 (
            .O(N__31708),
            .I(\b2v_inst5.count_rst_4_cascade_ ));
    InMux I__6971 (
            .O(N__31705),
            .I(N__31701));
    CascadeMux I__6970 (
            .O(N__31704),
            .I(N__31698));
    LocalMux I__6969 (
            .O(N__31701),
            .I(N__31694));
    InMux I__6968 (
            .O(N__31698),
            .I(N__31689));
    InMux I__6967 (
            .O(N__31697),
            .I(N__31689));
    Odrv4 I__6966 (
            .O(N__31694),
            .I(\b2v_inst5.countZ0Z_10 ));
    LocalMux I__6965 (
            .O(N__31689),
            .I(\b2v_inst5.countZ0Z_10 ));
    CascadeMux I__6964 (
            .O(N__31684),
            .I(\b2v_inst5.countZ0Z_10_cascade_ ));
    InMux I__6963 (
            .O(N__31681),
            .I(N__31675));
    InMux I__6962 (
            .O(N__31680),
            .I(N__31675));
    LocalMux I__6961 (
            .O(N__31675),
            .I(N__31672));
    Span4Mux_s0_h I__6960 (
            .O(N__31672),
            .I(N__31669));
    Odrv4 I__6959 (
            .O(N__31669),
            .I(\b2v_inst5.un2_count_1_cry_9_THRU_CO ));
    InMux I__6958 (
            .O(N__31666),
            .I(N__31663));
    LocalMux I__6957 (
            .O(N__31663),
            .I(\b2v_inst5.count_0_10 ));
    CascadeMux I__6956 (
            .O(N__31660),
            .I(\b2v_inst6.countZ0Z_8_cascade_ ));
    InMux I__6955 (
            .O(N__31657),
            .I(N__31651));
    InMux I__6954 (
            .O(N__31656),
            .I(N__31651));
    LocalMux I__6953 (
            .O(N__31651),
            .I(N__31648));
    Odrv12 I__6952 (
            .O(N__31648),
            .I(\b2v_inst6.un2_count_1_cry_7_THRU_CO ));
    InMux I__6951 (
            .O(N__31645),
            .I(N__31642));
    LocalMux I__6950 (
            .O(N__31642),
            .I(\b2v_inst6.count_3_8 ));
    CascadeMux I__6949 (
            .O(N__31639),
            .I(N__31636));
    InMux I__6948 (
            .O(N__31636),
            .I(N__31630));
    InMux I__6947 (
            .O(N__31635),
            .I(N__31625));
    InMux I__6946 (
            .O(N__31634),
            .I(N__31625));
    InMux I__6945 (
            .O(N__31633),
            .I(N__31622));
    LocalMux I__6944 (
            .O(N__31630),
            .I(\b2v_inst6.countZ0Z_9 ));
    LocalMux I__6943 (
            .O(N__31625),
            .I(\b2v_inst6.countZ0Z_9 ));
    LocalMux I__6942 (
            .O(N__31622),
            .I(\b2v_inst6.countZ0Z_9 ));
    InMux I__6941 (
            .O(N__31615),
            .I(N__31612));
    LocalMux I__6940 (
            .O(N__31612),
            .I(N__31608));
    InMux I__6939 (
            .O(N__31611),
            .I(N__31605));
    Odrv4 I__6938 (
            .O(N__31608),
            .I(\b2v_inst6.un2_count_1_cry_8_THRU_CO ));
    LocalMux I__6937 (
            .O(N__31605),
            .I(\b2v_inst6.un2_count_1_cry_8_THRU_CO ));
    InMux I__6936 (
            .O(N__31600),
            .I(N__31597));
    LocalMux I__6935 (
            .O(N__31597),
            .I(N__31594));
    Odrv4 I__6934 (
            .O(N__31594),
            .I(\b2v_inst6.count_3_9 ));
    CascadeMux I__6933 (
            .O(N__31591),
            .I(\b2v_inst36.N_2928_i_cascade_ ));
    InMux I__6932 (
            .O(N__31588),
            .I(N__31585));
    LocalMux I__6931 (
            .O(N__31585),
            .I(\b2v_inst36.count_1_13 ));
    InMux I__6930 (
            .O(N__31582),
            .I(N__31576));
    InMux I__6929 (
            .O(N__31581),
            .I(N__31576));
    LocalMux I__6928 (
            .O(N__31576),
            .I(N__31573));
    Odrv4 I__6927 (
            .O(N__31573),
            .I(\b2v_inst36.un2_count_1_cry_12_c_RNIS7LZ0Z1 ));
    CascadeMux I__6926 (
            .O(N__31570),
            .I(N__31566));
    InMux I__6925 (
            .O(N__31569),
            .I(N__31563));
    InMux I__6924 (
            .O(N__31566),
            .I(N__31560));
    LocalMux I__6923 (
            .O(N__31563),
            .I(N__31557));
    LocalMux I__6922 (
            .O(N__31560),
            .I(\b2v_inst36.countZ0Z_13 ));
    Odrv4 I__6921 (
            .O(N__31557),
            .I(\b2v_inst36.countZ0Z_13 ));
    CascadeMux I__6920 (
            .O(N__31552),
            .I(N__31549));
    InMux I__6919 (
            .O(N__31549),
            .I(N__31545));
    InMux I__6918 (
            .O(N__31548),
            .I(N__31542));
    LocalMux I__6917 (
            .O(N__31545),
            .I(N__31539));
    LocalMux I__6916 (
            .O(N__31542),
            .I(\b2v_inst36.countZ0Z_9 ));
    Odrv4 I__6915 (
            .O(N__31539),
            .I(\b2v_inst36.countZ0Z_9 ));
    CascadeMux I__6914 (
            .O(N__31534),
            .I(N__31531));
    InMux I__6913 (
            .O(N__31531),
            .I(N__31525));
    InMux I__6912 (
            .O(N__31530),
            .I(N__31525));
    LocalMux I__6911 (
            .O(N__31525),
            .I(N__31522));
    Span4Mux_s1_h I__6910 (
            .O(N__31522),
            .I(N__31519));
    Odrv4 I__6909 (
            .O(N__31519),
            .I(\b2v_inst36.un2_count_1_cry_8_c_RNIH8IZ0Z8 ));
    InMux I__6908 (
            .O(N__31516),
            .I(N__31513));
    LocalMux I__6907 (
            .O(N__31513),
            .I(\b2v_inst36.count_1_9 ));
    CascadeMux I__6906 (
            .O(N__31510),
            .I(\b2v_inst6.count_rst_8_cascade_ ));
    InMux I__6905 (
            .O(N__31507),
            .I(N__31501));
    InMux I__6904 (
            .O(N__31506),
            .I(N__31501));
    LocalMux I__6903 (
            .O(N__31501),
            .I(\b2v_inst6.count_rst_9 ));
    InMux I__6902 (
            .O(N__31498),
            .I(N__31495));
    LocalMux I__6901 (
            .O(N__31495),
            .I(N__31492));
    Odrv4 I__6900 (
            .O(N__31492),
            .I(\b2v_inst6.count_3_10 ));
    InMux I__6899 (
            .O(N__31489),
            .I(N__31485));
    CascadeMux I__6898 (
            .O(N__31488),
            .I(N__31481));
    LocalMux I__6897 (
            .O(N__31485),
            .I(N__31478));
    InMux I__6896 (
            .O(N__31484),
            .I(N__31475));
    InMux I__6895 (
            .O(N__31481),
            .I(N__31472));
    Span4Mux_s2_h I__6894 (
            .O(N__31478),
            .I(N__31469));
    LocalMux I__6893 (
            .O(N__31475),
            .I(N__31466));
    LocalMux I__6892 (
            .O(N__31472),
            .I(\b2v_inst6.countZ0Z_11 ));
    Odrv4 I__6891 (
            .O(N__31469),
            .I(\b2v_inst6.countZ0Z_11 ));
    Odrv12 I__6890 (
            .O(N__31466),
            .I(\b2v_inst6.countZ0Z_11 ));
    CascadeMux I__6889 (
            .O(N__31459),
            .I(\b2v_inst6.count_rst_6_cascade_ ));
    CascadeMux I__6888 (
            .O(N__31456),
            .I(N__31451));
    InMux I__6887 (
            .O(N__31455),
            .I(N__31448));
    InMux I__6886 (
            .O(N__31454),
            .I(N__31443));
    InMux I__6885 (
            .O(N__31451),
            .I(N__31443));
    LocalMux I__6884 (
            .O(N__31448),
            .I(N__31440));
    LocalMux I__6883 (
            .O(N__31443),
            .I(\b2v_inst6.countZ0Z_7 ));
    Odrv4 I__6882 (
            .O(N__31440),
            .I(\b2v_inst6.countZ0Z_7 ));
    InMux I__6881 (
            .O(N__31435),
            .I(N__31429));
    InMux I__6880 (
            .O(N__31434),
            .I(N__31429));
    LocalMux I__6879 (
            .O(N__31429),
            .I(N__31426));
    Odrv4 I__6878 (
            .O(N__31426),
            .I(\b2v_inst6.un2_count_1_cry_6_THRU_CO ));
    CascadeMux I__6877 (
            .O(N__31423),
            .I(\b2v_inst6.countZ0Z_7_cascade_ ));
    InMux I__6876 (
            .O(N__31420),
            .I(N__31417));
    LocalMux I__6875 (
            .O(N__31417),
            .I(\b2v_inst6.count_3_7 ));
    CascadeMux I__6874 (
            .O(N__31414),
            .I(\b2v_inst6.count_rst_7_cascade_ ));
    CascadeMux I__6873 (
            .O(N__31411),
            .I(N__31407));
    InMux I__6872 (
            .O(N__31410),
            .I(N__31403));
    InMux I__6871 (
            .O(N__31407),
            .I(N__31398));
    InMux I__6870 (
            .O(N__31406),
            .I(N__31398));
    LocalMux I__6869 (
            .O(N__31403),
            .I(N__31395));
    LocalMux I__6868 (
            .O(N__31398),
            .I(\b2v_inst6.countZ0Z_8 ));
    Odrv4 I__6867 (
            .O(N__31395),
            .I(\b2v_inst6.countZ0Z_8 ));
    InMux I__6866 (
            .O(N__31390),
            .I(\b2v_inst6.un2_count_1_cry_11 ));
    InMux I__6865 (
            .O(N__31387),
            .I(\b2v_inst6.un2_count_1_cry_12 ));
    InMux I__6864 (
            .O(N__31384),
            .I(\b2v_inst6.un2_count_1_cry_13 ));
    InMux I__6863 (
            .O(N__31381),
            .I(\b2v_inst6.un2_count_1_cry_14 ));
    CascadeMux I__6862 (
            .O(N__31378),
            .I(N__31375));
    InMux I__6861 (
            .O(N__31375),
            .I(N__31372));
    LocalMux I__6860 (
            .O(N__31372),
            .I(N__31368));
    InMux I__6859 (
            .O(N__31371),
            .I(N__31365));
    Span4Mux_s3_v I__6858 (
            .O(N__31368),
            .I(N__31362));
    LocalMux I__6857 (
            .O(N__31365),
            .I(N__31359));
    Odrv4 I__6856 (
            .O(N__31362),
            .I(\b2v_inst6.un2_count_1_cry_4_THRU_CO ));
    Odrv12 I__6855 (
            .O(N__31359),
            .I(\b2v_inst6.un2_count_1_cry_4_THRU_CO ));
    CascadeMux I__6854 (
            .O(N__31354),
            .I(\b2v_inst6.count_rst_4_cascade_ ));
    InMux I__6853 (
            .O(N__31351),
            .I(N__31348));
    LocalMux I__6852 (
            .O(N__31348),
            .I(N__31345));
    Span4Mux_s2_h I__6851 (
            .O(N__31345),
            .I(N__31342));
    Odrv4 I__6850 (
            .O(N__31342),
            .I(\b2v_inst6.count_3_5 ));
    CascadeMux I__6849 (
            .O(N__31339),
            .I(\b2v_inst6.count_rst_2_cascade_ ));
    InMux I__6848 (
            .O(N__31336),
            .I(\b2v_inst6.un2_count_1_cry_2 ));
    InMux I__6847 (
            .O(N__31333),
            .I(N__31327));
    InMux I__6846 (
            .O(N__31332),
            .I(N__31327));
    LocalMux I__6845 (
            .O(N__31327),
            .I(N__31324));
    Span4Mux_h I__6844 (
            .O(N__31324),
            .I(N__31321));
    Odrv4 I__6843 (
            .O(N__31321),
            .I(\b2v_inst6.un2_count_1_cry_3_THRU_CO ));
    InMux I__6842 (
            .O(N__31318),
            .I(\b2v_inst6.un2_count_1_cry_3 ));
    InMux I__6841 (
            .O(N__31315),
            .I(\b2v_inst6.un2_count_1_cry_4 ));
    InMux I__6840 (
            .O(N__31312),
            .I(\b2v_inst6.un2_count_1_cry_5 ));
    InMux I__6839 (
            .O(N__31309),
            .I(\b2v_inst6.un2_count_1_cry_6 ));
    InMux I__6838 (
            .O(N__31306),
            .I(\b2v_inst6.un2_count_1_cry_7 ));
    InMux I__6837 (
            .O(N__31303),
            .I(bfn_11_14_0_));
    InMux I__6836 (
            .O(N__31300),
            .I(\b2v_inst6.un2_count_1_cry_9 ));
    InMux I__6835 (
            .O(N__31297),
            .I(N__31291));
    InMux I__6834 (
            .O(N__31296),
            .I(N__31291));
    LocalMux I__6833 (
            .O(N__31291),
            .I(N__31288));
    Odrv4 I__6832 (
            .O(N__31288),
            .I(\b2v_inst6.un2_count_1_cry_10_THRU_CO ));
    InMux I__6831 (
            .O(N__31285),
            .I(\b2v_inst6.un2_count_1_cry_10 ));
    InMux I__6830 (
            .O(N__31282),
            .I(bfn_11_12_0_));
    InMux I__6829 (
            .O(N__31279),
            .I(\b2v_inst20.counter_1_cry_25 ));
    InMux I__6828 (
            .O(N__31276),
            .I(\b2v_inst20.counter_1_cry_26 ));
    InMux I__6827 (
            .O(N__31273),
            .I(\b2v_inst20.counter_1_cry_27 ));
    InMux I__6826 (
            .O(N__31270),
            .I(\b2v_inst20.counter_1_cry_28 ));
    InMux I__6825 (
            .O(N__31267),
            .I(\b2v_inst20.counter_1_cry_29 ));
    InMux I__6824 (
            .O(N__31264),
            .I(\b2v_inst20.counter_1_cry_30 ));
    InMux I__6823 (
            .O(N__31261),
            .I(\b2v_inst6.un2_count_1_cry_1 ));
    InMux I__6822 (
            .O(N__31258),
            .I(\b2v_inst20.counter_1_cry_15 ));
    InMux I__6821 (
            .O(N__31255),
            .I(bfn_11_11_0_));
    InMux I__6820 (
            .O(N__31252),
            .I(\b2v_inst20.counter_1_cry_17 ));
    InMux I__6819 (
            .O(N__31249),
            .I(\b2v_inst20.counter_1_cry_18 ));
    InMux I__6818 (
            .O(N__31246),
            .I(\b2v_inst20.counter_1_cry_19 ));
    InMux I__6817 (
            .O(N__31243),
            .I(\b2v_inst20.counter_1_cry_20 ));
    InMux I__6816 (
            .O(N__31240),
            .I(\b2v_inst20.counter_1_cry_21 ));
    InMux I__6815 (
            .O(N__31237),
            .I(\b2v_inst20.counter_1_cry_22 ));
    InMux I__6814 (
            .O(N__31234),
            .I(\b2v_inst20.counter_1_cry_23 ));
    InMux I__6813 (
            .O(N__31231),
            .I(N__31228));
    LocalMux I__6812 (
            .O(N__31228),
            .I(N__31224));
    InMux I__6811 (
            .O(N__31227),
            .I(N__31221));
    Span4Mux_h I__6810 (
            .O(N__31224),
            .I(N__31218));
    LocalMux I__6809 (
            .O(N__31221),
            .I(\b2v_inst20.counterZ0Z_7 ));
    Odrv4 I__6808 (
            .O(N__31218),
            .I(\b2v_inst20.counterZ0Z_7 ));
    InMux I__6807 (
            .O(N__31213),
            .I(\b2v_inst20.counter_1_cry_6 ));
    InMux I__6806 (
            .O(N__31210),
            .I(\b2v_inst20.counter_1_cry_7 ));
    InMux I__6805 (
            .O(N__31207),
            .I(bfn_11_10_0_));
    InMux I__6804 (
            .O(N__31204),
            .I(\b2v_inst20.counter_1_cry_9 ));
    InMux I__6803 (
            .O(N__31201),
            .I(\b2v_inst20.counter_1_cry_10 ));
    InMux I__6802 (
            .O(N__31198),
            .I(\b2v_inst20.counter_1_cry_11 ));
    InMux I__6801 (
            .O(N__31195),
            .I(\b2v_inst20.counter_1_cry_12 ));
    InMux I__6800 (
            .O(N__31192),
            .I(\b2v_inst20.counter_1_cry_13 ));
    InMux I__6799 (
            .O(N__31189),
            .I(\b2v_inst20.counter_1_cry_14 ));
    InMux I__6798 (
            .O(N__31186),
            .I(N__31183));
    LocalMux I__6797 (
            .O(N__31183),
            .I(N__31179));
    InMux I__6796 (
            .O(N__31182),
            .I(N__31176));
    Odrv4 I__6795 (
            .O(N__31179),
            .I(\b2v_inst5.countZ0Z_15 ));
    LocalMux I__6794 (
            .O(N__31176),
            .I(\b2v_inst5.countZ0Z_15 ));
    InMux I__6793 (
            .O(N__31171),
            .I(\b2v_inst5.un2_count_1_cry_14 ));
    InMux I__6792 (
            .O(N__31168),
            .I(N__31164));
    InMux I__6791 (
            .O(N__31167),
            .I(N__31161));
    LocalMux I__6790 (
            .O(N__31164),
            .I(N__31158));
    LocalMux I__6789 (
            .O(N__31161),
            .I(\b2v_inst5.count_rst ));
    Odrv12 I__6788 (
            .O(N__31158),
            .I(\b2v_inst5.count_rst ));
    InMux I__6787 (
            .O(N__31153),
            .I(N__31150));
    LocalMux I__6786 (
            .O(N__31150),
            .I(N__31147));
    Odrv12 I__6785 (
            .O(N__31147),
            .I(\b2v_inst5.count_0_15 ));
    InMux I__6784 (
            .O(N__31144),
            .I(N__31141));
    LocalMux I__6783 (
            .O(N__31141),
            .I(N__31137));
    InMux I__6782 (
            .O(N__31140),
            .I(N__31133));
    Span4Mux_s2_h I__6781 (
            .O(N__31137),
            .I(N__31130));
    InMux I__6780 (
            .O(N__31136),
            .I(N__31127));
    LocalMux I__6779 (
            .O(N__31133),
            .I(\b2v_inst20.counterZ0Z_1 ));
    Odrv4 I__6778 (
            .O(N__31130),
            .I(\b2v_inst20.counterZ0Z_1 ));
    LocalMux I__6777 (
            .O(N__31127),
            .I(\b2v_inst20.counterZ0Z_1 ));
    CascadeMux I__6776 (
            .O(N__31120),
            .I(N__31117));
    InMux I__6775 (
            .O(N__31117),
            .I(N__31114));
    LocalMux I__6774 (
            .O(N__31114),
            .I(N__31109));
    InMux I__6773 (
            .O(N__31113),
            .I(N__31105));
    InMux I__6772 (
            .O(N__31112),
            .I(N__31102));
    Span4Mux_s2_h I__6771 (
            .O(N__31109),
            .I(N__31099));
    InMux I__6770 (
            .O(N__31108),
            .I(N__31096));
    LocalMux I__6769 (
            .O(N__31105),
            .I(\b2v_inst20.counterZ0Z_0 ));
    LocalMux I__6768 (
            .O(N__31102),
            .I(\b2v_inst20.counterZ0Z_0 ));
    Odrv4 I__6767 (
            .O(N__31099),
            .I(\b2v_inst20.counterZ0Z_0 ));
    LocalMux I__6766 (
            .O(N__31096),
            .I(\b2v_inst20.counterZ0Z_0 ));
    InMux I__6765 (
            .O(N__31087),
            .I(N__31084));
    LocalMux I__6764 (
            .O(N__31084),
            .I(N__31080));
    InMux I__6763 (
            .O(N__31083),
            .I(N__31076));
    Span4Mux_s2_h I__6762 (
            .O(N__31080),
            .I(N__31073));
    InMux I__6761 (
            .O(N__31079),
            .I(N__31070));
    LocalMux I__6760 (
            .O(N__31076),
            .I(\b2v_inst20.counterZ0Z_2 ));
    Odrv4 I__6759 (
            .O(N__31073),
            .I(\b2v_inst20.counterZ0Z_2 ));
    LocalMux I__6758 (
            .O(N__31070),
            .I(\b2v_inst20.counterZ0Z_2 ));
    InMux I__6757 (
            .O(N__31063),
            .I(N__31060));
    LocalMux I__6756 (
            .O(N__31060),
            .I(N__31057));
    Span4Mux_h I__6755 (
            .O(N__31057),
            .I(N__31054));
    Odrv4 I__6754 (
            .O(N__31054),
            .I(\b2v_inst20.counter_1_cry_1_THRU_CO ));
    InMux I__6753 (
            .O(N__31051),
            .I(\b2v_inst20.counter_1_cry_1 ));
    InMux I__6752 (
            .O(N__31048),
            .I(N__31045));
    LocalMux I__6751 (
            .O(N__31045),
            .I(N__31040));
    CascadeMux I__6750 (
            .O(N__31044),
            .I(N__31037));
    InMux I__6749 (
            .O(N__31043),
            .I(N__31034));
    Span4Mux_s2_h I__6748 (
            .O(N__31040),
            .I(N__31031));
    InMux I__6747 (
            .O(N__31037),
            .I(N__31028));
    LocalMux I__6746 (
            .O(N__31034),
            .I(\b2v_inst20.counterZ0Z_3 ));
    Odrv4 I__6745 (
            .O(N__31031),
            .I(\b2v_inst20.counterZ0Z_3 ));
    LocalMux I__6744 (
            .O(N__31028),
            .I(\b2v_inst20.counterZ0Z_3 ));
    InMux I__6743 (
            .O(N__31021),
            .I(N__31018));
    LocalMux I__6742 (
            .O(N__31018),
            .I(N__31015));
    Span4Mux_h I__6741 (
            .O(N__31015),
            .I(N__31012));
    Odrv4 I__6740 (
            .O(N__31012),
            .I(\b2v_inst20.counter_1_cry_2_THRU_CO ));
    InMux I__6739 (
            .O(N__31009),
            .I(\b2v_inst20.counter_1_cry_2 ));
    InMux I__6738 (
            .O(N__31006),
            .I(N__31002));
    InMux I__6737 (
            .O(N__31005),
            .I(N__30998));
    LocalMux I__6736 (
            .O(N__31002),
            .I(N__30995));
    InMux I__6735 (
            .O(N__31001),
            .I(N__30992));
    LocalMux I__6734 (
            .O(N__30998),
            .I(\b2v_inst20.counterZ0Z_4 ));
    Odrv12 I__6733 (
            .O(N__30995),
            .I(\b2v_inst20.counterZ0Z_4 ));
    LocalMux I__6732 (
            .O(N__30992),
            .I(\b2v_inst20.counterZ0Z_4 ));
    InMux I__6731 (
            .O(N__30985),
            .I(N__30982));
    LocalMux I__6730 (
            .O(N__30982),
            .I(N__30979));
    Odrv12 I__6729 (
            .O(N__30979),
            .I(\b2v_inst20.counter_1_cry_3_THRU_CO ));
    InMux I__6728 (
            .O(N__30976),
            .I(\b2v_inst20.counter_1_cry_3 ));
    InMux I__6727 (
            .O(N__30973),
            .I(N__30970));
    LocalMux I__6726 (
            .O(N__30970),
            .I(N__30967));
    Span4Mux_s3_h I__6725 (
            .O(N__30967),
            .I(N__30962));
    InMux I__6724 (
            .O(N__30966),
            .I(N__30957));
    InMux I__6723 (
            .O(N__30965),
            .I(N__30957));
    Odrv4 I__6722 (
            .O(N__30962),
            .I(\b2v_inst20.counterZ0Z_5 ));
    LocalMux I__6721 (
            .O(N__30957),
            .I(\b2v_inst20.counterZ0Z_5 ));
    InMux I__6720 (
            .O(N__30952),
            .I(N__30949));
    LocalMux I__6719 (
            .O(N__30949),
            .I(N__30946));
    Span4Mux_v I__6718 (
            .O(N__30946),
            .I(N__30943));
    Odrv4 I__6717 (
            .O(N__30943),
            .I(\b2v_inst20.counter_1_cry_4_THRU_CO ));
    InMux I__6716 (
            .O(N__30940),
            .I(\b2v_inst20.counter_1_cry_4 ));
    InMux I__6715 (
            .O(N__30937),
            .I(N__30934));
    LocalMux I__6714 (
            .O(N__30934),
            .I(N__30930));
    CascadeMux I__6713 (
            .O(N__30933),
            .I(N__30926));
    Span4Mux_v I__6712 (
            .O(N__30930),
            .I(N__30923));
    InMux I__6711 (
            .O(N__30929),
            .I(N__30918));
    InMux I__6710 (
            .O(N__30926),
            .I(N__30918));
    Odrv4 I__6709 (
            .O(N__30923),
            .I(\b2v_inst20.counterZ0Z_6 ));
    LocalMux I__6708 (
            .O(N__30918),
            .I(\b2v_inst20.counterZ0Z_6 ));
    InMux I__6707 (
            .O(N__30913),
            .I(N__30910));
    LocalMux I__6706 (
            .O(N__30910),
            .I(N__30907));
    Span4Mux_v I__6705 (
            .O(N__30907),
            .I(N__30904));
    Span4Mux_h I__6704 (
            .O(N__30904),
            .I(N__30901));
    Odrv4 I__6703 (
            .O(N__30901),
            .I(\b2v_inst20.counter_1_cry_5_THRU_CO ));
    InMux I__6702 (
            .O(N__30898),
            .I(\b2v_inst20.counter_1_cry_5 ));
    CascadeMux I__6701 (
            .O(N__30895),
            .I(N__30892));
    InMux I__6700 (
            .O(N__30892),
            .I(N__30888));
    InMux I__6699 (
            .O(N__30891),
            .I(N__30885));
    LocalMux I__6698 (
            .O(N__30888),
            .I(N__30882));
    LocalMux I__6697 (
            .O(N__30885),
            .I(N__30879));
    Span4Mux_v I__6696 (
            .O(N__30882),
            .I(N__30876));
    Span4Mux_s2_h I__6695 (
            .O(N__30879),
            .I(N__30873));
    Odrv4 I__6694 (
            .O(N__30876),
            .I(\b2v_inst5.countZ0Z_7 ));
    Odrv4 I__6693 (
            .O(N__30873),
            .I(\b2v_inst5.countZ0Z_7 ));
    InMux I__6692 (
            .O(N__30868),
            .I(N__30864));
    InMux I__6691 (
            .O(N__30867),
            .I(N__30861));
    LocalMux I__6690 (
            .O(N__30864),
            .I(N__30858));
    LocalMux I__6689 (
            .O(N__30861),
            .I(N__30855));
    Span4Mux_h I__6688 (
            .O(N__30858),
            .I(N__30852));
    Odrv12 I__6687 (
            .O(N__30855),
            .I(\b2v_inst5.count_rst_7 ));
    Odrv4 I__6686 (
            .O(N__30852),
            .I(\b2v_inst5.count_rst_7 ));
    InMux I__6685 (
            .O(N__30847),
            .I(\b2v_inst5.un2_count_1_cry_6 ));
    InMux I__6684 (
            .O(N__30844),
            .I(\b2v_inst5.un2_count_1_cry_7 ));
    InMux I__6683 (
            .O(N__30841),
            .I(bfn_11_8_0_));
    InMux I__6682 (
            .O(N__30838),
            .I(\b2v_inst5.un2_count_1_cry_9 ));
    InMux I__6681 (
            .O(N__30835),
            .I(\b2v_inst5.un2_count_1_cry_10 ));
    CascadeMux I__6680 (
            .O(N__30832),
            .I(N__30829));
    InMux I__6679 (
            .O(N__30829),
            .I(N__30826));
    LocalMux I__6678 (
            .O(N__30826),
            .I(N__30823));
    Odrv4 I__6677 (
            .O(N__30823),
            .I(\b2v_inst5.un2_count_1_axb_12 ));
    InMux I__6676 (
            .O(N__30820),
            .I(N__30811));
    InMux I__6675 (
            .O(N__30819),
            .I(N__30811));
    InMux I__6674 (
            .O(N__30818),
            .I(N__30811));
    LocalMux I__6673 (
            .O(N__30811),
            .I(N__30808));
    Odrv4 I__6672 (
            .O(N__30808),
            .I(\b2v_inst5.count_rst_2 ));
    InMux I__6671 (
            .O(N__30805),
            .I(\b2v_inst5.un2_count_1_cry_11 ));
    InMux I__6670 (
            .O(N__30802),
            .I(\b2v_inst5.un2_count_1_cry_12 ));
    CascadeMux I__6669 (
            .O(N__30799),
            .I(N__30796));
    InMux I__6668 (
            .O(N__30796),
            .I(N__30793));
    LocalMux I__6667 (
            .O(N__30793),
            .I(N__30789));
    InMux I__6666 (
            .O(N__30792),
            .I(N__30786));
    Span4Mux_v I__6665 (
            .O(N__30789),
            .I(N__30783));
    LocalMux I__6664 (
            .O(N__30786),
            .I(N__30780));
    Odrv4 I__6663 (
            .O(N__30783),
            .I(\b2v_inst5.countZ0Z_14 ));
    Odrv12 I__6662 (
            .O(N__30780),
            .I(\b2v_inst5.countZ0Z_14 ));
    InMux I__6661 (
            .O(N__30775),
            .I(N__30771));
    InMux I__6660 (
            .O(N__30774),
            .I(N__30768));
    LocalMux I__6659 (
            .O(N__30771),
            .I(N__30765));
    LocalMux I__6658 (
            .O(N__30768),
            .I(N__30762));
    Odrv12 I__6657 (
            .O(N__30765),
            .I(\b2v_inst5.count_rst_0 ));
    Odrv4 I__6656 (
            .O(N__30762),
            .I(\b2v_inst5.count_rst_0 ));
    InMux I__6655 (
            .O(N__30757),
            .I(\b2v_inst5.un2_count_1_cry_13 ));
    InMux I__6654 (
            .O(N__30754),
            .I(N__30748));
    InMux I__6653 (
            .O(N__30753),
            .I(N__30748));
    LocalMux I__6652 (
            .O(N__30748),
            .I(\b2v_inst5.count_0_5 ));
    InMux I__6651 (
            .O(N__30745),
            .I(N__30741));
    InMux I__6650 (
            .O(N__30744),
            .I(N__30738));
    LocalMux I__6649 (
            .O(N__30741),
            .I(N__30735));
    LocalMux I__6648 (
            .O(N__30738),
            .I(N__30732));
    Span4Mux_v I__6647 (
            .O(N__30735),
            .I(N__30729));
    Odrv4 I__6646 (
            .O(N__30732),
            .I(\b2v_inst5.count_0_6 ));
    Odrv4 I__6645 (
            .O(N__30729),
            .I(\b2v_inst5.count_0_6 ));
    InMux I__6644 (
            .O(N__30724),
            .I(N__30721));
    LocalMux I__6643 (
            .O(N__30721),
            .I(\b2v_inst5.count_1_i_a2_2_0 ));
    InMux I__6642 (
            .O(N__30718),
            .I(\b2v_inst5.un2_count_1_cry_1 ));
    InMux I__6641 (
            .O(N__30715),
            .I(\b2v_inst5.un2_count_1_cry_2 ));
    InMux I__6640 (
            .O(N__30712),
            .I(\b2v_inst5.un2_count_1_cry_3 ));
    InMux I__6639 (
            .O(N__30709),
            .I(N__30706));
    LocalMux I__6638 (
            .O(N__30706),
            .I(\b2v_inst5.un2_count_1_axb_5 ));
    InMux I__6637 (
            .O(N__30703),
            .I(N__30694));
    InMux I__6636 (
            .O(N__30702),
            .I(N__30694));
    InMux I__6635 (
            .O(N__30701),
            .I(N__30694));
    LocalMux I__6634 (
            .O(N__30694),
            .I(\b2v_inst5.count_rst_9 ));
    InMux I__6633 (
            .O(N__30691),
            .I(\b2v_inst5.un2_count_1_cry_4 ));
    InMux I__6632 (
            .O(N__30688),
            .I(N__30685));
    LocalMux I__6631 (
            .O(N__30685),
            .I(N__30682));
    Span4Mux_s2_h I__6630 (
            .O(N__30682),
            .I(N__30679));
    Odrv4 I__6629 (
            .O(N__30679),
            .I(\b2v_inst5.un2_count_1_axb_6 ));
    InMux I__6628 (
            .O(N__30676),
            .I(N__30673));
    LocalMux I__6627 (
            .O(N__30673),
            .I(N__30670));
    Span4Mux_v I__6626 (
            .O(N__30670),
            .I(N__30666));
    InMux I__6625 (
            .O(N__30669),
            .I(N__30662));
    Sp12to4 I__6624 (
            .O(N__30666),
            .I(N__30659));
    InMux I__6623 (
            .O(N__30665),
            .I(N__30656));
    LocalMux I__6622 (
            .O(N__30662),
            .I(N__30653));
    Odrv12 I__6621 (
            .O(N__30659),
            .I(\b2v_inst5.count_rst_8 ));
    LocalMux I__6620 (
            .O(N__30656),
            .I(\b2v_inst5.count_rst_8 ));
    Odrv4 I__6619 (
            .O(N__30653),
            .I(\b2v_inst5.count_rst_8 ));
    InMux I__6618 (
            .O(N__30646),
            .I(\b2v_inst5.un2_count_1_cry_5 ));
    CascadeMux I__6617 (
            .O(N__30643),
            .I(N__30640));
    InMux I__6616 (
            .O(N__30640),
            .I(N__30634));
    CEMux I__6615 (
            .O(N__30639),
            .I(N__30634));
    LocalMux I__6614 (
            .O(N__30634),
            .I(N__30619));
    InMux I__6613 (
            .O(N__30633),
            .I(N__30610));
    InMux I__6612 (
            .O(N__30632),
            .I(N__30610));
    InMux I__6611 (
            .O(N__30631),
            .I(N__30610));
    InMux I__6610 (
            .O(N__30630),
            .I(N__30610));
    CEMux I__6609 (
            .O(N__30629),
            .I(N__30606));
    CEMux I__6608 (
            .O(N__30628),
            .I(N__30599));
    InMux I__6607 (
            .O(N__30627),
            .I(N__30589));
    InMux I__6606 (
            .O(N__30626),
            .I(N__30589));
    InMux I__6605 (
            .O(N__30625),
            .I(N__30589));
    InMux I__6604 (
            .O(N__30624),
            .I(N__30589));
    CEMux I__6603 (
            .O(N__30623),
            .I(N__30586));
    CEMux I__6602 (
            .O(N__30622),
            .I(N__30583));
    Span4Mux_s2_v I__6601 (
            .O(N__30619),
            .I(N__30578));
    LocalMux I__6600 (
            .O(N__30610),
            .I(N__30578));
    InMux I__6599 (
            .O(N__30609),
            .I(N__30575));
    LocalMux I__6598 (
            .O(N__30606),
            .I(N__30568));
    CEMux I__6597 (
            .O(N__30605),
            .I(N__30564));
    CEMux I__6596 (
            .O(N__30604),
            .I(N__30561));
    InMux I__6595 (
            .O(N__30603),
            .I(N__30556));
    InMux I__6594 (
            .O(N__30602),
            .I(N__30556));
    LocalMux I__6593 (
            .O(N__30599),
            .I(N__30553));
    CEMux I__6592 (
            .O(N__30598),
            .I(N__30550));
    LocalMux I__6591 (
            .O(N__30589),
            .I(N__30547));
    LocalMux I__6590 (
            .O(N__30586),
            .I(N__30538));
    LocalMux I__6589 (
            .O(N__30583),
            .I(N__30538));
    Span4Mux_v I__6588 (
            .O(N__30578),
            .I(N__30538));
    LocalMux I__6587 (
            .O(N__30575),
            .I(N__30538));
    InMux I__6586 (
            .O(N__30574),
            .I(N__30529));
    InMux I__6585 (
            .O(N__30573),
            .I(N__30529));
    InMux I__6584 (
            .O(N__30572),
            .I(N__30529));
    InMux I__6583 (
            .O(N__30571),
            .I(N__30529));
    Span4Mux_s2_h I__6582 (
            .O(N__30568),
            .I(N__30526));
    InMux I__6581 (
            .O(N__30567),
            .I(N__30523));
    LocalMux I__6580 (
            .O(N__30564),
            .I(N__30520));
    LocalMux I__6579 (
            .O(N__30561),
            .I(N__30515));
    LocalMux I__6578 (
            .O(N__30556),
            .I(N__30515));
    Span4Mux_s1_h I__6577 (
            .O(N__30553),
            .I(N__30512));
    LocalMux I__6576 (
            .O(N__30550),
            .I(N__30503));
    Span4Mux_s2_v I__6575 (
            .O(N__30547),
            .I(N__30503));
    Span4Mux_s2_v I__6574 (
            .O(N__30538),
            .I(N__30503));
    LocalMux I__6573 (
            .O(N__30529),
            .I(N__30503));
    Span4Mux_v I__6572 (
            .O(N__30526),
            .I(N__30498));
    LocalMux I__6571 (
            .O(N__30523),
            .I(N__30498));
    Span4Mux_h I__6570 (
            .O(N__30520),
            .I(N__30493));
    Span4Mux_s1_h I__6569 (
            .O(N__30515),
            .I(N__30493));
    Span4Mux_h I__6568 (
            .O(N__30512),
            .I(N__30490));
    Span4Mux_h I__6567 (
            .O(N__30503),
            .I(N__30487));
    Span4Mux_h I__6566 (
            .O(N__30498),
            .I(N__30482));
    Span4Mux_h I__6565 (
            .O(N__30493),
            .I(N__30482));
    Odrv4 I__6564 (
            .O(N__30490),
            .I(\b2v_inst16.count_en ));
    Odrv4 I__6563 (
            .O(N__30487),
            .I(\b2v_inst16.count_en ));
    Odrv4 I__6562 (
            .O(N__30482),
            .I(\b2v_inst16.count_en ));
    InMux I__6561 (
            .O(N__30475),
            .I(N__30472));
    LocalMux I__6560 (
            .O(N__30472),
            .I(N__30469));
    Span4Mux_v I__6559 (
            .O(N__30469),
            .I(N__30466));
    Odrv4 I__6558 (
            .O(N__30466),
            .I(\b2v_inst36.count_1_4 ));
    InMux I__6557 (
            .O(N__30463),
            .I(N__30459));
    InMux I__6556 (
            .O(N__30462),
            .I(N__30456));
    LocalMux I__6555 (
            .O(N__30459),
            .I(N__30453));
    LocalMux I__6554 (
            .O(N__30456),
            .I(N__30450));
    Span4Mux_v I__6553 (
            .O(N__30453),
            .I(N__30447));
    Odrv12 I__6552 (
            .O(N__30450),
            .I(\b2v_inst36.count_rst_10 ));
    Odrv4 I__6551 (
            .O(N__30447),
            .I(\b2v_inst36.count_rst_10 ));
    InMux I__6550 (
            .O(N__30442),
            .I(N__30438));
    InMux I__6549 (
            .O(N__30441),
            .I(N__30435));
    LocalMux I__6548 (
            .O(N__30438),
            .I(N__30432));
    LocalMux I__6547 (
            .O(N__30435),
            .I(N__30427));
    Span4Mux_h I__6546 (
            .O(N__30432),
            .I(N__30427));
    Odrv4 I__6545 (
            .O(N__30427),
            .I(\b2v_inst36.countZ0Z_4 ));
    CascadeMux I__6544 (
            .O(N__30424),
            .I(\b2v_inst5.N_2906_i_cascade_ ));
    CascadeMux I__6543 (
            .O(N__30421),
            .I(\b2v_inst5.count_1_i_a2_1_0_cascade_ ));
    InMux I__6542 (
            .O(N__30418),
            .I(N__30412));
    InMux I__6541 (
            .O(N__30417),
            .I(N__30412));
    LocalMux I__6540 (
            .O(N__30412),
            .I(\b2v_inst5.count_0_12 ));
    InMux I__6539 (
            .O(N__30409),
            .I(N__30406));
    LocalMux I__6538 (
            .O(N__30406),
            .I(\b2v_inst5.count_1_i_a2_0_0 ));
    InMux I__6537 (
            .O(N__30403),
            .I(N__30399));
    InMux I__6536 (
            .O(N__30402),
            .I(N__30396));
    LocalMux I__6535 (
            .O(N__30399),
            .I(N__30393));
    LocalMux I__6534 (
            .O(N__30396),
            .I(N__30390));
    Sp12to4 I__6533 (
            .O(N__30393),
            .I(N__30385));
    Span4Mux_v I__6532 (
            .O(N__30390),
            .I(N__30382));
    InMux I__6531 (
            .O(N__30389),
            .I(N__30379));
    InMux I__6530 (
            .O(N__30388),
            .I(N__30376));
    Span12Mux_v I__6529 (
            .O(N__30385),
            .I(N__30373));
    Odrv4 I__6528 (
            .O(N__30382),
            .I(\b2v_inst36.curr_stateZ0Z_0 ));
    LocalMux I__6527 (
            .O(N__30379),
            .I(\b2v_inst36.curr_stateZ0Z_0 ));
    LocalMux I__6526 (
            .O(N__30376),
            .I(\b2v_inst36.curr_stateZ0Z_0 ));
    Odrv12 I__6525 (
            .O(N__30373),
            .I(\b2v_inst36.curr_stateZ0Z_0 ));
    InMux I__6524 (
            .O(N__30364),
            .I(N__30361));
    LocalMux I__6523 (
            .O(N__30361),
            .I(\b2v_inst36.curr_state_4_0 ));
    InMux I__6522 (
            .O(N__30358),
            .I(N__30354));
    CascadeMux I__6521 (
            .O(N__30357),
            .I(N__30350));
    LocalMux I__6520 (
            .O(N__30354),
            .I(N__30346));
    CascadeMux I__6519 (
            .O(N__30353),
            .I(N__30343));
    InMux I__6518 (
            .O(N__30350),
            .I(N__30340));
    CascadeMux I__6517 (
            .O(N__30349),
            .I(N__30337));
    Span12Mux_v I__6516 (
            .O(N__30346),
            .I(N__30331));
    InMux I__6515 (
            .O(N__30343),
            .I(N__30328));
    LocalMux I__6514 (
            .O(N__30340),
            .I(N__30325));
    InMux I__6513 (
            .O(N__30337),
            .I(N__30316));
    InMux I__6512 (
            .O(N__30336),
            .I(N__30316));
    InMux I__6511 (
            .O(N__30335),
            .I(N__30316));
    InMux I__6510 (
            .O(N__30334),
            .I(N__30316));
    Odrv12 I__6509 (
            .O(N__30331),
            .I(\b2v_inst36.curr_stateZ0Z_1 ));
    LocalMux I__6508 (
            .O(N__30328),
            .I(\b2v_inst36.curr_stateZ0Z_1 ));
    Odrv4 I__6507 (
            .O(N__30325),
            .I(\b2v_inst36.curr_stateZ0Z_1 ));
    LocalMux I__6506 (
            .O(N__30316),
            .I(\b2v_inst36.curr_stateZ0Z_1 ));
    CascadeMux I__6505 (
            .O(N__30307),
            .I(N__30303));
    InMux I__6504 (
            .O(N__30306),
            .I(N__30295));
    InMux I__6503 (
            .O(N__30303),
            .I(N__30282));
    InMux I__6502 (
            .O(N__30302),
            .I(N__30282));
    InMux I__6501 (
            .O(N__30301),
            .I(N__30282));
    InMux I__6500 (
            .O(N__30300),
            .I(N__30282));
    InMux I__6499 (
            .O(N__30299),
            .I(N__30282));
    InMux I__6498 (
            .O(N__30298),
            .I(N__30282));
    LocalMux I__6497 (
            .O(N__30295),
            .I(N__30279));
    LocalMux I__6496 (
            .O(N__30282),
            .I(N__30276));
    Span4Mux_v I__6495 (
            .O(N__30279),
            .I(N__30273));
    Span4Mux_v I__6494 (
            .O(N__30276),
            .I(N__30270));
    Span4Mux_h I__6493 (
            .O(N__30273),
            .I(N__30265));
    Span4Mux_v I__6492 (
            .O(N__30270),
            .I(N__30265));
    Span4Mux_v I__6491 (
            .O(N__30265),
            .I(N__30262));
    Odrv4 I__6490 (
            .O(N__30262),
            .I(V33DSW_OK_c));
    InMux I__6489 (
            .O(N__30259),
            .I(N__30253));
    InMux I__6488 (
            .O(N__30258),
            .I(N__30246));
    InMux I__6487 (
            .O(N__30257),
            .I(N__30246));
    InMux I__6486 (
            .O(N__30256),
            .I(N__30246));
    LocalMux I__6485 (
            .O(N__30253),
            .I(N__30241));
    LocalMux I__6484 (
            .O(N__30246),
            .I(N__30241));
    Span4Mux_s3_h I__6483 (
            .O(N__30241),
            .I(N__30238));
    Span4Mux_v I__6482 (
            .O(N__30238),
            .I(N__30235));
    Span4Mux_h I__6481 (
            .O(N__30235),
            .I(N__30232));
    Odrv4 I__6480 (
            .O(N__30232),
            .I(\b2v_inst36.N_2925_i ));
    InMux I__6479 (
            .O(N__30229),
            .I(N__30226));
    LocalMux I__6478 (
            .O(N__30226),
            .I(N__30223));
    IoSpan4Mux I__6477 (
            .O(N__30223),
            .I(N__30220));
    IoSpan4Mux I__6476 (
            .O(N__30220),
            .I(N__30217));
    Odrv4 I__6475 (
            .O(N__30217),
            .I(\b2v_inst5.count_0_14 ));
    InMux I__6474 (
            .O(N__30214),
            .I(N__30211));
    LocalMux I__6473 (
            .O(N__30211),
            .I(N__30208));
    Span4Mux_v I__6472 (
            .O(N__30208),
            .I(N__30205));
    Span4Mux_h I__6471 (
            .O(N__30205),
            .I(N__30202));
    Odrv4 I__6470 (
            .O(N__30202),
            .I(\b2v_inst5.count_0_7 ));
    InMux I__6469 (
            .O(N__30199),
            .I(N__30195));
    InMux I__6468 (
            .O(N__30198),
            .I(N__30192));
    LocalMux I__6467 (
            .O(N__30195),
            .I(N__30187));
    LocalMux I__6466 (
            .O(N__30192),
            .I(N__30187));
    Span4Mux_s2_h I__6465 (
            .O(N__30187),
            .I(N__30184));
    Span4Mux_h I__6464 (
            .O(N__30184),
            .I(N__30181));
    Span4Mux_h I__6463 (
            .O(N__30181),
            .I(N__30178));
    Odrv4 I__6462 (
            .O(N__30178),
            .I(\b2v_inst16.countZ0Z_8 ));
    InMux I__6461 (
            .O(N__30175),
            .I(N__30169));
    InMux I__6460 (
            .O(N__30174),
            .I(N__30169));
    LocalMux I__6459 (
            .O(N__30169),
            .I(N__30166));
    Span4Mux_v I__6458 (
            .O(N__30166),
            .I(N__30163));
    Sp12to4 I__6457 (
            .O(N__30163),
            .I(N__30160));
    Odrv12 I__6456 (
            .O(N__30160),
            .I(\b2v_inst16.count_rst_13 ));
    InMux I__6455 (
            .O(N__30157),
            .I(N__30154));
    LocalMux I__6454 (
            .O(N__30154),
            .I(\b2v_inst16.count_4_8 ));
    InMux I__6453 (
            .O(N__30151),
            .I(N__30147));
    CascadeMux I__6452 (
            .O(N__30150),
            .I(N__30144));
    LocalMux I__6451 (
            .O(N__30147),
            .I(N__30141));
    InMux I__6450 (
            .O(N__30144),
            .I(N__30138));
    Span4Mux_s1_v I__6449 (
            .O(N__30141),
            .I(N__30135));
    LocalMux I__6448 (
            .O(N__30138),
            .I(N__30132));
    Span4Mux_h I__6447 (
            .O(N__30135),
            .I(N__30129));
    Span12Mux_s10_h I__6446 (
            .O(N__30132),
            .I(N__30126));
    Span4Mux_h I__6445 (
            .O(N__30129),
            .I(N__30123));
    Odrv12 I__6444 (
            .O(N__30126),
            .I(\b2v_inst16.countZ0Z_9 ));
    Odrv4 I__6443 (
            .O(N__30123),
            .I(\b2v_inst16.countZ0Z_9 ));
    InMux I__6442 (
            .O(N__30118),
            .I(N__30112));
    InMux I__6441 (
            .O(N__30117),
            .I(N__30112));
    LocalMux I__6440 (
            .O(N__30112),
            .I(N__30109));
    Span4Mux_s2_h I__6439 (
            .O(N__30109),
            .I(N__30106));
    Span4Mux_h I__6438 (
            .O(N__30106),
            .I(N__30103));
    Span4Mux_h I__6437 (
            .O(N__30103),
            .I(N__30100));
    Odrv4 I__6436 (
            .O(N__30100),
            .I(\b2v_inst16.count_rst_14 ));
    InMux I__6435 (
            .O(N__30097),
            .I(N__30094));
    LocalMux I__6434 (
            .O(N__30094),
            .I(\b2v_inst16.count_4_9 ));
    InMux I__6433 (
            .O(N__30091),
            .I(N__30088));
    LocalMux I__6432 (
            .O(N__30088),
            .I(N__30085));
    Span4Mux_s1_v I__6431 (
            .O(N__30085),
            .I(N__30081));
    InMux I__6430 (
            .O(N__30084),
            .I(N__30078));
    Odrv4 I__6429 (
            .O(N__30081),
            .I(\b2v_inst36.un2_count_1_cry_10_THRU_CO ));
    LocalMux I__6428 (
            .O(N__30078),
            .I(\b2v_inst36.un2_count_1_cry_10_THRU_CO ));
    CascadeMux I__6427 (
            .O(N__30073),
            .I(\b2v_inst36.countZ0Z_11_cascade_ ));
    InMux I__6426 (
            .O(N__30070),
            .I(N__30067));
    LocalMux I__6425 (
            .O(N__30067),
            .I(\b2v_inst36.count_1_11 ));
    CascadeMux I__6424 (
            .O(N__30064),
            .I(N__30061));
    InMux I__6423 (
            .O(N__30061),
            .I(N__30052));
    InMux I__6422 (
            .O(N__30060),
            .I(N__30052));
    InMux I__6421 (
            .O(N__30059),
            .I(N__30052));
    LocalMux I__6420 (
            .O(N__30052),
            .I(N__30049));
    Span4Mux_v I__6419 (
            .O(N__30049),
            .I(N__30046));
    Odrv4 I__6418 (
            .O(N__30046),
            .I(\b2v_inst36.count_rst_8 ));
    InMux I__6417 (
            .O(N__30043),
            .I(N__30037));
    InMux I__6416 (
            .O(N__30042),
            .I(N__30037));
    LocalMux I__6415 (
            .O(N__30037),
            .I(\b2v_inst36.count_1_6 ));
    InMux I__6414 (
            .O(N__30034),
            .I(N__30031));
    LocalMux I__6413 (
            .O(N__30031),
            .I(N__30028));
    Span4Mux_s2_v I__6412 (
            .O(N__30028),
            .I(N__30024));
    InMux I__6411 (
            .O(N__30027),
            .I(N__30021));
    Odrv4 I__6410 (
            .O(N__30024),
            .I(\b2v_inst36.countZ0Z_12 ));
    LocalMux I__6409 (
            .O(N__30021),
            .I(\b2v_inst36.countZ0Z_12 ));
    CascadeMux I__6408 (
            .O(N__30016),
            .I(\b2v_inst36.countZ0Z_6_cascade_ ));
    InMux I__6407 (
            .O(N__30013),
            .I(N__30010));
    LocalMux I__6406 (
            .O(N__30010),
            .I(\b2v_inst36.un12_clk_100khz_9 ));
    CascadeMux I__6405 (
            .O(N__30007),
            .I(\b2v_inst36.curr_stateZ0Z_1_cascade_ ));
    CascadeMux I__6404 (
            .O(N__30004),
            .I(\b2v_inst36.curr_state_7_0_cascade_ ));
    CascadeMux I__6403 (
            .O(N__30001),
            .I(\b2v_inst36.curr_stateZ0Z_0_cascade_ ));
    InMux I__6402 (
            .O(N__29998),
            .I(N__29995));
    LocalMux I__6401 (
            .O(N__29995),
            .I(N__29992));
    Span4Mux_h I__6400 (
            .O(N__29992),
            .I(N__29989));
    Span4Mux_v I__6399 (
            .O(N__29989),
            .I(N__29986));
    Odrv4 I__6398 (
            .O(N__29986),
            .I(\b2v_inst36.DSW_PWROK_0 ));
    InMux I__6397 (
            .O(N__29983),
            .I(N__29980));
    LocalMux I__6396 (
            .O(N__29980),
            .I(\b2v_inst36.curr_state_3_1 ));
    InMux I__6395 (
            .O(N__29977),
            .I(N__29974));
    LocalMux I__6394 (
            .O(N__29974),
            .I(\b2v_inst36.curr_state_7_1 ));
    CascadeMux I__6393 (
            .O(N__29971),
            .I(\b2v_inst36.count_rst_12_cascade_ ));
    InMux I__6392 (
            .O(N__29968),
            .I(N__29964));
    InMux I__6391 (
            .O(N__29967),
            .I(N__29960));
    LocalMux I__6390 (
            .O(N__29964),
            .I(N__29957));
    InMux I__6389 (
            .O(N__29963),
            .I(N__29954));
    LocalMux I__6388 (
            .O(N__29960),
            .I(N__29951));
    Odrv4 I__6387 (
            .O(N__29957),
            .I(\b2v_inst36.countZ0Z_2 ));
    LocalMux I__6386 (
            .O(N__29954),
            .I(\b2v_inst36.countZ0Z_2 ));
    Odrv4 I__6385 (
            .O(N__29951),
            .I(\b2v_inst36.countZ0Z_2 ));
    CascadeMux I__6384 (
            .O(N__29944),
            .I(\b2v_inst36.countZ0Z_2_cascade_ ));
    CascadeMux I__6383 (
            .O(N__29941),
            .I(N__29937));
    InMux I__6382 (
            .O(N__29940),
            .I(N__29934));
    InMux I__6381 (
            .O(N__29937),
            .I(N__29931));
    LocalMux I__6380 (
            .O(N__29934),
            .I(N__29926));
    LocalMux I__6379 (
            .O(N__29931),
            .I(N__29926));
    Span4Mux_s1_h I__6378 (
            .O(N__29926),
            .I(N__29923));
    Odrv4 I__6377 (
            .O(N__29923),
            .I(\b2v_inst36.un2_count_1_cry_1_THRU_CO ));
    InMux I__6376 (
            .O(N__29920),
            .I(N__29917));
    LocalMux I__6375 (
            .O(N__29917),
            .I(\b2v_inst36.count_1_2 ));
    CascadeMux I__6374 (
            .O(N__29914),
            .I(N__29910));
    InMux I__6373 (
            .O(N__29913),
            .I(N__29906));
    InMux I__6372 (
            .O(N__29910),
            .I(N__29900));
    InMux I__6371 (
            .O(N__29909),
            .I(N__29900));
    LocalMux I__6370 (
            .O(N__29906),
            .I(N__29897));
    InMux I__6369 (
            .O(N__29905),
            .I(N__29894));
    LocalMux I__6368 (
            .O(N__29900),
            .I(\b2v_inst36.countZ0Z_3 ));
    Odrv12 I__6367 (
            .O(N__29897),
            .I(\b2v_inst36.countZ0Z_3 ));
    LocalMux I__6366 (
            .O(N__29894),
            .I(\b2v_inst36.countZ0Z_3 ));
    InMux I__6365 (
            .O(N__29887),
            .I(N__29884));
    LocalMux I__6364 (
            .O(N__29884),
            .I(N__29880));
    InMux I__6363 (
            .O(N__29883),
            .I(N__29877));
    Odrv4 I__6362 (
            .O(N__29880),
            .I(\b2v_inst36.un2_count_1_cry_2_THRU_CO ));
    LocalMux I__6361 (
            .O(N__29877),
            .I(\b2v_inst36.un2_count_1_cry_2_THRU_CO ));
    InMux I__6360 (
            .O(N__29872),
            .I(N__29869));
    LocalMux I__6359 (
            .O(N__29869),
            .I(N__29866));
    Odrv12 I__6358 (
            .O(N__29866),
            .I(\b2v_inst36.count_1_3 ));
    InMux I__6357 (
            .O(N__29863),
            .I(N__29860));
    LocalMux I__6356 (
            .O(N__29860),
            .I(N__29855));
    InMux I__6355 (
            .O(N__29859),
            .I(N__29852));
    InMux I__6354 (
            .O(N__29858),
            .I(N__29849));
    Odrv12 I__6353 (
            .O(N__29855),
            .I(\b2v_inst36.countZ0Z_8 ));
    LocalMux I__6352 (
            .O(N__29852),
            .I(\b2v_inst36.countZ0Z_8 ));
    LocalMux I__6351 (
            .O(N__29849),
            .I(\b2v_inst36.countZ0Z_8 ));
    InMux I__6350 (
            .O(N__29842),
            .I(N__29838));
    CascadeMux I__6349 (
            .O(N__29841),
            .I(N__29835));
    LocalMux I__6348 (
            .O(N__29838),
            .I(N__29831));
    InMux I__6347 (
            .O(N__29835),
            .I(N__29828));
    InMux I__6346 (
            .O(N__29834),
            .I(N__29825));
    Odrv12 I__6345 (
            .O(N__29831),
            .I(\b2v_inst36.countZ0Z_10 ));
    LocalMux I__6344 (
            .O(N__29828),
            .I(\b2v_inst36.countZ0Z_10 ));
    LocalMux I__6343 (
            .O(N__29825),
            .I(\b2v_inst36.countZ0Z_10 ));
    CascadeMux I__6342 (
            .O(N__29818),
            .I(N__29814));
    CascadeMux I__6341 (
            .O(N__29817),
            .I(N__29811));
    InMux I__6340 (
            .O(N__29814),
            .I(N__29807));
    InMux I__6339 (
            .O(N__29811),
            .I(N__29804));
    InMux I__6338 (
            .O(N__29810),
            .I(N__29801));
    LocalMux I__6337 (
            .O(N__29807),
            .I(N__29798));
    LocalMux I__6336 (
            .O(N__29804),
            .I(\b2v_inst36.countZ0Z_1 ));
    LocalMux I__6335 (
            .O(N__29801),
            .I(\b2v_inst36.countZ0Z_1 ));
    Odrv4 I__6334 (
            .O(N__29798),
            .I(\b2v_inst36.countZ0Z_1 ));
    InMux I__6333 (
            .O(N__29791),
            .I(N__29788));
    LocalMux I__6332 (
            .O(N__29788),
            .I(N__29785));
    Span4Mux_v I__6331 (
            .O(N__29785),
            .I(N__29782));
    Odrv4 I__6330 (
            .O(N__29782),
            .I(\b2v_inst36.un12_clk_100khz_11 ));
    CascadeMux I__6329 (
            .O(N__29779),
            .I(\b2v_inst36.un12_clk_100khz_10_cascade_ ));
    InMux I__6328 (
            .O(N__29776),
            .I(N__29773));
    LocalMux I__6327 (
            .O(N__29773),
            .I(\b2v_inst36.un12_clk_100khz_8 ));
    InMux I__6326 (
            .O(N__29770),
            .I(N__29767));
    LocalMux I__6325 (
            .O(N__29767),
            .I(N__29764));
    Span4Mux_s1_v I__6324 (
            .O(N__29764),
            .I(N__29761));
    Odrv4 I__6323 (
            .O(N__29761),
            .I(\b2v_inst36.un2_count_1_axb_6 ));
    InMux I__6322 (
            .O(N__29758),
            .I(N__29755));
    LocalMux I__6321 (
            .O(N__29755),
            .I(N__29752));
    Odrv4 I__6320 (
            .O(N__29752),
            .I(\b2v_inst36.count_rst_3 ));
    CascadeMux I__6319 (
            .O(N__29749),
            .I(N__29746));
    InMux I__6318 (
            .O(N__29746),
            .I(N__29742));
    InMux I__6317 (
            .O(N__29745),
            .I(N__29738));
    LocalMux I__6316 (
            .O(N__29742),
            .I(N__29735));
    InMux I__6315 (
            .O(N__29741),
            .I(N__29732));
    LocalMux I__6314 (
            .O(N__29738),
            .I(N__29729));
    Odrv4 I__6313 (
            .O(N__29735),
            .I(\b2v_inst36.countZ0Z_11 ));
    LocalMux I__6312 (
            .O(N__29732),
            .I(\b2v_inst36.countZ0Z_11 ));
    Odrv4 I__6311 (
            .O(N__29729),
            .I(\b2v_inst36.countZ0Z_11 ));
    InMux I__6310 (
            .O(N__29722),
            .I(N__29718));
    InMux I__6309 (
            .O(N__29721),
            .I(N__29715));
    LocalMux I__6308 (
            .O(N__29718),
            .I(N__29710));
    LocalMux I__6307 (
            .O(N__29715),
            .I(N__29710));
    Odrv4 I__6306 (
            .O(N__29710),
            .I(VR_READY_VCCIN_c));
    CascadeMux I__6305 (
            .O(N__29707),
            .I(N__29703));
    InMux I__6304 (
            .O(N__29706),
            .I(N__29700));
    InMux I__6303 (
            .O(N__29703),
            .I(N__29697));
    LocalMux I__6302 (
            .O(N__29700),
            .I(N__29694));
    LocalMux I__6301 (
            .O(N__29697),
            .I(N__29691));
    Odrv4 I__6300 (
            .O(N__29694),
            .I(VR_READY_VCCINAUX_c));
    Odrv4 I__6299 (
            .O(N__29691),
            .I(VR_READY_VCCINAUX_c));
    IoInMux I__6298 (
            .O(N__29686),
            .I(N__29682));
    IoInMux I__6297 (
            .O(N__29685),
            .I(N__29679));
    LocalMux I__6296 (
            .O(N__29682),
            .I(N__29673));
    LocalMux I__6295 (
            .O(N__29679),
            .I(N__29673));
    CascadeMux I__6294 (
            .O(N__29678),
            .I(N__29667));
    IoSpan4Mux I__6293 (
            .O(N__29673),
            .I(N__29664));
    InMux I__6292 (
            .O(N__29672),
            .I(N__29661));
    CascadeMux I__6291 (
            .O(N__29671),
            .I(N__29655));
    CascadeMux I__6290 (
            .O(N__29670),
            .I(N__29649));
    InMux I__6289 (
            .O(N__29667),
            .I(N__29646));
    IoSpan4Mux I__6288 (
            .O(N__29664),
            .I(N__29643));
    LocalMux I__6287 (
            .O(N__29661),
            .I(N__29640));
    InMux I__6286 (
            .O(N__29660),
            .I(N__29635));
    InMux I__6285 (
            .O(N__29659),
            .I(N__29630));
    InMux I__6284 (
            .O(N__29658),
            .I(N__29627));
    InMux I__6283 (
            .O(N__29655),
            .I(N__29620));
    InMux I__6282 (
            .O(N__29654),
            .I(N__29620));
    InMux I__6281 (
            .O(N__29653),
            .I(N__29620));
    InMux I__6280 (
            .O(N__29652),
            .I(N__29616));
    InMux I__6279 (
            .O(N__29649),
            .I(N__29612));
    LocalMux I__6278 (
            .O(N__29646),
            .I(N__29609));
    Span4Mux_s2_h I__6277 (
            .O(N__29643),
            .I(N__29604));
    Span4Mux_v I__6276 (
            .O(N__29640),
            .I(N__29604));
    InMux I__6275 (
            .O(N__29639),
            .I(N__29601));
    InMux I__6274 (
            .O(N__29638),
            .I(N__29598));
    LocalMux I__6273 (
            .O(N__29635),
            .I(N__29595));
    InMux I__6272 (
            .O(N__29634),
            .I(N__29590));
    InMux I__6271 (
            .O(N__29633),
            .I(N__29590));
    LocalMux I__6270 (
            .O(N__29630),
            .I(N__29583));
    LocalMux I__6269 (
            .O(N__29627),
            .I(N__29583));
    LocalMux I__6268 (
            .O(N__29620),
            .I(N__29583));
    InMux I__6267 (
            .O(N__29619),
            .I(N__29580));
    LocalMux I__6266 (
            .O(N__29616),
            .I(N__29577));
    InMux I__6265 (
            .O(N__29615),
            .I(N__29574));
    LocalMux I__6264 (
            .O(N__29612),
            .I(N__29571));
    Span4Mux_v I__6263 (
            .O(N__29609),
            .I(N__29566));
    Span4Mux_h I__6262 (
            .O(N__29604),
            .I(N__29566));
    LocalMux I__6261 (
            .O(N__29601),
            .I(N__29553));
    LocalMux I__6260 (
            .O(N__29598),
            .I(N__29553));
    Span4Mux_h I__6259 (
            .O(N__29595),
            .I(N__29553));
    LocalMux I__6258 (
            .O(N__29590),
            .I(N__29553));
    Span4Mux_s3_v I__6257 (
            .O(N__29583),
            .I(N__29553));
    LocalMux I__6256 (
            .O(N__29580),
            .I(N__29553));
    Odrv12 I__6255 (
            .O(N__29577),
            .I(SYNTHESIZED_WIRE_48_i_0_o3_2));
    LocalMux I__6254 (
            .O(N__29574),
            .I(SYNTHESIZED_WIRE_48_i_0_o3_2));
    Odrv12 I__6253 (
            .O(N__29571),
            .I(SYNTHESIZED_WIRE_48_i_0_o3_2));
    Odrv4 I__6252 (
            .O(N__29566),
            .I(SYNTHESIZED_WIRE_48_i_0_o3_2));
    Odrv4 I__6251 (
            .O(N__29553),
            .I(SYNTHESIZED_WIRE_48_i_0_o3_2));
    CascadeMux I__6250 (
            .O(N__29542),
            .I(\b2v_inst6.N_413_cascade_ ));
    CascadeMux I__6249 (
            .O(N__29539),
            .I(\b2v_inst6.curr_state_7_1_cascade_ ));
    InMux I__6248 (
            .O(N__29536),
            .I(N__29529));
    InMux I__6247 (
            .O(N__29535),
            .I(N__29520));
    InMux I__6246 (
            .O(N__29534),
            .I(N__29520));
    InMux I__6245 (
            .O(N__29533),
            .I(N__29520));
    InMux I__6244 (
            .O(N__29532),
            .I(N__29520));
    LocalMux I__6243 (
            .O(N__29529),
            .I(\b2v_inst6.curr_stateZ0Z_1 ));
    LocalMux I__6242 (
            .O(N__29520),
            .I(\b2v_inst6.curr_stateZ0Z_1 ));
    CascadeMux I__6241 (
            .O(N__29515),
            .I(N__29507));
    InMux I__6240 (
            .O(N__29514),
            .I(N__29502));
    InMux I__6239 (
            .O(N__29513),
            .I(N__29493));
    InMux I__6238 (
            .O(N__29512),
            .I(N__29493));
    InMux I__6237 (
            .O(N__29511),
            .I(N__29493));
    InMux I__6236 (
            .O(N__29510),
            .I(N__29493));
    InMux I__6235 (
            .O(N__29507),
            .I(N__29486));
    InMux I__6234 (
            .O(N__29506),
            .I(N__29486));
    InMux I__6233 (
            .O(N__29505),
            .I(N__29486));
    LocalMux I__6232 (
            .O(N__29502),
            .I(\b2v_inst6.curr_stateZ0Z_0 ));
    LocalMux I__6231 (
            .O(N__29493),
            .I(\b2v_inst6.curr_stateZ0Z_0 ));
    LocalMux I__6230 (
            .O(N__29486),
            .I(\b2v_inst6.curr_stateZ0Z_0 ));
    CascadeMux I__6229 (
            .O(N__29479),
            .I(\b2v_inst6.curr_stateZ0Z_1_cascade_ ));
    InMux I__6228 (
            .O(N__29476),
            .I(N__29466));
    InMux I__6227 (
            .O(N__29475),
            .I(N__29466));
    InMux I__6226 (
            .O(N__29474),
            .I(N__29457));
    InMux I__6225 (
            .O(N__29473),
            .I(N__29457));
    InMux I__6224 (
            .O(N__29472),
            .I(N__29457));
    InMux I__6223 (
            .O(N__29471),
            .I(N__29457));
    LocalMux I__6222 (
            .O(N__29466),
            .I(\b2v_inst6.N_413 ));
    LocalMux I__6221 (
            .O(N__29457),
            .I(\b2v_inst6.N_413 ));
    InMux I__6220 (
            .O(N__29452),
            .I(N__29449));
    LocalMux I__6219 (
            .O(N__29449),
            .I(\b2v_inst6.curr_state_1_1 ));
    CascadeMux I__6218 (
            .O(N__29446),
            .I(\b2v_inst36.countZ0Z_1_cascade_ ));
    InMux I__6217 (
            .O(N__29443),
            .I(N__29440));
    LocalMux I__6216 (
            .O(N__29440),
            .I(\b2v_inst36.count_rst_13 ));
    InMux I__6215 (
            .O(N__29437),
            .I(N__29434));
    LocalMux I__6214 (
            .O(N__29434),
            .I(N__29431));
    Span4Mux_s1_v I__6213 (
            .O(N__29431),
            .I(N__29427));
    InMux I__6212 (
            .O(N__29430),
            .I(N__29424));
    Odrv4 I__6211 (
            .O(N__29427),
            .I(\b2v_inst36.countZ0Z_14 ));
    LocalMux I__6210 (
            .O(N__29424),
            .I(\b2v_inst36.countZ0Z_14 ));
    InMux I__6209 (
            .O(N__29419),
            .I(N__29416));
    LocalMux I__6208 (
            .O(N__29416),
            .I(N__29412));
    InMux I__6207 (
            .O(N__29415),
            .I(N__29409));
    Span4Mux_s3_h I__6206 (
            .O(N__29412),
            .I(N__29404));
    LocalMux I__6205 (
            .O(N__29409),
            .I(N__29404));
    Odrv4 I__6204 (
            .O(N__29404),
            .I(\b2v_inst36.countZ0Z_15 ));
    InMux I__6203 (
            .O(N__29401),
            .I(N__29398));
    LocalMux I__6202 (
            .O(N__29398),
            .I(\b2v_inst36.count_1_1 ));
    InMux I__6201 (
            .O(N__29395),
            .I(N__29392));
    LocalMux I__6200 (
            .O(N__29392),
            .I(\b2v_inst6.count_rst_10 ));
    CascadeMux I__6199 (
            .O(N__29389),
            .I(\b2v_inst6.count_rst_3_cascade_ ));
    CascadeMux I__6198 (
            .O(N__29386),
            .I(\b2v_inst6.countZ0Z_4_cascade_ ));
    InMux I__6197 (
            .O(N__29383),
            .I(N__29380));
    LocalMux I__6196 (
            .O(N__29380),
            .I(\b2v_inst6.count_3_4 ));
    CascadeMux I__6195 (
            .O(N__29377),
            .I(G_2746_cascade_));
    CascadeMux I__6194 (
            .O(N__29374),
            .I(\b2v_inst6.curr_stateZ0Z_0_cascade_ ));
    InMux I__6193 (
            .O(N__29371),
            .I(N__29368));
    LocalMux I__6192 (
            .O(N__29368),
            .I(\b2v_inst6.curr_state_2_0 ));
    InMux I__6191 (
            .O(N__29365),
            .I(N__29355));
    InMux I__6190 (
            .O(N__29364),
            .I(N__29355));
    InMux I__6189 (
            .O(N__29363),
            .I(N__29355));
    CascadeMux I__6188 (
            .O(N__29362),
            .I(N__29350));
    LocalMux I__6187 (
            .O(N__29355),
            .I(N__29347));
    InMux I__6186 (
            .O(N__29354),
            .I(N__29344));
    CascadeMux I__6185 (
            .O(N__29353),
            .I(N__29341));
    InMux I__6184 (
            .O(N__29350),
            .I(N__29338));
    Span4Mux_v I__6183 (
            .O(N__29347),
            .I(N__29335));
    LocalMux I__6182 (
            .O(N__29344),
            .I(N__29332));
    InMux I__6181 (
            .O(N__29341),
            .I(N__29329));
    LocalMux I__6180 (
            .O(N__29338),
            .I(N__29325));
    Span4Mux_h I__6179 (
            .O(N__29335),
            .I(N__29318));
    Span4Mux_v I__6178 (
            .O(N__29332),
            .I(N__29318));
    LocalMux I__6177 (
            .O(N__29329),
            .I(N__29318));
    InMux I__6176 (
            .O(N__29328),
            .I(N__29315));
    Span4Mux_v I__6175 (
            .O(N__29325),
            .I(N__29311));
    Span4Mux_h I__6174 (
            .O(N__29318),
            .I(N__29308));
    LocalMux I__6173 (
            .O(N__29315),
            .I(N__29305));
    InMux I__6172 (
            .O(N__29314),
            .I(N__29302));
    Odrv4 I__6171 (
            .O(N__29311),
            .I(\b2v_inst11.N_158 ));
    Odrv4 I__6170 (
            .O(N__29308),
            .I(\b2v_inst11.N_158 ));
    Odrv12 I__6169 (
            .O(N__29305),
            .I(\b2v_inst11.N_158 ));
    LocalMux I__6168 (
            .O(N__29302),
            .I(\b2v_inst11.N_158 ));
    CascadeMux I__6167 (
            .O(N__29293),
            .I(N__29290));
    InMux I__6166 (
            .O(N__29290),
            .I(N__29287));
    LocalMux I__6165 (
            .O(N__29287),
            .I(N__29281));
    InMux I__6164 (
            .O(N__29286),
            .I(N__29278));
    InMux I__6163 (
            .O(N__29285),
            .I(N__29274));
    InMux I__6162 (
            .O(N__29284),
            .I(N__29269));
    Span4Mux_v I__6161 (
            .O(N__29281),
            .I(N__29265));
    LocalMux I__6160 (
            .O(N__29278),
            .I(N__29262));
    InMux I__6159 (
            .O(N__29277),
            .I(N__29259));
    LocalMux I__6158 (
            .O(N__29274),
            .I(N__29256));
    InMux I__6157 (
            .O(N__29273),
            .I(N__29251));
    InMux I__6156 (
            .O(N__29272),
            .I(N__29251));
    LocalMux I__6155 (
            .O(N__29269),
            .I(N__29243));
    InMux I__6154 (
            .O(N__29268),
            .I(N__29240));
    Span4Mux_s1_v I__6153 (
            .O(N__29265),
            .I(N__29228));
    Span4Mux_v I__6152 (
            .O(N__29262),
            .I(N__29228));
    LocalMux I__6151 (
            .O(N__29259),
            .I(N__29228));
    Span4Mux_s3_h I__6150 (
            .O(N__29256),
            .I(N__29223));
    LocalMux I__6149 (
            .O(N__29251),
            .I(N__29223));
    CascadeMux I__6148 (
            .O(N__29250),
            .I(N__29218));
    CascadeMux I__6147 (
            .O(N__29249),
            .I(N__29211));
    CascadeMux I__6146 (
            .O(N__29248),
            .I(N__29208));
    CascadeMux I__6145 (
            .O(N__29247),
            .I(N__29205));
    CascadeMux I__6144 (
            .O(N__29246),
            .I(N__29202));
    Span4Mux_s2_v I__6143 (
            .O(N__29243),
            .I(N__29197));
    LocalMux I__6142 (
            .O(N__29240),
            .I(N__29194));
    InMux I__6141 (
            .O(N__29239),
            .I(N__29191));
    InMux I__6140 (
            .O(N__29238),
            .I(N__29186));
    InMux I__6139 (
            .O(N__29237),
            .I(N__29186));
    InMux I__6138 (
            .O(N__29236),
            .I(N__29183));
    InMux I__6137 (
            .O(N__29235),
            .I(N__29180));
    Span4Mux_h I__6136 (
            .O(N__29228),
            .I(N__29175));
    Span4Mux_h I__6135 (
            .O(N__29223),
            .I(N__29175));
    InMux I__6134 (
            .O(N__29222),
            .I(N__29164));
    InMux I__6133 (
            .O(N__29221),
            .I(N__29164));
    InMux I__6132 (
            .O(N__29218),
            .I(N__29164));
    InMux I__6131 (
            .O(N__29217),
            .I(N__29164));
    InMux I__6130 (
            .O(N__29216),
            .I(N__29164));
    InMux I__6129 (
            .O(N__29215),
            .I(N__29147));
    InMux I__6128 (
            .O(N__29214),
            .I(N__29147));
    InMux I__6127 (
            .O(N__29211),
            .I(N__29147));
    InMux I__6126 (
            .O(N__29208),
            .I(N__29147));
    InMux I__6125 (
            .O(N__29205),
            .I(N__29147));
    InMux I__6124 (
            .O(N__29202),
            .I(N__29147));
    InMux I__6123 (
            .O(N__29201),
            .I(N__29147));
    InMux I__6122 (
            .O(N__29200),
            .I(N__29147));
    Odrv4 I__6121 (
            .O(N__29197),
            .I(\b2v_inst11.N_3046_i ));
    Odrv12 I__6120 (
            .O(N__29194),
            .I(\b2v_inst11.N_3046_i ));
    LocalMux I__6119 (
            .O(N__29191),
            .I(\b2v_inst11.N_3046_i ));
    LocalMux I__6118 (
            .O(N__29186),
            .I(\b2v_inst11.N_3046_i ));
    LocalMux I__6117 (
            .O(N__29183),
            .I(\b2v_inst11.N_3046_i ));
    LocalMux I__6116 (
            .O(N__29180),
            .I(\b2v_inst11.N_3046_i ));
    Odrv4 I__6115 (
            .O(N__29175),
            .I(\b2v_inst11.N_3046_i ));
    LocalMux I__6114 (
            .O(N__29164),
            .I(\b2v_inst11.N_3046_i ));
    LocalMux I__6113 (
            .O(N__29147),
            .I(\b2v_inst11.N_3046_i ));
    InMux I__6112 (
            .O(N__29128),
            .I(N__29125));
    LocalMux I__6111 (
            .O(N__29125),
            .I(\b2v_inst11.g3_0 ));
    CascadeMux I__6110 (
            .O(N__29122),
            .I(\b2v_inst11.g2_0_cascade_ ));
    IoInMux I__6109 (
            .O(N__29119),
            .I(N__29116));
    LocalMux I__6108 (
            .O(N__29116),
            .I(N__29113));
    IoSpan4Mux I__6107 (
            .O(N__29113),
            .I(N__29108));
    InMux I__6106 (
            .O(N__29112),
            .I(N__29103));
    InMux I__6105 (
            .O(N__29111),
            .I(N__29103));
    Span4Mux_s3_h I__6104 (
            .O(N__29108),
            .I(N__29100));
    LocalMux I__6103 (
            .O(N__29103),
            .I(N__29096));
    Span4Mux_v I__6102 (
            .O(N__29100),
            .I(N__29089));
    InMux I__6101 (
            .O(N__29099),
            .I(N__29086));
    Sp12to4 I__6100 (
            .O(N__29096),
            .I(N__29082));
    InMux I__6099 (
            .O(N__29095),
            .I(N__29079));
    InMux I__6098 (
            .O(N__29094),
            .I(N__29076));
    InMux I__6097 (
            .O(N__29093),
            .I(N__29073));
    InMux I__6096 (
            .O(N__29092),
            .I(N__29068));
    Span4Mux_v I__6095 (
            .O(N__29089),
            .I(N__29063));
    LocalMux I__6094 (
            .O(N__29086),
            .I(N__29063));
    InMux I__6093 (
            .O(N__29085),
            .I(N__29060));
    Span12Mux_s7_h I__6092 (
            .O(N__29082),
            .I(N__29055));
    LocalMux I__6091 (
            .O(N__29079),
            .I(N__29055));
    LocalMux I__6090 (
            .O(N__29076),
            .I(N__29050));
    LocalMux I__6089 (
            .O(N__29073),
            .I(N__29050));
    InMux I__6088 (
            .O(N__29072),
            .I(N__29047));
    InMux I__6087 (
            .O(N__29071),
            .I(N__29044));
    LocalMux I__6086 (
            .O(N__29068),
            .I(N__29037));
    Span4Mux_h I__6085 (
            .O(N__29063),
            .I(N__29037));
    LocalMux I__6084 (
            .O(N__29060),
            .I(N__29037));
    Span12Mux_s2_v I__6083 (
            .O(N__29055),
            .I(N__29034));
    Odrv4 I__6082 (
            .O(N__29050),
            .I(RSMRSTn_RNI8DFE));
    LocalMux I__6081 (
            .O(N__29047),
            .I(RSMRSTn_RNI8DFE));
    LocalMux I__6080 (
            .O(N__29044),
            .I(RSMRSTn_RNI8DFE));
    Odrv4 I__6079 (
            .O(N__29037),
            .I(RSMRSTn_RNI8DFE));
    Odrv12 I__6078 (
            .O(N__29034),
            .I(RSMRSTn_RNI8DFE));
    InMux I__6077 (
            .O(N__29023),
            .I(N__29020));
    LocalMux I__6076 (
            .O(N__29020),
            .I(N__29017));
    Span4Mux_s3_v I__6075 (
            .O(N__29017),
            .I(N__29014));
    Odrv4 I__6074 (
            .O(N__29014),
            .I(\b2v_inst11.N_228_N_0 ));
    InMux I__6073 (
            .O(N__29011),
            .I(N__29008));
    LocalMux I__6072 (
            .O(N__29008),
            .I(N__29005));
    Odrv4 I__6071 (
            .O(N__29005),
            .I(\b2v_inst6.delayed_vccin_vccinaux_okZ0 ));
    InMux I__6070 (
            .O(N__29002),
            .I(N__28999));
    LocalMux I__6069 (
            .O(N__28999),
            .I(\b2v_inst11.g1_4_2_0 ));
    CascadeMux I__6068 (
            .O(N__28996),
            .I(N__28987));
    CascadeMux I__6067 (
            .O(N__28995),
            .I(N__28984));
    InMux I__6066 (
            .O(N__28994),
            .I(N__28981));
    InMux I__6065 (
            .O(N__28993),
            .I(N__28978));
    CascadeMux I__6064 (
            .O(N__28992),
            .I(N__28975));
    InMux I__6063 (
            .O(N__28991),
            .I(N__28966));
    InMux I__6062 (
            .O(N__28990),
            .I(N__28966));
    InMux I__6061 (
            .O(N__28987),
            .I(N__28963));
    InMux I__6060 (
            .O(N__28984),
            .I(N__28959));
    LocalMux I__6059 (
            .O(N__28981),
            .I(N__28950));
    LocalMux I__6058 (
            .O(N__28978),
            .I(N__28947));
    InMux I__6057 (
            .O(N__28975),
            .I(N__28944));
    CascadeMux I__6056 (
            .O(N__28974),
            .I(N__28941));
    CascadeMux I__6055 (
            .O(N__28973),
            .I(N__28937));
    InMux I__6054 (
            .O(N__28972),
            .I(N__28931));
    InMux I__6053 (
            .O(N__28971),
            .I(N__28927));
    LocalMux I__6052 (
            .O(N__28966),
            .I(N__28924));
    LocalMux I__6051 (
            .O(N__28963),
            .I(N__28921));
    CascadeMux I__6050 (
            .O(N__28962),
            .I(N__28918));
    LocalMux I__6049 (
            .O(N__28959),
            .I(N__28915));
    InMux I__6048 (
            .O(N__28958),
            .I(N__28910));
    InMux I__6047 (
            .O(N__28957),
            .I(N__28910));
    InMux I__6046 (
            .O(N__28956),
            .I(N__28901));
    InMux I__6045 (
            .O(N__28955),
            .I(N__28901));
    InMux I__6044 (
            .O(N__28954),
            .I(N__28901));
    InMux I__6043 (
            .O(N__28953),
            .I(N__28901));
    Span4Mux_v I__6042 (
            .O(N__28950),
            .I(N__28896));
    Span4Mux_v I__6041 (
            .O(N__28947),
            .I(N__28896));
    LocalMux I__6040 (
            .O(N__28944),
            .I(N__28893));
    InMux I__6039 (
            .O(N__28941),
            .I(N__28888));
    InMux I__6038 (
            .O(N__28940),
            .I(N__28888));
    InMux I__6037 (
            .O(N__28937),
            .I(N__28879));
    InMux I__6036 (
            .O(N__28936),
            .I(N__28879));
    InMux I__6035 (
            .O(N__28935),
            .I(N__28879));
    InMux I__6034 (
            .O(N__28934),
            .I(N__28879));
    LocalMux I__6033 (
            .O(N__28931),
            .I(N__28876));
    InMux I__6032 (
            .O(N__28930),
            .I(N__28873));
    LocalMux I__6031 (
            .O(N__28927),
            .I(N__28866));
    Span4Mux_v I__6030 (
            .O(N__28924),
            .I(N__28866));
    Span4Mux_s3_v I__6029 (
            .O(N__28921),
            .I(N__28866));
    InMux I__6028 (
            .O(N__28918),
            .I(N__28863));
    Span4Mux_v I__6027 (
            .O(N__28915),
            .I(N__28856));
    LocalMux I__6026 (
            .O(N__28910),
            .I(N__28856));
    LocalMux I__6025 (
            .O(N__28901),
            .I(N__28856));
    Odrv4 I__6024 (
            .O(N__28896),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    Odrv12 I__6023 (
            .O(N__28893),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    LocalMux I__6022 (
            .O(N__28888),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    LocalMux I__6021 (
            .O(N__28879),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    Odrv4 I__6020 (
            .O(N__28876),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    LocalMux I__6019 (
            .O(N__28873),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    Odrv4 I__6018 (
            .O(N__28866),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    LocalMux I__6017 (
            .O(N__28863),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    Odrv4 I__6016 (
            .O(N__28856),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    CascadeMux I__6015 (
            .O(N__28837),
            .I(N__28833));
    InMux I__6014 (
            .O(N__28836),
            .I(N__28825));
    InMux I__6013 (
            .O(N__28833),
            .I(N__28822));
    InMux I__6012 (
            .O(N__28832),
            .I(N__28819));
    InMux I__6011 (
            .O(N__28831),
            .I(N__28814));
    InMux I__6010 (
            .O(N__28830),
            .I(N__28814));
    InMux I__6009 (
            .O(N__28829),
            .I(N__28811));
    InMux I__6008 (
            .O(N__28828),
            .I(N__28808));
    LocalMux I__6007 (
            .O(N__28825),
            .I(N__28805));
    LocalMux I__6006 (
            .O(N__28822),
            .I(N__28802));
    LocalMux I__6005 (
            .O(N__28819),
            .I(N__28799));
    LocalMux I__6004 (
            .O(N__28814),
            .I(N__28795));
    LocalMux I__6003 (
            .O(N__28811),
            .I(N__28792));
    LocalMux I__6002 (
            .O(N__28808),
            .I(N__28789));
    Span4Mux_h I__6001 (
            .O(N__28805),
            .I(N__28784));
    Span4Mux_h I__6000 (
            .O(N__28802),
            .I(N__28784));
    Span4Mux_v I__5999 (
            .O(N__28799),
            .I(N__28781));
    InMux I__5998 (
            .O(N__28798),
            .I(N__28778));
    Span4Mux_v I__5997 (
            .O(N__28795),
            .I(N__28773));
    Span4Mux_v I__5996 (
            .O(N__28792),
            .I(N__28773));
    Odrv4 I__5995 (
            .O(N__28789),
            .I(N_19_i));
    Odrv4 I__5994 (
            .O(N__28784),
            .I(N_19_i));
    Odrv4 I__5993 (
            .O(N__28781),
            .I(N_19_i));
    LocalMux I__5992 (
            .O(N__28778),
            .I(N_19_i));
    Odrv4 I__5991 (
            .O(N__28773),
            .I(N_19_i));
    InMux I__5990 (
            .O(N__28762),
            .I(N__28756));
    InMux I__5989 (
            .O(N__28761),
            .I(N__28756));
    LocalMux I__5988 (
            .O(N__28756),
            .I(\b2v_inst11.g0_8_0_0 ));
    CascadeMux I__5987 (
            .O(N__28753),
            .I(N__28748));
    CascadeMux I__5986 (
            .O(N__28752),
            .I(N__28741));
    CascadeMux I__5985 (
            .O(N__28751),
            .I(N__28736));
    InMux I__5984 (
            .O(N__28748),
            .I(N__28733));
    InMux I__5983 (
            .O(N__28747),
            .I(N__28728));
    InMux I__5982 (
            .O(N__28746),
            .I(N__28725));
    InMux I__5981 (
            .O(N__28745),
            .I(N__28722));
    InMux I__5980 (
            .O(N__28744),
            .I(N__28717));
    InMux I__5979 (
            .O(N__28741),
            .I(N__28717));
    InMux I__5978 (
            .O(N__28740),
            .I(N__28712));
    InMux I__5977 (
            .O(N__28739),
            .I(N__28712));
    InMux I__5976 (
            .O(N__28736),
            .I(N__28709));
    LocalMux I__5975 (
            .O(N__28733),
            .I(N__28702));
    InMux I__5974 (
            .O(N__28732),
            .I(N__28697));
    InMux I__5973 (
            .O(N__28731),
            .I(N__28697));
    LocalMux I__5972 (
            .O(N__28728),
            .I(N__28692));
    LocalMux I__5971 (
            .O(N__28725),
            .I(N__28692));
    LocalMux I__5970 (
            .O(N__28722),
            .I(N__28685));
    LocalMux I__5969 (
            .O(N__28717),
            .I(N__28685));
    LocalMux I__5968 (
            .O(N__28712),
            .I(N__28685));
    LocalMux I__5967 (
            .O(N__28709),
            .I(N__28682));
    InMux I__5966 (
            .O(N__28708),
            .I(N__28679));
    InMux I__5965 (
            .O(N__28707),
            .I(N__28675));
    InMux I__5964 (
            .O(N__28706),
            .I(N__28669));
    InMux I__5963 (
            .O(N__28705),
            .I(N__28669));
    Span4Mux_v I__5962 (
            .O(N__28702),
            .I(N__28663));
    LocalMux I__5961 (
            .O(N__28697),
            .I(N__28663));
    Span4Mux_v I__5960 (
            .O(N__28692),
            .I(N__28654));
    Span4Mux_h I__5959 (
            .O(N__28685),
            .I(N__28654));
    Span4Mux_v I__5958 (
            .O(N__28682),
            .I(N__28654));
    LocalMux I__5957 (
            .O(N__28679),
            .I(N__28654));
    InMux I__5956 (
            .O(N__28678),
            .I(N__28651));
    LocalMux I__5955 (
            .O(N__28675),
            .I(N__28648));
    InMux I__5954 (
            .O(N__28674),
            .I(N__28645));
    LocalMux I__5953 (
            .O(N__28669),
            .I(N__28642));
    InMux I__5952 (
            .O(N__28668),
            .I(N__28639));
    IoSpan4Mux I__5951 (
            .O(N__28663),
            .I(N__28636));
    Span4Mux_h I__5950 (
            .O(N__28654),
            .I(N__28633));
    LocalMux I__5949 (
            .O(N__28651),
            .I(N__28630));
    Span4Mux_h I__5948 (
            .O(N__28648),
            .I(N__28625));
    LocalMux I__5947 (
            .O(N__28645),
            .I(N__28625));
    Span4Mux_h I__5946 (
            .O(N__28642),
            .I(N__28620));
    LocalMux I__5945 (
            .O(N__28639),
            .I(N__28620));
    IoSpan4Mux I__5944 (
            .O(N__28636),
            .I(N__28617));
    Span4Mux_v I__5943 (
            .O(N__28633),
            .I(N__28614));
    IoSpan4Mux I__5942 (
            .O(N__28630),
            .I(N__28611));
    IoSpan4Mux I__5941 (
            .O(N__28625),
            .I(N__28606));
    IoSpan4Mux I__5940 (
            .O(N__28620),
            .I(N__28606));
    Odrv4 I__5939 (
            .O(N__28617),
            .I(SLP_S4n_c));
    Odrv4 I__5938 (
            .O(N__28614),
            .I(SLP_S4n_c));
    Odrv4 I__5937 (
            .O(N__28611),
            .I(SLP_S4n_c));
    Odrv4 I__5936 (
            .O(N__28606),
            .I(SLP_S4n_c));
    InMux I__5935 (
            .O(N__28597),
            .I(N__28594));
    LocalMux I__5934 (
            .O(N__28594),
            .I(N__28588));
    InMux I__5933 (
            .O(N__28593),
            .I(N__28583));
    InMux I__5932 (
            .O(N__28592),
            .I(N__28583));
    InMux I__5931 (
            .O(N__28591),
            .I(N__28578));
    Span4Mux_h I__5930 (
            .O(N__28588),
            .I(N__28567));
    LocalMux I__5929 (
            .O(N__28583),
            .I(N__28567));
    InMux I__5928 (
            .O(N__28582),
            .I(N__28564));
    InMux I__5927 (
            .O(N__28581),
            .I(N__28561));
    LocalMux I__5926 (
            .O(N__28578),
            .I(N__28556));
    InMux I__5925 (
            .O(N__28577),
            .I(N__28553));
    InMux I__5924 (
            .O(N__28576),
            .I(N__28550));
    InMux I__5923 (
            .O(N__28575),
            .I(N__28545));
    InMux I__5922 (
            .O(N__28574),
            .I(N__28542));
    InMux I__5921 (
            .O(N__28573),
            .I(N__28539));
    InMux I__5920 (
            .O(N__28572),
            .I(N__28536));
    Span4Mux_v I__5919 (
            .O(N__28567),
            .I(N__28529));
    LocalMux I__5918 (
            .O(N__28564),
            .I(N__28529));
    LocalMux I__5917 (
            .O(N__28561),
            .I(N__28529));
    InMux I__5916 (
            .O(N__28560),
            .I(N__28524));
    InMux I__5915 (
            .O(N__28559),
            .I(N__28524));
    Span4Mux_v I__5914 (
            .O(N__28556),
            .I(N__28519));
    LocalMux I__5913 (
            .O(N__28553),
            .I(N__28519));
    LocalMux I__5912 (
            .O(N__28550),
            .I(N__28516));
    InMux I__5911 (
            .O(N__28549),
            .I(N__28511));
    InMux I__5910 (
            .O(N__28548),
            .I(N__28511));
    LocalMux I__5909 (
            .O(N__28545),
            .I(N__28504));
    LocalMux I__5908 (
            .O(N__28542),
            .I(N__28504));
    LocalMux I__5907 (
            .O(N__28539),
            .I(N__28504));
    LocalMux I__5906 (
            .O(N__28536),
            .I(N__28501));
    Span4Mux_h I__5905 (
            .O(N__28529),
            .I(N__28496));
    LocalMux I__5904 (
            .O(N__28524),
            .I(N__28496));
    Span4Mux_v I__5903 (
            .O(N__28519),
            .I(N__28489));
    Span4Mux_h I__5902 (
            .O(N__28516),
            .I(N__28489));
    LocalMux I__5901 (
            .O(N__28511),
            .I(N__28489));
    Span12Mux_s9_h I__5900 (
            .O(N__28504),
            .I(N__28485));
    Span4Mux_v I__5899 (
            .O(N__28501),
            .I(N__28482));
    IoSpan4Mux I__5898 (
            .O(N__28496),
            .I(N__28479));
    Span4Mux_h I__5897 (
            .O(N__28489),
            .I(N__28476));
    InMux I__5896 (
            .O(N__28488),
            .I(N__28473));
    Odrv12 I__5895 (
            .O(N__28485),
            .I(GPIO_FPGA_PCH_5_c));
    Odrv4 I__5894 (
            .O(N__28482),
            .I(GPIO_FPGA_PCH_5_c));
    Odrv4 I__5893 (
            .O(N__28479),
            .I(GPIO_FPGA_PCH_5_c));
    Odrv4 I__5892 (
            .O(N__28476),
            .I(GPIO_FPGA_PCH_5_c));
    LocalMux I__5891 (
            .O(N__28473),
            .I(GPIO_FPGA_PCH_5_c));
    InMux I__5890 (
            .O(N__28462),
            .I(N__28447));
    InMux I__5889 (
            .O(N__28461),
            .I(N__28447));
    InMux I__5888 (
            .O(N__28460),
            .I(N__28447));
    InMux I__5887 (
            .O(N__28459),
            .I(N__28440));
    InMux I__5886 (
            .O(N__28458),
            .I(N__28440));
    InMux I__5885 (
            .O(N__28457),
            .I(N__28440));
    InMux I__5884 (
            .O(N__28456),
            .I(N__28435));
    InMux I__5883 (
            .O(N__28455),
            .I(N__28435));
    InMux I__5882 (
            .O(N__28454),
            .I(N__28430));
    LocalMux I__5881 (
            .O(N__28447),
            .I(N__28426));
    LocalMux I__5880 (
            .O(N__28440),
            .I(N__28423));
    LocalMux I__5879 (
            .O(N__28435),
            .I(N__28420));
    InMux I__5878 (
            .O(N__28434),
            .I(N__28417));
    CascadeMux I__5877 (
            .O(N__28433),
            .I(N__28414));
    LocalMux I__5876 (
            .O(N__28430),
            .I(N__28409));
    InMux I__5875 (
            .O(N__28429),
            .I(N__28406));
    Span4Mux_s3_v I__5874 (
            .O(N__28426),
            .I(N__28396));
    Span4Mux_s3_h I__5873 (
            .O(N__28423),
            .I(N__28396));
    Span4Mux_v I__5872 (
            .O(N__28420),
            .I(N__28396));
    LocalMux I__5871 (
            .O(N__28417),
            .I(N__28392));
    InMux I__5870 (
            .O(N__28414),
            .I(N__28389));
    InMux I__5869 (
            .O(N__28413),
            .I(N__28386));
    InMux I__5868 (
            .O(N__28412),
            .I(N__28383));
    Span4Mux_s3_v I__5867 (
            .O(N__28409),
            .I(N__28378));
    LocalMux I__5866 (
            .O(N__28406),
            .I(N__28378));
    InMux I__5865 (
            .O(N__28405),
            .I(N__28371));
    InMux I__5864 (
            .O(N__28404),
            .I(N__28371));
    InMux I__5863 (
            .O(N__28403),
            .I(N__28371));
    Span4Mux_h I__5862 (
            .O(N__28396),
            .I(N__28368));
    InMux I__5861 (
            .O(N__28395),
            .I(N__28365));
    Odrv4 I__5860 (
            .O(N__28392),
            .I(\b2v_inst11.func_state ));
    LocalMux I__5859 (
            .O(N__28389),
            .I(\b2v_inst11.func_state ));
    LocalMux I__5858 (
            .O(N__28386),
            .I(\b2v_inst11.func_state ));
    LocalMux I__5857 (
            .O(N__28383),
            .I(\b2v_inst11.func_state ));
    Odrv4 I__5856 (
            .O(N__28378),
            .I(\b2v_inst11.func_state ));
    LocalMux I__5855 (
            .O(N__28371),
            .I(\b2v_inst11.func_state ));
    Odrv4 I__5854 (
            .O(N__28368),
            .I(\b2v_inst11.func_state ));
    LocalMux I__5853 (
            .O(N__28365),
            .I(\b2v_inst11.func_state ));
    InMux I__5852 (
            .O(N__28348),
            .I(N__28340));
    InMux I__5851 (
            .O(N__28347),
            .I(N__28337));
    CascadeMux I__5850 (
            .O(N__28346),
            .I(N__28333));
    CascadeMux I__5849 (
            .O(N__28345),
            .I(N__28329));
    CascadeMux I__5848 (
            .O(N__28344),
            .I(N__28326));
    CascadeMux I__5847 (
            .O(N__28343),
            .I(N__28323));
    LocalMux I__5846 (
            .O(N__28340),
            .I(N__28317));
    LocalMux I__5845 (
            .O(N__28337),
            .I(N__28317));
    InMux I__5844 (
            .O(N__28336),
            .I(N__28312));
    InMux I__5843 (
            .O(N__28333),
            .I(N__28312));
    InMux I__5842 (
            .O(N__28332),
            .I(N__28304));
    InMux I__5841 (
            .O(N__28329),
            .I(N__28301));
    InMux I__5840 (
            .O(N__28326),
            .I(N__28298));
    InMux I__5839 (
            .O(N__28323),
            .I(N__28293));
    InMux I__5838 (
            .O(N__28322),
            .I(N__28293));
    Span4Mux_h I__5837 (
            .O(N__28317),
            .I(N__28287));
    LocalMux I__5836 (
            .O(N__28312),
            .I(N__28284));
    InMux I__5835 (
            .O(N__28311),
            .I(N__28277));
    InMux I__5834 (
            .O(N__28310),
            .I(N__28277));
    InMux I__5833 (
            .O(N__28309),
            .I(N__28277));
    CascadeMux I__5832 (
            .O(N__28308),
            .I(N__28273));
    InMux I__5831 (
            .O(N__28307),
            .I(N__28270));
    LocalMux I__5830 (
            .O(N__28304),
            .I(N__28265));
    LocalMux I__5829 (
            .O(N__28301),
            .I(N__28265));
    LocalMux I__5828 (
            .O(N__28298),
            .I(N__28260));
    LocalMux I__5827 (
            .O(N__28293),
            .I(N__28260));
    InMux I__5826 (
            .O(N__28292),
            .I(N__28257));
    InMux I__5825 (
            .O(N__28291),
            .I(N__28254));
    CascadeMux I__5824 (
            .O(N__28290),
            .I(N__28249));
    Span4Mux_v I__5823 (
            .O(N__28287),
            .I(N__28244));
    Span4Mux_h I__5822 (
            .O(N__28284),
            .I(N__28244));
    LocalMux I__5821 (
            .O(N__28277),
            .I(N__28241));
    InMux I__5820 (
            .O(N__28276),
            .I(N__28238));
    InMux I__5819 (
            .O(N__28273),
            .I(N__28235));
    LocalMux I__5818 (
            .O(N__28270),
            .I(N__28232));
    Span4Mux_h I__5817 (
            .O(N__28265),
            .I(N__28223));
    Span4Mux_h I__5816 (
            .O(N__28260),
            .I(N__28223));
    LocalMux I__5815 (
            .O(N__28257),
            .I(N__28223));
    LocalMux I__5814 (
            .O(N__28254),
            .I(N__28223));
    InMux I__5813 (
            .O(N__28253),
            .I(N__28220));
    InMux I__5812 (
            .O(N__28252),
            .I(N__28216));
    InMux I__5811 (
            .O(N__28249),
            .I(N__28213));
    IoSpan4Mux I__5810 (
            .O(N__28244),
            .I(N__28210));
    Span4Mux_v I__5809 (
            .O(N__28241),
            .I(N__28203));
    LocalMux I__5808 (
            .O(N__28238),
            .I(N__28203));
    LocalMux I__5807 (
            .O(N__28235),
            .I(N__28203));
    Span4Mux_v I__5806 (
            .O(N__28232),
            .I(N__28196));
    Span4Mux_h I__5805 (
            .O(N__28223),
            .I(N__28196));
    LocalMux I__5804 (
            .O(N__28220),
            .I(N__28196));
    InMux I__5803 (
            .O(N__28219),
            .I(N__28193));
    LocalMux I__5802 (
            .O(N__28216),
            .I(N__28188));
    LocalMux I__5801 (
            .O(N__28213),
            .I(N__28188));
    Span4Mux_s0_v I__5800 (
            .O(N__28210),
            .I(N__28179));
    Span4Mux_h I__5799 (
            .O(N__28203),
            .I(N__28179));
    Span4Mux_v I__5798 (
            .O(N__28196),
            .I(N__28179));
    LocalMux I__5797 (
            .O(N__28193),
            .I(N__28179));
    Span12Mux_s10_h I__5796 (
            .O(N__28188),
            .I(N__28176));
    Span4Mux_h I__5795 (
            .O(N__28179),
            .I(N__28173));
    Odrv12 I__5794 (
            .O(N__28176),
            .I(SLP_S3n_c));
    Odrv4 I__5793 (
            .O(N__28173),
            .I(SLP_S3n_c));
    InMux I__5792 (
            .O(N__28168),
            .I(N__28160));
    InMux I__5791 (
            .O(N__28167),
            .I(N__28154));
    InMux I__5790 (
            .O(N__28166),
            .I(N__28148));
    InMux I__5789 (
            .O(N__28165),
            .I(N__28148));
    InMux I__5788 (
            .O(N__28164),
            .I(N__28143));
    InMux I__5787 (
            .O(N__28163),
            .I(N__28143));
    LocalMux I__5786 (
            .O(N__28160),
            .I(N__28137));
    InMux I__5785 (
            .O(N__28159),
            .I(N__28130));
    InMux I__5784 (
            .O(N__28158),
            .I(N__28130));
    InMux I__5783 (
            .O(N__28157),
            .I(N__28130));
    LocalMux I__5782 (
            .O(N__28154),
            .I(N__28127));
    InMux I__5781 (
            .O(N__28153),
            .I(N__28124));
    LocalMux I__5780 (
            .O(N__28148),
            .I(N__28119));
    LocalMux I__5779 (
            .O(N__28143),
            .I(N__28119));
    InMux I__5778 (
            .O(N__28142),
            .I(N__28114));
    InMux I__5777 (
            .O(N__28141),
            .I(N__28111));
    InMux I__5776 (
            .O(N__28140),
            .I(N__28108));
    Span4Mux_v I__5775 (
            .O(N__28137),
            .I(N__28102));
    LocalMux I__5774 (
            .O(N__28130),
            .I(N__28102));
    Span4Mux_v I__5773 (
            .O(N__28127),
            .I(N__28097));
    LocalMux I__5772 (
            .O(N__28124),
            .I(N__28097));
    Span4Mux_v I__5771 (
            .O(N__28119),
            .I(N__28093));
    InMux I__5770 (
            .O(N__28118),
            .I(N__28090));
    InMux I__5769 (
            .O(N__28117),
            .I(N__28087));
    LocalMux I__5768 (
            .O(N__28114),
            .I(N__28080));
    LocalMux I__5767 (
            .O(N__28111),
            .I(N__28080));
    LocalMux I__5766 (
            .O(N__28108),
            .I(N__28080));
    InMux I__5765 (
            .O(N__28107),
            .I(N__28077));
    Span4Mux_s2_v I__5764 (
            .O(N__28102),
            .I(N__28074));
    Span4Mux_h I__5763 (
            .O(N__28097),
            .I(N__28071));
    InMux I__5762 (
            .O(N__28096),
            .I(N__28068));
    Sp12to4 I__5761 (
            .O(N__28093),
            .I(N__28063));
    LocalMux I__5760 (
            .O(N__28090),
            .I(N__28063));
    LocalMux I__5759 (
            .O(N__28087),
            .I(N__28056));
    Span4Mux_v I__5758 (
            .O(N__28080),
            .I(N__28056));
    LocalMux I__5757 (
            .O(N__28077),
            .I(N__28056));
    Span4Mux_h I__5756 (
            .O(N__28074),
            .I(N__28053));
    Span4Mux_h I__5755 (
            .O(N__28071),
            .I(N__28048));
    LocalMux I__5754 (
            .O(N__28068),
            .I(N__28048));
    Odrv12 I__5753 (
            .O(N__28063),
            .I(\b2v_inst11.count_clk_RNIZ0Z_3 ));
    Odrv4 I__5752 (
            .O(N__28056),
            .I(\b2v_inst11.count_clk_RNIZ0Z_3 ));
    Odrv4 I__5751 (
            .O(N__28053),
            .I(\b2v_inst11.count_clk_RNIZ0Z_3 ));
    Odrv4 I__5750 (
            .O(N__28048),
            .I(\b2v_inst11.count_clk_RNIZ0Z_3 ));
    CascadeMux I__5749 (
            .O(N__28039),
            .I(\b2v_inst11.g1_2_1_cascade_ ));
    CascadeMux I__5748 (
            .O(N__28036),
            .I(N__28033));
    InMux I__5747 (
            .O(N__28033),
            .I(N__28025));
    CascadeMux I__5746 (
            .O(N__28032),
            .I(N__28021));
    InMux I__5745 (
            .O(N__28031),
            .I(N__28003));
    InMux I__5744 (
            .O(N__28030),
            .I(N__28003));
    InMux I__5743 (
            .O(N__28029),
            .I(N__28003));
    CascadeMux I__5742 (
            .O(N__28028),
            .I(N__28000));
    LocalMux I__5741 (
            .O(N__28025),
            .I(N__27996));
    InMux I__5740 (
            .O(N__28024),
            .I(N__27991));
    InMux I__5739 (
            .O(N__28021),
            .I(N__27991));
    CascadeMux I__5738 (
            .O(N__28020),
            .I(N__27988));
    InMux I__5737 (
            .O(N__28019),
            .I(N__27982));
    InMux I__5736 (
            .O(N__28018),
            .I(N__27975));
    InMux I__5735 (
            .O(N__28017),
            .I(N__27975));
    InMux I__5734 (
            .O(N__28016),
            .I(N__27975));
    InMux I__5733 (
            .O(N__28015),
            .I(N__27972));
    InMux I__5732 (
            .O(N__28014),
            .I(N__27969));
    CascadeMux I__5731 (
            .O(N__28013),
            .I(N__27966));
    InMux I__5730 (
            .O(N__28012),
            .I(N__27958));
    InMux I__5729 (
            .O(N__28011),
            .I(N__27958));
    InMux I__5728 (
            .O(N__28010),
            .I(N__27958));
    LocalMux I__5727 (
            .O(N__28003),
            .I(N__27953));
    InMux I__5726 (
            .O(N__28000),
            .I(N__27950));
    InMux I__5725 (
            .O(N__27999),
            .I(N__27947));
    Span4Mux_v I__5724 (
            .O(N__27996),
            .I(N__27942));
    LocalMux I__5723 (
            .O(N__27991),
            .I(N__27942));
    InMux I__5722 (
            .O(N__27988),
            .I(N__27939));
    InMux I__5721 (
            .O(N__27987),
            .I(N__27936));
    InMux I__5720 (
            .O(N__27986),
            .I(N__27931));
    InMux I__5719 (
            .O(N__27985),
            .I(N__27931));
    LocalMux I__5718 (
            .O(N__27982),
            .I(N__27928));
    LocalMux I__5717 (
            .O(N__27975),
            .I(N__27921));
    LocalMux I__5716 (
            .O(N__27972),
            .I(N__27921));
    LocalMux I__5715 (
            .O(N__27969),
            .I(N__27921));
    InMux I__5714 (
            .O(N__27966),
            .I(N__27916));
    InMux I__5713 (
            .O(N__27965),
            .I(N__27916));
    LocalMux I__5712 (
            .O(N__27958),
            .I(N__27913));
    InMux I__5711 (
            .O(N__27957),
            .I(N__27909));
    InMux I__5710 (
            .O(N__27956),
            .I(N__27906));
    Span4Mux_v I__5709 (
            .O(N__27953),
            .I(N__27897));
    LocalMux I__5708 (
            .O(N__27950),
            .I(N__27897));
    LocalMux I__5707 (
            .O(N__27947),
            .I(N__27897));
    Span4Mux_v I__5706 (
            .O(N__27942),
            .I(N__27897));
    LocalMux I__5705 (
            .O(N__27939),
            .I(N__27890));
    LocalMux I__5704 (
            .O(N__27936),
            .I(N__27890));
    LocalMux I__5703 (
            .O(N__27931),
            .I(N__27890));
    Span4Mux_v I__5702 (
            .O(N__27928),
            .I(N__27883));
    Span4Mux_h I__5701 (
            .O(N__27921),
            .I(N__27883));
    LocalMux I__5700 (
            .O(N__27916),
            .I(N__27883));
    Span4Mux_h I__5699 (
            .O(N__27913),
            .I(N__27880));
    InMux I__5698 (
            .O(N__27912),
            .I(N__27877));
    LocalMux I__5697 (
            .O(N__27909),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    LocalMux I__5696 (
            .O(N__27906),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv4 I__5695 (
            .O(N__27897),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv4 I__5694 (
            .O(N__27890),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv4 I__5693 (
            .O(N__27883),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv4 I__5692 (
            .O(N__27880),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    LocalMux I__5691 (
            .O(N__27877),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    InMux I__5690 (
            .O(N__27862),
            .I(N__27859));
    LocalMux I__5689 (
            .O(N__27859),
            .I(N__27856));
    Odrv4 I__5688 (
            .O(N__27856),
            .I(\b2v_inst11.g1_2 ));
    CascadeMux I__5687 (
            .O(N__27853),
            .I(\b2v_inst6.countZ0Z_11_cascade_ ));
    InMux I__5686 (
            .O(N__27850),
            .I(N__27847));
    LocalMux I__5685 (
            .O(N__27847),
            .I(\b2v_inst6.count_3_11 ));
    CascadeMux I__5684 (
            .O(N__27844),
            .I(N__27840));
    InMux I__5683 (
            .O(N__27843),
            .I(N__27835));
    InMux I__5682 (
            .O(N__27840),
            .I(N__27835));
    LocalMux I__5681 (
            .O(N__27835),
            .I(\b2v_inst6.curr_state_RNIDMSJ1Z0Z_1 ));
    InMux I__5680 (
            .O(N__27832),
            .I(N__27829));
    LocalMux I__5679 (
            .O(N__27829),
            .I(b2v_inst11_count_off_1_sqmuxa_0_0_0));
    InMux I__5678 (
            .O(N__27826),
            .I(N__27823));
    LocalMux I__5677 (
            .O(N__27823),
            .I(G_26_0_a5_1_0));
    CascadeMux I__5676 (
            .O(N__27820),
            .I(G_26_0_a5_2_1_cascade_));
    InMux I__5675 (
            .O(N__27817),
            .I(N__27814));
    LocalMux I__5674 (
            .O(N__27814),
            .I(G_26_0_0));
    InMux I__5673 (
            .O(N__27811),
            .I(N__27808));
    LocalMux I__5672 (
            .O(N__27808),
            .I(N__27805));
    Span4Mux_h I__5671 (
            .O(N__27805),
            .I(N__27802));
    Odrv4 I__5670 (
            .O(N__27802),
            .I(\b2v_inst11.g2_0_1 ));
    InMux I__5669 (
            .O(N__27799),
            .I(N__27796));
    LocalMux I__5668 (
            .O(N__27796),
            .I(\b2v_inst11.un1_dutycycle_172_m4 ));
    CascadeMux I__5667 (
            .O(N__27793),
            .I(b2v_inst11_un1_dutycycle_172_m3_0_0_0_cascade_));
    InMux I__5666 (
            .O(N__27790),
            .I(N__27787));
    LocalMux I__5665 (
            .O(N__27787),
            .I(N__27784));
    Odrv4 I__5664 (
            .O(N__27784),
            .I(\b2v_inst11.g2_1 ));
    CascadeMux I__5663 (
            .O(N__27781),
            .I(N__27773));
    InMux I__5662 (
            .O(N__27780),
            .I(N__27767));
    InMux I__5661 (
            .O(N__27779),
            .I(N__27764));
    InMux I__5660 (
            .O(N__27778),
            .I(N__27761));
    InMux I__5659 (
            .O(N__27777),
            .I(N__27755));
    InMux I__5658 (
            .O(N__27776),
            .I(N__27747));
    InMux I__5657 (
            .O(N__27773),
            .I(N__27742));
    InMux I__5656 (
            .O(N__27772),
            .I(N__27742));
    InMux I__5655 (
            .O(N__27771),
            .I(N__27738));
    InMux I__5654 (
            .O(N__27770),
            .I(N__27735));
    LocalMux I__5653 (
            .O(N__27767),
            .I(N__27728));
    LocalMux I__5652 (
            .O(N__27764),
            .I(N__27728));
    LocalMux I__5651 (
            .O(N__27761),
            .I(N__27728));
    InMux I__5650 (
            .O(N__27760),
            .I(N__27721));
    InMux I__5649 (
            .O(N__27759),
            .I(N__27721));
    InMux I__5648 (
            .O(N__27758),
            .I(N__27721));
    LocalMux I__5647 (
            .O(N__27755),
            .I(N__27718));
    InMux I__5646 (
            .O(N__27754),
            .I(N__27715));
    InMux I__5645 (
            .O(N__27753),
            .I(N__27710));
    InMux I__5644 (
            .O(N__27752),
            .I(N__27710));
    InMux I__5643 (
            .O(N__27751),
            .I(N__27707));
    InMux I__5642 (
            .O(N__27750),
            .I(N__27704));
    LocalMux I__5641 (
            .O(N__27747),
            .I(N__27699));
    LocalMux I__5640 (
            .O(N__27742),
            .I(N__27699));
    CascadeMux I__5639 (
            .O(N__27741),
            .I(N__27696));
    LocalMux I__5638 (
            .O(N__27738),
            .I(N__27689));
    LocalMux I__5637 (
            .O(N__27735),
            .I(N__27686));
    Span4Mux_v I__5636 (
            .O(N__27728),
            .I(N__27681));
    LocalMux I__5635 (
            .O(N__27721),
            .I(N__27681));
    Span4Mux_h I__5634 (
            .O(N__27718),
            .I(N__27676));
    LocalMux I__5633 (
            .O(N__27715),
            .I(N__27676));
    LocalMux I__5632 (
            .O(N__27710),
            .I(N__27667));
    LocalMux I__5631 (
            .O(N__27707),
            .I(N__27667));
    LocalMux I__5630 (
            .O(N__27704),
            .I(N__27667));
    Span4Mux_s2_v I__5629 (
            .O(N__27699),
            .I(N__27667));
    InMux I__5628 (
            .O(N__27696),
            .I(N__27664));
    InMux I__5627 (
            .O(N__27695),
            .I(N__27661));
    InMux I__5626 (
            .O(N__27694),
            .I(N__27654));
    InMux I__5625 (
            .O(N__27693),
            .I(N__27654));
    InMux I__5624 (
            .O(N__27692),
            .I(N__27654));
    Span4Mux_s3_v I__5623 (
            .O(N__27689),
            .I(N__27645));
    Span4Mux_s3_v I__5622 (
            .O(N__27686),
            .I(N__27645));
    Span4Mux_h I__5621 (
            .O(N__27681),
            .I(N__27645));
    Span4Mux_h I__5620 (
            .O(N__27676),
            .I(N__27645));
    Span4Mux_v I__5619 (
            .O(N__27667),
            .I(N__27642));
    LocalMux I__5618 (
            .O(N__27664),
            .I(N__27637));
    LocalMux I__5617 (
            .O(N__27661),
            .I(N__27637));
    LocalMux I__5616 (
            .O(N__27654),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z2 ));
    Odrv4 I__5615 (
            .O(N__27645),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z2 ));
    Odrv4 I__5614 (
            .O(N__27642),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z2 ));
    Odrv4 I__5613 (
            .O(N__27637),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z2 ));
    CascadeMux I__5612 (
            .O(N__27628),
            .I(\b2v_inst11.g4_cascade_ ));
    IoInMux I__5611 (
            .O(N__27625),
            .I(N__27621));
    InMux I__5610 (
            .O(N__27624),
            .I(N__27614));
    LocalMux I__5609 (
            .O(N__27621),
            .I(N__27611));
    CascadeMux I__5608 (
            .O(N__27620),
            .I(N__27607));
    InMux I__5607 (
            .O(N__27619),
            .I(N__27600));
    InMux I__5606 (
            .O(N__27618),
            .I(N__27588));
    InMux I__5605 (
            .O(N__27617),
            .I(N__27588));
    LocalMux I__5604 (
            .O(N__27614),
            .I(N__27582));
    IoSpan4Mux I__5603 (
            .O(N__27611),
            .I(N__27582));
    InMux I__5602 (
            .O(N__27610),
            .I(N__27575));
    InMux I__5601 (
            .O(N__27607),
            .I(N__27575));
    InMux I__5600 (
            .O(N__27606),
            .I(N__27575));
    InMux I__5599 (
            .O(N__27605),
            .I(N__27570));
    InMux I__5598 (
            .O(N__27604),
            .I(N__27570));
    InMux I__5597 (
            .O(N__27603),
            .I(N__27567));
    LocalMux I__5596 (
            .O(N__27600),
            .I(N__27564));
    InMux I__5595 (
            .O(N__27599),
            .I(N__27561));
    InMux I__5594 (
            .O(N__27598),
            .I(N__27558));
    InMux I__5593 (
            .O(N__27597),
            .I(N__27551));
    InMux I__5592 (
            .O(N__27596),
            .I(N__27551));
    InMux I__5591 (
            .O(N__27595),
            .I(N__27551));
    InMux I__5590 (
            .O(N__27594),
            .I(N__27540));
    InMux I__5589 (
            .O(N__27593),
            .I(N__27540));
    LocalMux I__5588 (
            .O(N__27588),
            .I(N__27537));
    InMux I__5587 (
            .O(N__27587),
            .I(N__27532));
    Span4Mux_s3_v I__5586 (
            .O(N__27582),
            .I(N__27529));
    LocalMux I__5585 (
            .O(N__27575),
            .I(N__27524));
    LocalMux I__5584 (
            .O(N__27570),
            .I(N__27524));
    LocalMux I__5583 (
            .O(N__27567),
            .I(N__27521));
    Span4Mux_s3_v I__5582 (
            .O(N__27564),
            .I(N__27514));
    LocalMux I__5581 (
            .O(N__27561),
            .I(N__27514));
    LocalMux I__5580 (
            .O(N__27558),
            .I(N__27514));
    LocalMux I__5579 (
            .O(N__27551),
            .I(N__27511));
    InMux I__5578 (
            .O(N__27550),
            .I(N__27504));
    InMux I__5577 (
            .O(N__27549),
            .I(N__27504));
    InMux I__5576 (
            .O(N__27548),
            .I(N__27504));
    InMux I__5575 (
            .O(N__27547),
            .I(N__27499));
    InMux I__5574 (
            .O(N__27546),
            .I(N__27499));
    InMux I__5573 (
            .O(N__27545),
            .I(N__27496));
    LocalMux I__5572 (
            .O(N__27540),
            .I(N__27493));
    Span4Mux_h I__5571 (
            .O(N__27537),
            .I(N__27490));
    InMux I__5570 (
            .O(N__27536),
            .I(N__27485));
    InMux I__5569 (
            .O(N__27535),
            .I(N__27485));
    LocalMux I__5568 (
            .O(N__27532),
            .I(N__27482));
    Span4Mux_h I__5567 (
            .O(N__27529),
            .I(N__27467));
    Span4Mux_s3_v I__5566 (
            .O(N__27524),
            .I(N__27467));
    Span4Mux_s3_v I__5565 (
            .O(N__27521),
            .I(N__27467));
    Span4Mux_h I__5564 (
            .O(N__27514),
            .I(N__27467));
    Span4Mux_h I__5563 (
            .O(N__27511),
            .I(N__27467));
    LocalMux I__5562 (
            .O(N__27504),
            .I(N__27467));
    LocalMux I__5561 (
            .O(N__27499),
            .I(N__27467));
    LocalMux I__5560 (
            .O(N__27496),
            .I(N__27464));
    Odrv4 I__5559 (
            .O(N__27493),
            .I(b2v_inst16_delayed_vddq_pwrgd_en));
    Odrv4 I__5558 (
            .O(N__27490),
            .I(b2v_inst16_delayed_vddq_pwrgd_en));
    LocalMux I__5557 (
            .O(N__27485),
            .I(b2v_inst16_delayed_vddq_pwrgd_en));
    Odrv12 I__5556 (
            .O(N__27482),
            .I(b2v_inst16_delayed_vddq_pwrgd_en));
    Odrv4 I__5555 (
            .O(N__27467),
            .I(b2v_inst16_delayed_vddq_pwrgd_en));
    Odrv4 I__5554 (
            .O(N__27464),
            .I(b2v_inst16_delayed_vddq_pwrgd_en));
    InMux I__5553 (
            .O(N__27451),
            .I(N__27445));
    InMux I__5552 (
            .O(N__27450),
            .I(N__27445));
    LocalMux I__5551 (
            .O(N__27445),
            .I(\b2v_inst11.N_5 ));
    InMux I__5550 (
            .O(N__27442),
            .I(N__27439));
    LocalMux I__5549 (
            .O(N__27439),
            .I(\b2v_inst11.un1_clk_100khz_52_and_i_a2_1_xZ0 ));
    CascadeMux I__5548 (
            .O(N__27436),
            .I(N__27432));
    CascadeMux I__5547 (
            .O(N__27435),
            .I(N__27429));
    InMux I__5546 (
            .O(N__27432),
            .I(N__27423));
    InMux I__5545 (
            .O(N__27429),
            .I(N__27418));
    InMux I__5544 (
            .O(N__27428),
            .I(N__27418));
    CascadeMux I__5543 (
            .O(N__27427),
            .I(N__27414));
    InMux I__5542 (
            .O(N__27426),
            .I(N__27410));
    LocalMux I__5541 (
            .O(N__27423),
            .I(N__27403));
    LocalMux I__5540 (
            .O(N__27418),
            .I(N__27403));
    InMux I__5539 (
            .O(N__27417),
            .I(N__27400));
    InMux I__5538 (
            .O(N__27414),
            .I(N__27397));
    CascadeMux I__5537 (
            .O(N__27413),
            .I(N__27394));
    LocalMux I__5536 (
            .O(N__27410),
            .I(N__27391));
    InMux I__5535 (
            .O(N__27409),
            .I(N__27386));
    InMux I__5534 (
            .O(N__27408),
            .I(N__27383));
    Span4Mux_v I__5533 (
            .O(N__27403),
            .I(N__27379));
    LocalMux I__5532 (
            .O(N__27400),
            .I(N__27374));
    LocalMux I__5531 (
            .O(N__27397),
            .I(N__27374));
    InMux I__5530 (
            .O(N__27394),
            .I(N__27371));
    Span12Mux_v I__5529 (
            .O(N__27391),
            .I(N__27368));
    InMux I__5528 (
            .O(N__27390),
            .I(N__27365));
    InMux I__5527 (
            .O(N__27389),
            .I(N__27362));
    LocalMux I__5526 (
            .O(N__27386),
            .I(N__27359));
    LocalMux I__5525 (
            .O(N__27383),
            .I(N__27356));
    InMux I__5524 (
            .O(N__27382),
            .I(N__27353));
    Span4Mux_v I__5523 (
            .O(N__27379),
            .I(N__27346));
    Span4Mux_s3_v I__5522 (
            .O(N__27374),
            .I(N__27346));
    LocalMux I__5521 (
            .O(N__27371),
            .I(N__27346));
    Odrv12 I__5520 (
            .O(N__27368),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    LocalMux I__5519 (
            .O(N__27365),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    LocalMux I__5518 (
            .O(N__27362),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    Odrv4 I__5517 (
            .O(N__27359),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    Odrv4 I__5516 (
            .O(N__27356),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    LocalMux I__5515 (
            .O(N__27353),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    Odrv4 I__5514 (
            .O(N__27346),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    InMux I__5513 (
            .O(N__27331),
            .I(N__27325));
    InMux I__5512 (
            .O(N__27330),
            .I(N__27325));
    LocalMux I__5511 (
            .O(N__27325),
            .I(\b2v_inst11.N_12 ));
    CascadeMux I__5510 (
            .O(N__27322),
            .I(N__27319));
    InMux I__5509 (
            .O(N__27319),
            .I(N__27308));
    InMux I__5508 (
            .O(N__27318),
            .I(N__27297));
    InMux I__5507 (
            .O(N__27317),
            .I(N__27297));
    InMux I__5506 (
            .O(N__27316),
            .I(N__27289));
    InMux I__5505 (
            .O(N__27315),
            .I(N__27284));
    InMux I__5504 (
            .O(N__27314),
            .I(N__27284));
    InMux I__5503 (
            .O(N__27313),
            .I(N__27279));
    InMux I__5502 (
            .O(N__27312),
            .I(N__27279));
    InMux I__5501 (
            .O(N__27311),
            .I(N__27276));
    LocalMux I__5500 (
            .O(N__27308),
            .I(N__27271));
    InMux I__5499 (
            .O(N__27307),
            .I(N__27266));
    InMux I__5498 (
            .O(N__27306),
            .I(N__27266));
    InMux I__5497 (
            .O(N__27305),
            .I(N__27263));
    InMux I__5496 (
            .O(N__27304),
            .I(N__27259));
    InMux I__5495 (
            .O(N__27303),
            .I(N__27252));
    InMux I__5494 (
            .O(N__27302),
            .I(N__27252));
    LocalMux I__5493 (
            .O(N__27297),
            .I(N__27249));
    InMux I__5492 (
            .O(N__27296),
            .I(N__27240));
    InMux I__5491 (
            .O(N__27295),
            .I(N__27240));
    InMux I__5490 (
            .O(N__27294),
            .I(N__27240));
    InMux I__5489 (
            .O(N__27293),
            .I(N__27240));
    InMux I__5488 (
            .O(N__27292),
            .I(N__27237));
    LocalMux I__5487 (
            .O(N__27289),
            .I(N__27221));
    LocalMux I__5486 (
            .O(N__27284),
            .I(N__27221));
    LocalMux I__5485 (
            .O(N__27279),
            .I(N__27221));
    LocalMux I__5484 (
            .O(N__27276),
            .I(N__27218));
    InMux I__5483 (
            .O(N__27275),
            .I(N__27213));
    InMux I__5482 (
            .O(N__27274),
            .I(N__27213));
    Span4Mux_v I__5481 (
            .O(N__27271),
            .I(N__27206));
    LocalMux I__5480 (
            .O(N__27266),
            .I(N__27206));
    LocalMux I__5479 (
            .O(N__27263),
            .I(N__27206));
    InMux I__5478 (
            .O(N__27262),
            .I(N__27203));
    LocalMux I__5477 (
            .O(N__27259),
            .I(N__27200));
    InMux I__5476 (
            .O(N__27258),
            .I(N__27195));
    InMux I__5475 (
            .O(N__27257),
            .I(N__27195));
    LocalMux I__5474 (
            .O(N__27252),
            .I(N__27188));
    Span4Mux_v I__5473 (
            .O(N__27249),
            .I(N__27188));
    LocalMux I__5472 (
            .O(N__27240),
            .I(N__27188));
    LocalMux I__5471 (
            .O(N__27237),
            .I(N__27185));
    InMux I__5470 (
            .O(N__27236),
            .I(N__27182));
    InMux I__5469 (
            .O(N__27235),
            .I(N__27179));
    InMux I__5468 (
            .O(N__27234),
            .I(N__27168));
    InMux I__5467 (
            .O(N__27233),
            .I(N__27168));
    InMux I__5466 (
            .O(N__27232),
            .I(N__27168));
    InMux I__5465 (
            .O(N__27231),
            .I(N__27168));
    InMux I__5464 (
            .O(N__27230),
            .I(N__27168));
    InMux I__5463 (
            .O(N__27229),
            .I(N__27163));
    InMux I__5462 (
            .O(N__27228),
            .I(N__27163));
    Span4Mux_v I__5461 (
            .O(N__27221),
            .I(N__27160));
    Span4Mux_v I__5460 (
            .O(N__27218),
            .I(N__27153));
    LocalMux I__5459 (
            .O(N__27213),
            .I(N__27153));
    Span4Mux_v I__5458 (
            .O(N__27206),
            .I(N__27153));
    LocalMux I__5457 (
            .O(N__27203),
            .I(N__27148));
    Span4Mux_h I__5456 (
            .O(N__27200),
            .I(N__27148));
    LocalMux I__5455 (
            .O(N__27195),
            .I(N__27141));
    Span4Mux_h I__5454 (
            .O(N__27188),
            .I(N__27141));
    Span4Mux_h I__5453 (
            .O(N__27185),
            .I(N__27141));
    LocalMux I__5452 (
            .O(N__27182),
            .I(\b2v_inst11.func_state_RNINJ641_0Z0Z_1 ));
    LocalMux I__5451 (
            .O(N__27179),
            .I(\b2v_inst11.func_state_RNINJ641_0Z0Z_1 ));
    LocalMux I__5450 (
            .O(N__27168),
            .I(\b2v_inst11.func_state_RNINJ641_0Z0Z_1 ));
    LocalMux I__5449 (
            .O(N__27163),
            .I(\b2v_inst11.func_state_RNINJ641_0Z0Z_1 ));
    Odrv4 I__5448 (
            .O(N__27160),
            .I(\b2v_inst11.func_state_RNINJ641_0Z0Z_1 ));
    Odrv4 I__5447 (
            .O(N__27153),
            .I(\b2v_inst11.func_state_RNINJ641_0Z0Z_1 ));
    Odrv4 I__5446 (
            .O(N__27148),
            .I(\b2v_inst11.func_state_RNINJ641_0Z0Z_1 ));
    Odrv4 I__5445 (
            .O(N__27141),
            .I(\b2v_inst11.func_state_RNINJ641_0Z0Z_1 ));
    InMux I__5444 (
            .O(N__27124),
            .I(N__27121));
    LocalMux I__5443 (
            .O(N__27121),
            .I(N_4));
    InMux I__5442 (
            .O(N__27118),
            .I(N__27115));
    LocalMux I__5441 (
            .O(N__27115),
            .I(N__27112));
    Odrv4 I__5440 (
            .O(N__27112),
            .I(G_26_0_a5_2));
    CascadeMux I__5439 (
            .O(N__27109),
            .I(N__27104));
    InMux I__5438 (
            .O(N__27108),
            .I(N__27098));
    InMux I__5437 (
            .O(N__27107),
            .I(N__27098));
    InMux I__5436 (
            .O(N__27104),
            .I(N__27093));
    InMux I__5435 (
            .O(N__27103),
            .I(N__27093));
    LocalMux I__5434 (
            .O(N__27098),
            .I(N__27084));
    LocalMux I__5433 (
            .O(N__27093),
            .I(N__27081));
    InMux I__5432 (
            .O(N__27092),
            .I(N__27078));
    InMux I__5431 (
            .O(N__27091),
            .I(N__27075));
    CascadeMux I__5430 (
            .O(N__27090),
            .I(N__27072));
    InMux I__5429 (
            .O(N__27089),
            .I(N__27065));
    InMux I__5428 (
            .O(N__27088),
            .I(N__27065));
    InMux I__5427 (
            .O(N__27087),
            .I(N__27062));
    Span4Mux_v I__5426 (
            .O(N__27084),
            .I(N__27053));
    Span4Mux_h I__5425 (
            .O(N__27081),
            .I(N__27053));
    LocalMux I__5424 (
            .O(N__27078),
            .I(N__27053));
    LocalMux I__5423 (
            .O(N__27075),
            .I(N__27053));
    InMux I__5422 (
            .O(N__27072),
            .I(N__27050));
    InMux I__5421 (
            .O(N__27071),
            .I(N__27045));
    InMux I__5420 (
            .O(N__27070),
            .I(N__27045));
    LocalMux I__5419 (
            .O(N__27065),
            .I(curr_state_RNI5VS71_0_1));
    LocalMux I__5418 (
            .O(N__27062),
            .I(curr_state_RNI5VS71_0_1));
    Odrv4 I__5417 (
            .O(N__27053),
            .I(curr_state_RNI5VS71_0_1));
    LocalMux I__5416 (
            .O(N__27050),
            .I(curr_state_RNI5VS71_0_1));
    LocalMux I__5415 (
            .O(N__27045),
            .I(curr_state_RNI5VS71_0_1));
    InMux I__5414 (
            .O(N__27034),
            .I(N__27031));
    LocalMux I__5413 (
            .O(N__27031),
            .I(N__27022));
    InMux I__5412 (
            .O(N__27030),
            .I(N__27016));
    InMux I__5411 (
            .O(N__27029),
            .I(N__27016));
    InMux I__5410 (
            .O(N__27028),
            .I(N__27013));
    InMux I__5409 (
            .O(N__27027),
            .I(N__27008));
    InMux I__5408 (
            .O(N__27026),
            .I(N__27008));
    CascadeMux I__5407 (
            .O(N__27025),
            .I(N__27005));
    Span12Mux_s7_v I__5406 (
            .O(N__27022),
            .I(N__27001));
    InMux I__5405 (
            .O(N__27021),
            .I(N__26998));
    LocalMux I__5404 (
            .O(N__27016),
            .I(N__26995));
    LocalMux I__5403 (
            .O(N__27013),
            .I(N__26990));
    LocalMux I__5402 (
            .O(N__27008),
            .I(N__26990));
    InMux I__5401 (
            .O(N__27005),
            .I(N__26987));
    InMux I__5400 (
            .O(N__27004),
            .I(N__26984));
    Odrv12 I__5399 (
            .O(N__27001),
            .I(RSMRSTn_0));
    LocalMux I__5398 (
            .O(N__26998),
            .I(RSMRSTn_0));
    Odrv4 I__5397 (
            .O(N__26995),
            .I(RSMRSTn_0));
    Odrv12 I__5396 (
            .O(N__26990),
            .I(RSMRSTn_0));
    LocalMux I__5395 (
            .O(N__26987),
            .I(RSMRSTn_0));
    LocalMux I__5394 (
            .O(N__26984),
            .I(RSMRSTn_0));
    CascadeMux I__5393 (
            .O(N__26971),
            .I(\b2v_inst11.N_234_cascade_ ));
    CascadeMux I__5392 (
            .O(N__26968),
            .I(\b2v_inst11.un1_clk_100khz_52_and_i_0_0_cascade_ ));
    CascadeMux I__5391 (
            .O(N__26965),
            .I(N__26961));
    InMux I__5390 (
            .O(N__26964),
            .I(N__26956));
    InMux I__5389 (
            .O(N__26961),
            .I(N__26951));
    InMux I__5388 (
            .O(N__26960),
            .I(N__26946));
    InMux I__5387 (
            .O(N__26959),
            .I(N__26946));
    LocalMux I__5386 (
            .O(N__26956),
            .I(N__26943));
    InMux I__5385 (
            .O(N__26955),
            .I(N__26937));
    InMux I__5384 (
            .O(N__26954),
            .I(N__26937));
    LocalMux I__5383 (
            .O(N__26951),
            .I(N__26934));
    LocalMux I__5382 (
            .O(N__26946),
            .I(N__26931));
    Span4Mux_v I__5381 (
            .O(N__26943),
            .I(N__26928));
    InMux I__5380 (
            .O(N__26942),
            .I(N__26920));
    LocalMux I__5379 (
            .O(N__26937),
            .I(N__26917));
    Span4Mux_v I__5378 (
            .O(N__26934),
            .I(N__26912));
    Span4Mux_v I__5377 (
            .O(N__26931),
            .I(N__26912));
    Span4Mux_h I__5376 (
            .O(N__26928),
            .I(N__26909));
    InMux I__5375 (
            .O(N__26927),
            .I(N__26906));
    InMux I__5374 (
            .O(N__26926),
            .I(N__26899));
    InMux I__5373 (
            .O(N__26925),
            .I(N__26899));
    InMux I__5372 (
            .O(N__26924),
            .I(N__26899));
    InMux I__5371 (
            .O(N__26923),
            .I(N__26896));
    LocalMux I__5370 (
            .O(N__26920),
            .I(SYNTHESIZED_WIRE_47keep_rep1));
    Odrv12 I__5369 (
            .O(N__26917),
            .I(SYNTHESIZED_WIRE_47keep_rep1));
    Odrv4 I__5368 (
            .O(N__26912),
            .I(SYNTHESIZED_WIRE_47keep_rep1));
    Odrv4 I__5367 (
            .O(N__26909),
            .I(SYNTHESIZED_WIRE_47keep_rep1));
    LocalMux I__5366 (
            .O(N__26906),
            .I(SYNTHESIZED_WIRE_47keep_rep1));
    LocalMux I__5365 (
            .O(N__26899),
            .I(SYNTHESIZED_WIRE_47keep_rep1));
    LocalMux I__5364 (
            .O(N__26896),
            .I(SYNTHESIZED_WIRE_47keep_rep1));
    CascadeMux I__5363 (
            .O(N__26881),
            .I(N__26874));
    InMux I__5362 (
            .O(N__26880),
            .I(N__26868));
    InMux I__5361 (
            .O(N__26879),
            .I(N__26868));
    InMux I__5360 (
            .O(N__26878),
            .I(N__26863));
    InMux I__5359 (
            .O(N__26877),
            .I(N__26860));
    InMux I__5358 (
            .O(N__26874),
            .I(N__26855));
    InMux I__5357 (
            .O(N__26873),
            .I(N__26855));
    LocalMux I__5356 (
            .O(N__26868),
            .I(N__26852));
    CascadeMux I__5355 (
            .O(N__26867),
            .I(N__26845));
    InMux I__5354 (
            .O(N__26866),
            .I(N__26840));
    LocalMux I__5353 (
            .O(N__26863),
            .I(N__26837));
    LocalMux I__5352 (
            .O(N__26860),
            .I(N__26834));
    LocalMux I__5351 (
            .O(N__26855),
            .I(N__26831));
    Span4Mux_h I__5350 (
            .O(N__26852),
            .I(N__26828));
    InMux I__5349 (
            .O(N__26851),
            .I(N__26822));
    InMux I__5348 (
            .O(N__26850),
            .I(N__26822));
    InMux I__5347 (
            .O(N__26849),
            .I(N__26811));
    InMux I__5346 (
            .O(N__26848),
            .I(N__26811));
    InMux I__5345 (
            .O(N__26845),
            .I(N__26811));
    InMux I__5344 (
            .O(N__26844),
            .I(N__26811));
    InMux I__5343 (
            .O(N__26843),
            .I(N__26811));
    LocalMux I__5342 (
            .O(N__26840),
            .I(N__26806));
    Span4Mux_v I__5341 (
            .O(N__26837),
            .I(N__26806));
    Span4Mux_v I__5340 (
            .O(N__26834),
            .I(N__26801));
    Span4Mux_h I__5339 (
            .O(N__26831),
            .I(N__26801));
    Span4Mux_h I__5338 (
            .O(N__26828),
            .I(N__26798));
    InMux I__5337 (
            .O(N__26827),
            .I(N__26795));
    LocalMux I__5336 (
            .O(N__26822),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    LocalMux I__5335 (
            .O(N__26811),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    Odrv4 I__5334 (
            .O(N__26806),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    Odrv4 I__5333 (
            .O(N__26801),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    Odrv4 I__5332 (
            .O(N__26798),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    LocalMux I__5331 (
            .O(N__26795),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    CascadeMux I__5330 (
            .O(N__26782),
            .I(N__26776));
    CascadeMux I__5329 (
            .O(N__26781),
            .I(N__26773));
    InMux I__5328 (
            .O(N__26780),
            .I(N__26770));
    CascadeMux I__5327 (
            .O(N__26779),
            .I(N__26767));
    InMux I__5326 (
            .O(N__26776),
            .I(N__26761));
    InMux I__5325 (
            .O(N__26773),
            .I(N__26758));
    LocalMux I__5324 (
            .O(N__26770),
            .I(N__26754));
    InMux I__5323 (
            .O(N__26767),
            .I(N__26749));
    InMux I__5322 (
            .O(N__26766),
            .I(N__26749));
    InMux I__5321 (
            .O(N__26765),
            .I(N__26746));
    CascadeMux I__5320 (
            .O(N__26764),
            .I(N__26743));
    LocalMux I__5319 (
            .O(N__26761),
            .I(N__26739));
    LocalMux I__5318 (
            .O(N__26758),
            .I(N__26736));
    CascadeMux I__5317 (
            .O(N__26757),
            .I(N__26733));
    Span4Mux_h I__5316 (
            .O(N__26754),
            .I(N__26729));
    LocalMux I__5315 (
            .O(N__26749),
            .I(N__26724));
    LocalMux I__5314 (
            .O(N__26746),
            .I(N__26724));
    InMux I__5313 (
            .O(N__26743),
            .I(N__26721));
    InMux I__5312 (
            .O(N__26742),
            .I(N__26718));
    Span4Mux_v I__5311 (
            .O(N__26739),
            .I(N__26713));
    Span4Mux_v I__5310 (
            .O(N__26736),
            .I(N__26713));
    InMux I__5309 (
            .O(N__26733),
            .I(N__26708));
    InMux I__5308 (
            .O(N__26732),
            .I(N__26708));
    Span4Mux_v I__5307 (
            .O(N__26729),
            .I(N__26703));
    Span4Mux_h I__5306 (
            .O(N__26724),
            .I(N__26703));
    LocalMux I__5305 (
            .O(N__26721),
            .I(dutycycle_RNIIOE3D_0_5));
    LocalMux I__5304 (
            .O(N__26718),
            .I(dutycycle_RNIIOE3D_0_5));
    Odrv4 I__5303 (
            .O(N__26713),
            .I(dutycycle_RNIIOE3D_0_5));
    LocalMux I__5302 (
            .O(N__26708),
            .I(dutycycle_RNIIOE3D_0_5));
    Odrv4 I__5301 (
            .O(N__26703),
            .I(dutycycle_RNIIOE3D_0_5));
    InMux I__5300 (
            .O(N__26692),
            .I(bfn_9_10_0_));
    CascadeMux I__5299 (
            .O(N__26689),
            .I(N__26686));
    InMux I__5298 (
            .O(N__26686),
            .I(N__26683));
    LocalMux I__5297 (
            .O(N__26683),
            .I(\b2v_inst20.un4_counter_1_and ));
    InMux I__5296 (
            .O(N__26680),
            .I(N__26677));
    LocalMux I__5295 (
            .O(N__26677),
            .I(N__26674));
    Span4Mux_v I__5294 (
            .O(N__26674),
            .I(N__26671));
    Odrv4 I__5293 (
            .O(N__26671),
            .I(\b2v_inst11.dutycycle_RNITBKN1Z0Z_7 ));
    InMux I__5292 (
            .O(N__26668),
            .I(N__26664));
    InMux I__5291 (
            .O(N__26667),
            .I(N__26661));
    LocalMux I__5290 (
            .O(N__26664),
            .I(N_229));
    LocalMux I__5289 (
            .O(N__26661),
            .I(N_229));
    CascadeMux I__5288 (
            .O(N__26656),
            .I(\b2v_inst5.count_enZ0_cascade_ ));
    CascadeMux I__5287 (
            .O(N__26653),
            .I(N__26650));
    InMux I__5286 (
            .O(N__26650),
            .I(N__26646));
    CascadeMux I__5285 (
            .O(N__26649),
            .I(N__26643));
    LocalMux I__5284 (
            .O(N__26646),
            .I(N__26639));
    InMux I__5283 (
            .O(N__26643),
            .I(N__26633));
    InMux I__5282 (
            .O(N__26642),
            .I(N__26633));
    Span4Mux_h I__5281 (
            .O(N__26639),
            .I(N__26630));
    InMux I__5280 (
            .O(N__26638),
            .I(N__26627));
    LocalMux I__5279 (
            .O(N__26633),
            .I(\b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    Odrv4 I__5278 (
            .O(N__26630),
            .I(\b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    LocalMux I__5277 (
            .O(N__26627),
            .I(\b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    InMux I__5276 (
            .O(N__26620),
            .I(N__26617));
    LocalMux I__5275 (
            .O(N__26617),
            .I(N__26614));
    Odrv4 I__5274 (
            .O(N__26614),
            .I(\b2v_inst11.g0_2_1 ));
    InMux I__5273 (
            .O(N__26611),
            .I(N__26607));
    InMux I__5272 (
            .O(N__26610),
            .I(N__26603));
    LocalMux I__5271 (
            .O(N__26607),
            .I(N__26600));
    InMux I__5270 (
            .O(N__26606),
            .I(N__26597));
    LocalMux I__5269 (
            .O(N__26603),
            .I(N__26594));
    Odrv4 I__5268 (
            .O(N__26600),
            .I(\b2v_inst11.pwm_outZ0 ));
    LocalMux I__5267 (
            .O(N__26597),
            .I(\b2v_inst11.pwm_outZ0 ));
    Odrv4 I__5266 (
            .O(N__26594),
            .I(\b2v_inst11.pwm_outZ0 ));
    SRMux I__5265 (
            .O(N__26587),
            .I(N__26584));
    LocalMux I__5264 (
            .O(N__26584),
            .I(N__26581));
    Span4Mux_v I__5263 (
            .O(N__26581),
            .I(N__26578));
    Odrv4 I__5262 (
            .O(N__26578),
            .I(\b2v_inst11.pwm_out_1_sqmuxa ));
    CascadeMux I__5261 (
            .O(N__26575),
            .I(N__26572));
    InMux I__5260 (
            .O(N__26572),
            .I(N__26569));
    LocalMux I__5259 (
            .O(N__26569),
            .I(\b2v_inst20.un4_counter_0_and ));
    CascadeMux I__5258 (
            .O(N__26566),
            .I(\b2v_inst11.count_RNIZ0Z_1_cascade_ ));
    InMux I__5257 (
            .O(N__26563),
            .I(N__26560));
    LocalMux I__5256 (
            .O(N__26560),
            .I(N__26556));
    CascadeMux I__5255 (
            .O(N__26559),
            .I(N__26552));
    Span12Mux_s8_h I__5254 (
            .O(N__26556),
            .I(N__26549));
    InMux I__5253 (
            .O(N__26555),
            .I(N__26546));
    InMux I__5252 (
            .O(N__26552),
            .I(N__26543));
    Odrv12 I__5251 (
            .O(N__26549),
            .I(\b2v_inst11.countZ0Z_1 ));
    LocalMux I__5250 (
            .O(N__26546),
            .I(\b2v_inst11.countZ0Z_1 ));
    LocalMux I__5249 (
            .O(N__26543),
            .I(\b2v_inst11.countZ0Z_1 ));
    InMux I__5248 (
            .O(N__26536),
            .I(N__26532));
    InMux I__5247 (
            .O(N__26535),
            .I(N__26528));
    LocalMux I__5246 (
            .O(N__26532),
            .I(N__26525));
    InMux I__5245 (
            .O(N__26531),
            .I(N__26522));
    LocalMux I__5244 (
            .O(N__26528),
            .I(N__26519));
    Span4Mux_v I__5243 (
            .O(N__26525),
            .I(N__26512));
    LocalMux I__5242 (
            .O(N__26522),
            .I(N__26512));
    Span4Mux_h I__5241 (
            .O(N__26519),
            .I(N__26509));
    InMux I__5240 (
            .O(N__26518),
            .I(N__26506));
    InMux I__5239 (
            .O(N__26517),
            .I(N__26503));
    Odrv4 I__5238 (
            .O(N__26512),
            .I(\b2v_inst11.countZ0Z_0 ));
    Odrv4 I__5237 (
            .O(N__26509),
            .I(\b2v_inst11.countZ0Z_0 ));
    LocalMux I__5236 (
            .O(N__26506),
            .I(\b2v_inst11.countZ0Z_0 ));
    LocalMux I__5235 (
            .O(N__26503),
            .I(\b2v_inst11.countZ0Z_0 ));
    CascadeMux I__5234 (
            .O(N__26494),
            .I(\b2v_inst11.countZ0Z_1_cascade_ ));
    InMux I__5233 (
            .O(N__26491),
            .I(N__26470));
    InMux I__5232 (
            .O(N__26490),
            .I(N__26470));
    InMux I__5231 (
            .O(N__26489),
            .I(N__26470));
    InMux I__5230 (
            .O(N__26488),
            .I(N__26470));
    InMux I__5229 (
            .O(N__26487),
            .I(N__26465));
    InMux I__5228 (
            .O(N__26486),
            .I(N__26465));
    InMux I__5227 (
            .O(N__26485),
            .I(N__26455));
    InMux I__5226 (
            .O(N__26484),
            .I(N__26455));
    InMux I__5225 (
            .O(N__26483),
            .I(N__26455));
    InMux I__5224 (
            .O(N__26482),
            .I(N__26446));
    InMux I__5223 (
            .O(N__26481),
            .I(N__26446));
    InMux I__5222 (
            .O(N__26480),
            .I(N__26446));
    InMux I__5221 (
            .O(N__26479),
            .I(N__26446));
    LocalMux I__5220 (
            .O(N__26470),
            .I(N__26441));
    LocalMux I__5219 (
            .O(N__26465),
            .I(N__26441));
    InMux I__5218 (
            .O(N__26464),
            .I(N__26433));
    InMux I__5217 (
            .O(N__26463),
            .I(N__26433));
    InMux I__5216 (
            .O(N__26462),
            .I(N__26433));
    LocalMux I__5215 (
            .O(N__26455),
            .I(N__26428));
    LocalMux I__5214 (
            .O(N__26446),
            .I(N__26428));
    Span4Mux_h I__5213 (
            .O(N__26441),
            .I(N__26425));
    InMux I__5212 (
            .O(N__26440),
            .I(N__26422));
    LocalMux I__5211 (
            .O(N__26433),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    Odrv4 I__5210 (
            .O(N__26428),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    Odrv4 I__5209 (
            .O(N__26425),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    LocalMux I__5208 (
            .O(N__26422),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    InMux I__5207 (
            .O(N__26413),
            .I(N__26410));
    LocalMux I__5206 (
            .O(N__26410),
            .I(\b2v_inst11.count_0_1 ));
    InMux I__5205 (
            .O(N__26407),
            .I(N__26404));
    LocalMux I__5204 (
            .O(N__26404),
            .I(N__26400));
    InMux I__5203 (
            .O(N__26403),
            .I(N__26397));
    Span4Mux_h I__5202 (
            .O(N__26400),
            .I(N__26393));
    LocalMux I__5201 (
            .O(N__26397),
            .I(N__26390));
    InMux I__5200 (
            .O(N__26396),
            .I(N__26387));
    Odrv4 I__5199 (
            .O(N__26393),
            .I(\b2v_inst11.countZ0Z_8 ));
    Odrv4 I__5198 (
            .O(N__26390),
            .I(\b2v_inst11.countZ0Z_8 ));
    LocalMux I__5197 (
            .O(N__26387),
            .I(\b2v_inst11.countZ0Z_8 ));
    InMux I__5196 (
            .O(N__26380),
            .I(N__26374));
    InMux I__5195 (
            .O(N__26379),
            .I(N__26374));
    LocalMux I__5194 (
            .O(N__26374),
            .I(\b2v_inst11.un1_count_cry_7_c_RNIOU0EZ0 ));
    InMux I__5193 (
            .O(N__26371),
            .I(N__26368));
    LocalMux I__5192 (
            .O(N__26368),
            .I(\b2v_inst11.count_0_8 ));
    CascadeMux I__5191 (
            .O(N__26365),
            .I(N__26361));
    InMux I__5190 (
            .O(N__26364),
            .I(N__26358));
    InMux I__5189 (
            .O(N__26361),
            .I(N__26355));
    LocalMux I__5188 (
            .O(N__26358),
            .I(N__26351));
    LocalMux I__5187 (
            .O(N__26355),
            .I(N__26348));
    CascadeMux I__5186 (
            .O(N__26354),
            .I(N__26345));
    Span4Mux_h I__5185 (
            .O(N__26351),
            .I(N__26342));
    Span4Mux_s3_h I__5184 (
            .O(N__26348),
            .I(N__26339));
    InMux I__5183 (
            .O(N__26345),
            .I(N__26336));
    Odrv4 I__5182 (
            .O(N__26342),
            .I(\b2v_inst11.countZ0Z_9 ));
    Odrv4 I__5181 (
            .O(N__26339),
            .I(\b2v_inst11.countZ0Z_9 ));
    LocalMux I__5180 (
            .O(N__26336),
            .I(\b2v_inst11.countZ0Z_9 ));
    InMux I__5179 (
            .O(N__26329),
            .I(N__26323));
    InMux I__5178 (
            .O(N__26328),
            .I(N__26323));
    LocalMux I__5177 (
            .O(N__26323),
            .I(\b2v_inst11.un1_count_cry_8_c_RNIP02EZ0 ));
    InMux I__5176 (
            .O(N__26320),
            .I(N__26317));
    LocalMux I__5175 (
            .O(N__26317),
            .I(\b2v_inst11.count_0_9 ));
    InMux I__5174 (
            .O(N__26314),
            .I(N__26311));
    LocalMux I__5173 (
            .O(N__26311),
            .I(\b2v_inst5.curr_state_3_0 ));
    CascadeMux I__5172 (
            .O(N__26308),
            .I(N__26302));
    InMux I__5171 (
            .O(N__26307),
            .I(N__26298));
    InMux I__5170 (
            .O(N__26306),
            .I(N__26289));
    InMux I__5169 (
            .O(N__26305),
            .I(N__26289));
    InMux I__5168 (
            .O(N__26302),
            .I(N__26289));
    InMux I__5167 (
            .O(N__26301),
            .I(N__26289));
    LocalMux I__5166 (
            .O(N__26298),
            .I(\b2v_inst5.curr_stateZ0Z_0 ));
    LocalMux I__5165 (
            .O(N__26289),
            .I(\b2v_inst5.curr_stateZ0Z_0 ));
    InMux I__5164 (
            .O(N__26284),
            .I(N__26279));
    InMux I__5163 (
            .O(N__26283),
            .I(N__26274));
    InMux I__5162 (
            .O(N__26282),
            .I(N__26274));
    LocalMux I__5161 (
            .O(N__26279),
            .I(G_2727));
    LocalMux I__5160 (
            .O(N__26274),
            .I(G_2727));
    CascadeMux I__5159 (
            .O(N__26269),
            .I(\b2v_inst5.curr_stateZ0Z_0_cascade_ ));
    InMux I__5158 (
            .O(N__26266),
            .I(N__26263));
    LocalMux I__5157 (
            .O(N__26263),
            .I(\b2v_inst5.m4_0 ));
    InMux I__5156 (
            .O(N__26260),
            .I(N__26257));
    LocalMux I__5155 (
            .O(N__26257),
            .I(N__26254));
    Span4Mux_h I__5154 (
            .O(N__26254),
            .I(N__26250));
    InMux I__5153 (
            .O(N__26253),
            .I(N__26247));
    Span4Mux_v I__5152 (
            .O(N__26250),
            .I(N__26244));
    LocalMux I__5151 (
            .O(N__26247),
            .I(N__26241));
    Odrv4 I__5150 (
            .O(N__26244),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1 ));
    Odrv12 I__5149 (
            .O(N__26241),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1 ));
    InMux I__5148 (
            .O(N__26236),
            .I(N__26225));
    InMux I__5147 (
            .O(N__26235),
            .I(N__26225));
    InMux I__5146 (
            .O(N__26234),
            .I(N__26220));
    InMux I__5145 (
            .O(N__26233),
            .I(N__26216));
    InMux I__5144 (
            .O(N__26232),
            .I(N__26207));
    CascadeMux I__5143 (
            .O(N__26231),
            .I(N__26204));
    CascadeMux I__5142 (
            .O(N__26230),
            .I(N__26200));
    LocalMux I__5141 (
            .O(N__26225),
            .I(N__26196));
    CascadeMux I__5140 (
            .O(N__26224),
            .I(N__26193));
    InMux I__5139 (
            .O(N__26223),
            .I(N__26190));
    LocalMux I__5138 (
            .O(N__26220),
            .I(N__26184));
    InMux I__5137 (
            .O(N__26219),
            .I(N__26181));
    LocalMux I__5136 (
            .O(N__26216),
            .I(N__26175));
    InMux I__5135 (
            .O(N__26215),
            .I(N__26168));
    InMux I__5134 (
            .O(N__26214),
            .I(N__26168));
    InMux I__5133 (
            .O(N__26213),
            .I(N__26168));
    InMux I__5132 (
            .O(N__26212),
            .I(N__26163));
    InMux I__5131 (
            .O(N__26211),
            .I(N__26163));
    InMux I__5130 (
            .O(N__26210),
            .I(N__26160));
    LocalMux I__5129 (
            .O(N__26207),
            .I(N__26157));
    InMux I__5128 (
            .O(N__26204),
            .I(N__26148));
    InMux I__5127 (
            .O(N__26203),
            .I(N__26148));
    InMux I__5126 (
            .O(N__26200),
            .I(N__26148));
    InMux I__5125 (
            .O(N__26199),
            .I(N__26148));
    Span4Mux_v I__5124 (
            .O(N__26196),
            .I(N__26145));
    InMux I__5123 (
            .O(N__26193),
            .I(N__26142));
    LocalMux I__5122 (
            .O(N__26190),
            .I(N__26139));
    InMux I__5121 (
            .O(N__26189),
            .I(N__26134));
    InMux I__5120 (
            .O(N__26188),
            .I(N__26134));
    InMux I__5119 (
            .O(N__26187),
            .I(N__26131));
    Span4Mux_h I__5118 (
            .O(N__26184),
            .I(N__26126));
    LocalMux I__5117 (
            .O(N__26181),
            .I(N__26126));
    InMux I__5116 (
            .O(N__26180),
            .I(N__26119));
    InMux I__5115 (
            .O(N__26179),
            .I(N__26119));
    InMux I__5114 (
            .O(N__26178),
            .I(N__26119));
    Span4Mux_h I__5113 (
            .O(N__26175),
            .I(N__26112));
    LocalMux I__5112 (
            .O(N__26168),
            .I(N__26112));
    LocalMux I__5111 (
            .O(N__26163),
            .I(N__26112));
    LocalMux I__5110 (
            .O(N__26160),
            .I(N__26105));
    Span4Mux_v I__5109 (
            .O(N__26157),
            .I(N__26105));
    LocalMux I__5108 (
            .O(N__26148),
            .I(N__26105));
    Odrv4 I__5107 (
            .O(N__26145),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    LocalMux I__5106 (
            .O(N__26142),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    Odrv12 I__5105 (
            .O(N__26139),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    LocalMux I__5104 (
            .O(N__26134),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    LocalMux I__5103 (
            .O(N__26131),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    Odrv4 I__5102 (
            .O(N__26126),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    LocalMux I__5101 (
            .O(N__26119),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    Odrv4 I__5100 (
            .O(N__26112),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    Odrv4 I__5099 (
            .O(N__26105),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    InMux I__5098 (
            .O(N__26086),
            .I(N__26080));
    InMux I__5097 (
            .O(N__26085),
            .I(N__26080));
    LocalMux I__5096 (
            .O(N__26080),
            .I(\b2v_inst11.un1_count_cry_2_c_RNIJKRDZ0 ));
    InMux I__5095 (
            .O(N__26077),
            .I(N__26074));
    LocalMux I__5094 (
            .O(N__26074),
            .I(\b2v_inst11.count_0_3 ));
    InMux I__5093 (
            .O(N__26071),
            .I(N__26067));
    CascadeMux I__5092 (
            .O(N__26070),
            .I(N__26063));
    LocalMux I__5091 (
            .O(N__26067),
            .I(N__26060));
    InMux I__5090 (
            .O(N__26066),
            .I(N__26057));
    InMux I__5089 (
            .O(N__26063),
            .I(N__26054));
    Odrv4 I__5088 (
            .O(N__26060),
            .I(\b2v_inst11.countZ0Z_13 ));
    LocalMux I__5087 (
            .O(N__26057),
            .I(\b2v_inst11.countZ0Z_13 ));
    LocalMux I__5086 (
            .O(N__26054),
            .I(\b2v_inst11.countZ0Z_13 ));
    CascadeMux I__5085 (
            .O(N__26047),
            .I(N__26044));
    InMux I__5084 (
            .O(N__26044),
            .I(N__26038));
    InMux I__5083 (
            .O(N__26043),
            .I(N__26038));
    LocalMux I__5082 (
            .O(N__26038),
            .I(\b2v_inst11.un1_count_cry_12_c_RNI48TZ0Z6 ));
    InMux I__5081 (
            .O(N__26035),
            .I(N__26032));
    LocalMux I__5080 (
            .O(N__26032),
            .I(\b2v_inst11.count_0_13 ));
    InMux I__5079 (
            .O(N__26029),
            .I(N__26026));
    LocalMux I__5078 (
            .O(N__26026),
            .I(N__26022));
    CascadeMux I__5077 (
            .O(N__26025),
            .I(N__26018));
    Span4Mux_v I__5076 (
            .O(N__26022),
            .I(N__26015));
    InMux I__5075 (
            .O(N__26021),
            .I(N__26012));
    InMux I__5074 (
            .O(N__26018),
            .I(N__26009));
    Odrv4 I__5073 (
            .O(N__26015),
            .I(\b2v_inst11.countZ0Z_4 ));
    LocalMux I__5072 (
            .O(N__26012),
            .I(\b2v_inst11.countZ0Z_4 ));
    LocalMux I__5071 (
            .O(N__26009),
            .I(\b2v_inst11.countZ0Z_4 ));
    InMux I__5070 (
            .O(N__26002),
            .I(N__25996));
    InMux I__5069 (
            .O(N__26001),
            .I(N__25996));
    LocalMux I__5068 (
            .O(N__25996),
            .I(\b2v_inst11.un1_count_cry_3_c_RNIKMSDZ0 ));
    InMux I__5067 (
            .O(N__25993),
            .I(N__25990));
    LocalMux I__5066 (
            .O(N__25990),
            .I(\b2v_inst11.count_0_4 ));
    InMux I__5065 (
            .O(N__25987),
            .I(N__25984));
    LocalMux I__5064 (
            .O(N__25984),
            .I(N__25980));
    CascadeMux I__5063 (
            .O(N__25983),
            .I(N__25976));
    Span4Mux_v I__5062 (
            .O(N__25980),
            .I(N__25973));
    InMux I__5061 (
            .O(N__25979),
            .I(N__25970));
    InMux I__5060 (
            .O(N__25976),
            .I(N__25967));
    Odrv4 I__5059 (
            .O(N__25973),
            .I(\b2v_inst11.countZ0Z_5 ));
    LocalMux I__5058 (
            .O(N__25970),
            .I(\b2v_inst11.countZ0Z_5 ));
    LocalMux I__5057 (
            .O(N__25967),
            .I(\b2v_inst11.countZ0Z_5 ));
    InMux I__5056 (
            .O(N__25960),
            .I(N__25954));
    InMux I__5055 (
            .O(N__25959),
            .I(N__25954));
    LocalMux I__5054 (
            .O(N__25954),
            .I(\b2v_inst11.un1_count_cry_4_c_RNILOTDZ0 ));
    InMux I__5053 (
            .O(N__25951),
            .I(N__25948));
    LocalMux I__5052 (
            .O(N__25948),
            .I(\b2v_inst11.count_0_5 ));
    InMux I__5051 (
            .O(N__25945),
            .I(N__25942));
    LocalMux I__5050 (
            .O(N__25942),
            .I(N__25939));
    Span4Mux_v I__5049 (
            .O(N__25939),
            .I(N__25936));
    Odrv4 I__5048 (
            .O(N__25936),
            .I(\b2v_inst11.count_0_0 ));
    InMux I__5047 (
            .O(N__25933),
            .I(N__25930));
    LocalMux I__5046 (
            .O(N__25930),
            .I(N__25927));
    Odrv4 I__5045 (
            .O(N__25927),
            .I(\b2v_inst11.count_RNI_2_0 ));
    CascadeMux I__5044 (
            .O(N__25924),
            .I(\b2v_inst11.countZ0Z_0_cascade_ ));
    CascadeMux I__5043 (
            .O(N__25921),
            .I(N__25916));
    InMux I__5042 (
            .O(N__25920),
            .I(N__25913));
    InMux I__5041 (
            .O(N__25919),
            .I(N__25910));
    InMux I__5040 (
            .O(N__25916),
            .I(N__25907));
    LocalMux I__5039 (
            .O(N__25913),
            .I(N__25904));
    LocalMux I__5038 (
            .O(N__25910),
            .I(N__25899));
    LocalMux I__5037 (
            .O(N__25907),
            .I(N__25899));
    Odrv4 I__5036 (
            .O(N__25904),
            .I(\b2v_inst11.countZ0Z_2 ));
    Odrv4 I__5035 (
            .O(N__25899),
            .I(\b2v_inst11.countZ0Z_2 ));
    InMux I__5034 (
            .O(N__25894),
            .I(N__25890));
    CascadeMux I__5033 (
            .O(N__25893),
            .I(N__25886));
    LocalMux I__5032 (
            .O(N__25890),
            .I(N__25883));
    InMux I__5031 (
            .O(N__25889),
            .I(N__25880));
    InMux I__5030 (
            .O(N__25886),
            .I(N__25877));
    Odrv4 I__5029 (
            .O(N__25883),
            .I(\b2v_inst11.countZ0Z_7 ));
    LocalMux I__5028 (
            .O(N__25880),
            .I(\b2v_inst11.countZ0Z_7 ));
    LocalMux I__5027 (
            .O(N__25877),
            .I(\b2v_inst11.countZ0Z_7 ));
    InMux I__5026 (
            .O(N__25870),
            .I(N__25867));
    LocalMux I__5025 (
            .O(N__25867),
            .I(N__25863));
    InMux I__5024 (
            .O(N__25866),
            .I(N__25859));
    Span12Mux_s11_v I__5023 (
            .O(N__25863),
            .I(N__25856));
    InMux I__5022 (
            .O(N__25862),
            .I(N__25853));
    LocalMux I__5021 (
            .O(N__25859),
            .I(\b2v_inst11.countZ0Z_15 ));
    Odrv12 I__5020 (
            .O(N__25856),
            .I(\b2v_inst11.countZ0Z_15 ));
    LocalMux I__5019 (
            .O(N__25853),
            .I(\b2v_inst11.countZ0Z_15 ));
    InMux I__5018 (
            .O(N__25846),
            .I(N__25843));
    LocalMux I__5017 (
            .O(N__25843),
            .I(N__25839));
    InMux I__5016 (
            .O(N__25842),
            .I(N__25836));
    Span4Mux_v I__5015 (
            .O(N__25839),
            .I(N__25832));
    LocalMux I__5014 (
            .O(N__25836),
            .I(N__25829));
    InMux I__5013 (
            .O(N__25835),
            .I(N__25826));
    Odrv4 I__5012 (
            .O(N__25832),
            .I(\b2v_inst11.countZ0Z_11 ));
    Odrv4 I__5011 (
            .O(N__25829),
            .I(\b2v_inst11.countZ0Z_11 ));
    LocalMux I__5010 (
            .O(N__25826),
            .I(\b2v_inst11.countZ0Z_11 ));
    InMux I__5009 (
            .O(N__25819),
            .I(N__25816));
    LocalMux I__5008 (
            .O(N__25816),
            .I(N__25811));
    InMux I__5007 (
            .O(N__25815),
            .I(N__25808));
    CascadeMux I__5006 (
            .O(N__25814),
            .I(N__25805));
    Span4Mux_v I__5005 (
            .O(N__25811),
            .I(N__25802));
    LocalMux I__5004 (
            .O(N__25808),
            .I(N__25799));
    InMux I__5003 (
            .O(N__25805),
            .I(N__25796));
    Odrv4 I__5002 (
            .O(N__25802),
            .I(\b2v_inst11.countZ0Z_10 ));
    Odrv4 I__5001 (
            .O(N__25799),
            .I(\b2v_inst11.countZ0Z_10 ));
    LocalMux I__5000 (
            .O(N__25796),
            .I(\b2v_inst11.countZ0Z_10 ));
    InMux I__4999 (
            .O(N__25789),
            .I(N__25784));
    CascadeMux I__4998 (
            .O(N__25788),
            .I(N__25781));
    InMux I__4997 (
            .O(N__25787),
            .I(N__25778));
    LocalMux I__4996 (
            .O(N__25784),
            .I(N__25775));
    InMux I__4995 (
            .O(N__25781),
            .I(N__25772));
    LocalMux I__4994 (
            .O(N__25778),
            .I(\b2v_inst11.countZ0Z_12 ));
    Odrv4 I__4993 (
            .O(N__25775),
            .I(\b2v_inst11.countZ0Z_12 ));
    LocalMux I__4992 (
            .O(N__25772),
            .I(\b2v_inst11.countZ0Z_12 ));
    InMux I__4991 (
            .O(N__25765),
            .I(N__25762));
    LocalMux I__4990 (
            .O(N__25762),
            .I(\b2v_inst11.un79_clk_100khzlt6 ));
    CascadeMux I__4989 (
            .O(N__25759),
            .I(N__25754));
    InMux I__4988 (
            .O(N__25758),
            .I(N__25751));
    InMux I__4987 (
            .O(N__25757),
            .I(N__25748));
    InMux I__4986 (
            .O(N__25754),
            .I(N__25745));
    LocalMux I__4985 (
            .O(N__25751),
            .I(\b2v_inst11.countZ0Z_6 ));
    LocalMux I__4984 (
            .O(N__25748),
            .I(\b2v_inst11.countZ0Z_6 ));
    LocalMux I__4983 (
            .O(N__25745),
            .I(\b2v_inst11.countZ0Z_6 ));
    CascadeMux I__4982 (
            .O(N__25738),
            .I(\b2v_inst11.un79_clk_100khzlto15_5_cascade_ ));
    CascadeMux I__4981 (
            .O(N__25735),
            .I(N__25732));
    InMux I__4980 (
            .O(N__25732),
            .I(N__25727));
    InMux I__4979 (
            .O(N__25731),
            .I(N__25724));
    InMux I__4978 (
            .O(N__25730),
            .I(N__25721));
    LocalMux I__4977 (
            .O(N__25727),
            .I(N__25718));
    LocalMux I__4976 (
            .O(N__25724),
            .I(\b2v_inst11.countZ0Z_14 ));
    LocalMux I__4975 (
            .O(N__25721),
            .I(\b2v_inst11.countZ0Z_14 ));
    Odrv4 I__4974 (
            .O(N__25718),
            .I(\b2v_inst11.countZ0Z_14 ));
    CascadeMux I__4973 (
            .O(N__25711),
            .I(\b2v_inst11.un79_clk_100khzlto15_7_cascade_ ));
    InMux I__4972 (
            .O(N__25708),
            .I(N__25705));
    LocalMux I__4971 (
            .O(N__25705),
            .I(\b2v_inst11.un79_clk_100khzlto15_4 ));
    CascadeMux I__4970 (
            .O(N__25702),
            .I(N__25697));
    InMux I__4969 (
            .O(N__25701),
            .I(N__25693));
    InMux I__4968 (
            .O(N__25700),
            .I(N__25686));
    InMux I__4967 (
            .O(N__25697),
            .I(N__25686));
    InMux I__4966 (
            .O(N__25696),
            .I(N__25686));
    LocalMux I__4965 (
            .O(N__25693),
            .I(N__25683));
    LocalMux I__4964 (
            .O(N__25686),
            .I(N__25680));
    Span4Mux_v I__4963 (
            .O(N__25683),
            .I(N__25676));
    Span4Mux_h I__4962 (
            .O(N__25680),
            .I(N__25673));
    InMux I__4961 (
            .O(N__25679),
            .I(N__25670));
    Odrv4 I__4960 (
            .O(N__25676),
            .I(\b2v_inst11.count_RNIZ0Z_13 ));
    Odrv4 I__4959 (
            .O(N__25673),
            .I(\b2v_inst11.count_RNIZ0Z_13 ));
    LocalMux I__4958 (
            .O(N__25670),
            .I(\b2v_inst11.count_RNIZ0Z_13 ));
    InMux I__4957 (
            .O(N__25663),
            .I(N__25657));
    InMux I__4956 (
            .O(N__25662),
            .I(N__25657));
    LocalMux I__4955 (
            .O(N__25657),
            .I(N__25649));
    InMux I__4954 (
            .O(N__25656),
            .I(N__25646));
    InMux I__4953 (
            .O(N__25655),
            .I(N__25637));
    InMux I__4952 (
            .O(N__25654),
            .I(N__25637));
    InMux I__4951 (
            .O(N__25653),
            .I(N__25637));
    InMux I__4950 (
            .O(N__25652),
            .I(N__25637));
    Span4Mux_v I__4949 (
            .O(N__25649),
            .I(N__25634));
    LocalMux I__4948 (
            .O(N__25646),
            .I(\b2v_inst11.curr_stateZ0Z_0 ));
    LocalMux I__4947 (
            .O(N__25637),
            .I(\b2v_inst11.curr_stateZ0Z_0 ));
    Odrv4 I__4946 (
            .O(N__25634),
            .I(\b2v_inst11.curr_stateZ0Z_0 ));
    CascadeMux I__4945 (
            .O(N__25627),
            .I(\b2v_inst11.count_RNIZ0Z_13_cascade_ ));
    InMux I__4944 (
            .O(N__25624),
            .I(N__25621));
    LocalMux I__4943 (
            .O(N__25621),
            .I(N__25617));
    CascadeMux I__4942 (
            .O(N__25620),
            .I(N__25613));
    Span4Mux_v I__4941 (
            .O(N__25617),
            .I(N__25610));
    InMux I__4940 (
            .O(N__25616),
            .I(N__25607));
    InMux I__4939 (
            .O(N__25613),
            .I(N__25604));
    Odrv4 I__4938 (
            .O(N__25610),
            .I(\b2v_inst11.countZ0Z_3 ));
    LocalMux I__4937 (
            .O(N__25607),
            .I(\b2v_inst11.countZ0Z_3 ));
    LocalMux I__4936 (
            .O(N__25604),
            .I(\b2v_inst11.countZ0Z_3 ));
    CascadeMux I__4935 (
            .O(N__25597),
            .I(N__25591));
    CascadeMux I__4934 (
            .O(N__25596),
            .I(N__25586));
    InMux I__4933 (
            .O(N__25595),
            .I(N__25583));
    InMux I__4932 (
            .O(N__25594),
            .I(N__25578));
    InMux I__4931 (
            .O(N__25591),
            .I(N__25578));
    InMux I__4930 (
            .O(N__25590),
            .I(N__25575));
    InMux I__4929 (
            .O(N__25589),
            .I(N__25572));
    InMux I__4928 (
            .O(N__25586),
            .I(N__25567));
    LocalMux I__4927 (
            .O(N__25583),
            .I(N__25562));
    LocalMux I__4926 (
            .O(N__25578),
            .I(N__25562));
    LocalMux I__4925 (
            .O(N__25575),
            .I(N__25559));
    LocalMux I__4924 (
            .O(N__25572),
            .I(N__25556));
    InMux I__4923 (
            .O(N__25571),
            .I(N__25553));
    CascadeMux I__4922 (
            .O(N__25570),
            .I(N__25545));
    LocalMux I__4921 (
            .O(N__25567),
            .I(N__25540));
    Span4Mux_h I__4920 (
            .O(N__25562),
            .I(N__25540));
    Span12Mux_s5_h I__4919 (
            .O(N__25559),
            .I(N__25537));
    Span4Mux_v I__4918 (
            .O(N__25556),
            .I(N__25534));
    LocalMux I__4917 (
            .O(N__25553),
            .I(N__25531));
    InMux I__4916 (
            .O(N__25552),
            .I(N__25528));
    InMux I__4915 (
            .O(N__25551),
            .I(N__25525));
    InMux I__4914 (
            .O(N__25550),
            .I(N__25520));
    InMux I__4913 (
            .O(N__25549),
            .I(N__25520));
    InMux I__4912 (
            .O(N__25548),
            .I(N__25517));
    InMux I__4911 (
            .O(N__25545),
            .I(N__25514));
    Span4Mux_v I__4910 (
            .O(N__25540),
            .I(N__25511));
    Odrv12 I__4909 (
            .O(N__25537),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    Odrv4 I__4908 (
            .O(N__25534),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    Odrv4 I__4907 (
            .O(N__25531),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    LocalMux I__4906 (
            .O(N__25528),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    LocalMux I__4905 (
            .O(N__25525),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    LocalMux I__4904 (
            .O(N__25520),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    LocalMux I__4903 (
            .O(N__25517),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    LocalMux I__4902 (
            .O(N__25514),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    Odrv4 I__4901 (
            .O(N__25511),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    InMux I__4900 (
            .O(N__25492),
            .I(N__25489));
    LocalMux I__4899 (
            .O(N__25489),
            .I(\b2v_inst11.mult1_un159_sum_cry_2_s ));
    CascadeMux I__4898 (
            .O(N__25486),
            .I(N__25483));
    InMux I__4897 (
            .O(N__25483),
            .I(N__25480));
    LocalMux I__4896 (
            .O(N__25480),
            .I(\b2v_inst11.mult1_un159_sum_cry_3_s ));
    InMux I__4895 (
            .O(N__25477),
            .I(N__25474));
    LocalMux I__4894 (
            .O(N__25474),
            .I(\b2v_inst11.mult1_un159_sum_cry_4_s ));
    CascadeMux I__4893 (
            .O(N__25471),
            .I(N__25468));
    InMux I__4892 (
            .O(N__25468),
            .I(N__25457));
    InMux I__4891 (
            .O(N__25467),
            .I(N__25457));
    InMux I__4890 (
            .O(N__25466),
            .I(N__25457));
    InMux I__4889 (
            .O(N__25465),
            .I(N__25454));
    InMux I__4888 (
            .O(N__25464),
            .I(N__25451));
    LocalMux I__4887 (
            .O(N__25457),
            .I(\b2v_inst11.mult1_un159_sum_s_7 ));
    LocalMux I__4886 (
            .O(N__25454),
            .I(\b2v_inst11.mult1_un159_sum_s_7 ));
    LocalMux I__4885 (
            .O(N__25451),
            .I(\b2v_inst11.mult1_un159_sum_s_7 ));
    CascadeMux I__4884 (
            .O(N__25444),
            .I(N__25440));
    InMux I__4883 (
            .O(N__25443),
            .I(N__25432));
    InMux I__4882 (
            .O(N__25440),
            .I(N__25432));
    InMux I__4881 (
            .O(N__25439),
            .I(N__25432));
    LocalMux I__4880 (
            .O(N__25432),
            .I(G_2890));
    CascadeMux I__4879 (
            .O(N__25429),
            .I(N__25426));
    InMux I__4878 (
            .O(N__25426),
            .I(N__25423));
    LocalMux I__4877 (
            .O(N__25423),
            .I(N__25420));
    Odrv4 I__4876 (
            .O(N__25420),
            .I(\b2v_inst11.mult1_un159_sum_cry_5_s ));
    InMux I__4875 (
            .O(N__25417),
            .I(N__25414));
    LocalMux I__4874 (
            .O(N__25414),
            .I(\b2v_inst11.mult1_un166_sum_axb_6 ));
    InMux I__4873 (
            .O(N__25411),
            .I(\b2v_inst11.mult1_un166_sum_cry_5 ));
    InMux I__4872 (
            .O(N__25408),
            .I(N__25405));
    LocalMux I__4871 (
            .O(N__25405),
            .I(N__25402));
    Span4Mux_v I__4870 (
            .O(N__25402),
            .I(N__25399));
    Odrv4 I__4869 (
            .O(N__25399),
            .I(\b2v_inst11.un85_clk_100khz_0 ));
    InMux I__4868 (
            .O(N__25396),
            .I(N__25393));
    LocalMux I__4867 (
            .O(N__25393),
            .I(N__25386));
    CascadeMux I__4866 (
            .O(N__25392),
            .I(N__25380));
    InMux I__4865 (
            .O(N__25391),
            .I(N__25376));
    InMux I__4864 (
            .O(N__25390),
            .I(N__25371));
    InMux I__4863 (
            .O(N__25389),
            .I(N__25371));
    Span4Mux_v I__4862 (
            .O(N__25386),
            .I(N__25368));
    InMux I__4861 (
            .O(N__25385),
            .I(N__25365));
    InMux I__4860 (
            .O(N__25384),
            .I(N__25361));
    InMux I__4859 (
            .O(N__25383),
            .I(N__25355));
    InMux I__4858 (
            .O(N__25380),
            .I(N__25355));
    InMux I__4857 (
            .O(N__25379),
            .I(N__25352));
    LocalMux I__4856 (
            .O(N__25376),
            .I(N__25347));
    LocalMux I__4855 (
            .O(N__25371),
            .I(N__25347));
    Span4Mux_h I__4854 (
            .O(N__25368),
            .I(N__25341));
    LocalMux I__4853 (
            .O(N__25365),
            .I(N__25341));
    InMux I__4852 (
            .O(N__25364),
            .I(N__25338));
    LocalMux I__4851 (
            .O(N__25361),
            .I(N__25334));
    CascadeMux I__4850 (
            .O(N__25360),
            .I(N__25330));
    LocalMux I__4849 (
            .O(N__25355),
            .I(N__25327));
    LocalMux I__4848 (
            .O(N__25352),
            .I(N__25322));
    Span4Mux_v I__4847 (
            .O(N__25347),
            .I(N__25322));
    InMux I__4846 (
            .O(N__25346),
            .I(N__25319));
    Span4Mux_v I__4845 (
            .O(N__25341),
            .I(N__25315));
    LocalMux I__4844 (
            .O(N__25338),
            .I(N__25312));
    CascadeMux I__4843 (
            .O(N__25337),
            .I(N__25309));
    Span4Mux_v I__4842 (
            .O(N__25334),
            .I(N__25305));
    InMux I__4841 (
            .O(N__25333),
            .I(N__25300));
    InMux I__4840 (
            .O(N__25330),
            .I(N__25300));
    Span4Mux_h I__4839 (
            .O(N__25327),
            .I(N__25293));
    Span4Mux_v I__4838 (
            .O(N__25322),
            .I(N__25293));
    LocalMux I__4837 (
            .O(N__25319),
            .I(N__25293));
    InMux I__4836 (
            .O(N__25318),
            .I(N__25290));
    Span4Mux_v I__4835 (
            .O(N__25315),
            .I(N__25285));
    Span4Mux_s3_v I__4834 (
            .O(N__25312),
            .I(N__25285));
    InMux I__4833 (
            .O(N__25309),
            .I(N__25282));
    InMux I__4832 (
            .O(N__25308),
            .I(N__25279));
    Span4Mux_v I__4831 (
            .O(N__25305),
            .I(N__25274));
    LocalMux I__4830 (
            .O(N__25300),
            .I(N__25274));
    Span4Mux_s3_v I__4829 (
            .O(N__25293),
            .I(N__25271));
    LocalMux I__4828 (
            .O(N__25290),
            .I(N__25268));
    Odrv4 I__4827 (
            .O(N__25285),
            .I(\b2v_inst11.dutycycle ));
    LocalMux I__4826 (
            .O(N__25282),
            .I(\b2v_inst11.dutycycle ));
    LocalMux I__4825 (
            .O(N__25279),
            .I(\b2v_inst11.dutycycle ));
    Odrv4 I__4824 (
            .O(N__25274),
            .I(\b2v_inst11.dutycycle ));
    Odrv4 I__4823 (
            .O(N__25271),
            .I(\b2v_inst11.dutycycle ));
    Odrv4 I__4822 (
            .O(N__25268),
            .I(\b2v_inst11.dutycycle ));
    CascadeMux I__4821 (
            .O(N__25255),
            .I(N__25252));
    InMux I__4820 (
            .O(N__25252),
            .I(N__25249));
    LocalMux I__4819 (
            .O(N__25249),
            .I(\b2v_inst11.mult1_un159_sum_i ));
    InMux I__4818 (
            .O(N__25246),
            .I(\b2v_inst36.un2_count_1_cry_13 ));
    InMux I__4817 (
            .O(N__25243),
            .I(\b2v_inst36.un2_count_1_cry_14 ));
    InMux I__4816 (
            .O(N__25240),
            .I(N__25237));
    LocalMux I__4815 (
            .O(N__25237),
            .I(\b2v_inst36.count_1_12 ));
    CascadeMux I__4814 (
            .O(N__25234),
            .I(\b2v_inst36.count_en_cascade_ ));
    InMux I__4813 (
            .O(N__25231),
            .I(N__25225));
    InMux I__4812 (
            .O(N__25230),
            .I(N__25225));
    LocalMux I__4811 (
            .O(N__25225),
            .I(\b2v_inst36.count_rst_2 ));
    InMux I__4810 (
            .O(N__25222),
            .I(N__25218));
    InMux I__4809 (
            .O(N__25221),
            .I(N__25215));
    LocalMux I__4808 (
            .O(N__25218),
            .I(\b2v_inst36.count_rst_0 ));
    LocalMux I__4807 (
            .O(N__25215),
            .I(\b2v_inst36.count_rst_0 ));
    InMux I__4806 (
            .O(N__25210),
            .I(N__25207));
    LocalMux I__4805 (
            .O(N__25207),
            .I(N__25204));
    Odrv4 I__4804 (
            .O(N__25204),
            .I(\b2v_inst36.count_1_14 ));
    CascadeMux I__4803 (
            .O(N__25201),
            .I(N__25198));
    InMux I__4802 (
            .O(N__25198),
            .I(N__25192));
    InMux I__4801 (
            .O(N__25197),
            .I(N__25192));
    LocalMux I__4800 (
            .O(N__25192),
            .I(\b2v_inst36.count_rst ));
    InMux I__4799 (
            .O(N__25189),
            .I(N__25186));
    LocalMux I__4798 (
            .O(N__25186),
            .I(\b2v_inst36.count_1_15 ));
    InMux I__4797 (
            .O(N__25183),
            .I(\b2v_inst36.un2_count_1_cry_5 ));
    InMux I__4796 (
            .O(N__25180),
            .I(N__25176));
    CascadeMux I__4795 (
            .O(N__25179),
            .I(N__25173));
    LocalMux I__4794 (
            .O(N__25176),
            .I(N__25169));
    InMux I__4793 (
            .O(N__25173),
            .I(N__25166));
    InMux I__4792 (
            .O(N__25172),
            .I(N__25163));
    Odrv4 I__4791 (
            .O(N__25169),
            .I(\b2v_inst36.countZ0Z_7 ));
    LocalMux I__4790 (
            .O(N__25166),
            .I(\b2v_inst36.countZ0Z_7 ));
    LocalMux I__4789 (
            .O(N__25163),
            .I(\b2v_inst36.countZ0Z_7 ));
    InMux I__4788 (
            .O(N__25156),
            .I(N__25153));
    LocalMux I__4787 (
            .O(N__25153),
            .I(N__25149));
    InMux I__4786 (
            .O(N__25152),
            .I(N__25146));
    Odrv4 I__4785 (
            .O(N__25149),
            .I(\b2v_inst36.un2_count_1_cry_6_THRU_CO ));
    LocalMux I__4784 (
            .O(N__25146),
            .I(\b2v_inst36.un2_count_1_cry_6_THRU_CO ));
    InMux I__4783 (
            .O(N__25141),
            .I(\b2v_inst36.un2_count_1_cry_6 ));
    CascadeMux I__4782 (
            .O(N__25138),
            .I(N__25134));
    InMux I__4781 (
            .O(N__25137),
            .I(N__25131));
    InMux I__4780 (
            .O(N__25134),
            .I(N__25128));
    LocalMux I__4779 (
            .O(N__25131),
            .I(\b2v_inst36.un2_count_1_cry_7_THRU_CO ));
    LocalMux I__4778 (
            .O(N__25128),
            .I(\b2v_inst36.un2_count_1_cry_7_THRU_CO ));
    InMux I__4777 (
            .O(N__25123),
            .I(\b2v_inst36.un2_count_1_cry_7 ));
    InMux I__4776 (
            .O(N__25120),
            .I(bfn_9_2_0_));
    InMux I__4775 (
            .O(N__25117),
            .I(N__25111));
    InMux I__4774 (
            .O(N__25116),
            .I(N__25111));
    LocalMux I__4773 (
            .O(N__25111),
            .I(\b2v_inst36.un2_count_1_cry_9_THRU_CO ));
    InMux I__4772 (
            .O(N__25108),
            .I(\b2v_inst36.un2_count_1_cry_9 ));
    InMux I__4771 (
            .O(N__25105),
            .I(\b2v_inst36.un2_count_1_cry_10 ));
    InMux I__4770 (
            .O(N__25102),
            .I(\b2v_inst36.un2_count_1_cry_11 ));
    InMux I__4769 (
            .O(N__25099),
            .I(\b2v_inst36.un2_count_1_cry_12 ));
    IoInMux I__4768 (
            .O(N__25096),
            .I(N__25093));
    LocalMux I__4767 (
            .O(N__25093),
            .I(N__25090));
    IoSpan4Mux I__4766 (
            .O(N__25090),
            .I(N__25087));
    Span4Mux_s3_h I__4765 (
            .O(N__25087),
            .I(N__25082));
    InMux I__4764 (
            .O(N__25086),
            .I(N__25079));
    CascadeMux I__4763 (
            .O(N__25085),
            .I(N__25074));
    Span4Mux_v I__4762 (
            .O(N__25082),
            .I(N__25068));
    LocalMux I__4761 (
            .O(N__25079),
            .I(N__25068));
    InMux I__4760 (
            .O(N__25078),
            .I(N__25056));
    InMux I__4759 (
            .O(N__25077),
            .I(N__25056));
    InMux I__4758 (
            .O(N__25074),
            .I(N__25056));
    InMux I__4757 (
            .O(N__25073),
            .I(N__25056));
    Span4Mux_v I__4756 (
            .O(N__25068),
            .I(N__25052));
    InMux I__4755 (
            .O(N__25067),
            .I(N__25047));
    InMux I__4754 (
            .O(N__25066),
            .I(N__25047));
    InMux I__4753 (
            .O(N__25065),
            .I(N__25044));
    LocalMux I__4752 (
            .O(N__25056),
            .I(N__25041));
    InMux I__4751 (
            .O(N__25055),
            .I(N__25038));
    Span4Mux_s0_v I__4750 (
            .O(N__25052),
            .I(N__25033));
    LocalMux I__4749 (
            .O(N__25047),
            .I(N__25033));
    LocalMux I__4748 (
            .O(N__25044),
            .I(N__25030));
    Span4Mux_h I__4747 (
            .O(N__25041),
            .I(N__25027));
    LocalMux I__4746 (
            .O(N__25038),
            .I(N__25022));
    Span4Mux_h I__4745 (
            .O(N__25033),
            .I(N__25022));
    Span4Mux_h I__4744 (
            .O(N__25030),
            .I(N__25019));
    Span4Mux_v I__4743 (
            .O(N__25027),
            .I(N__25016));
    Span4Mux_v I__4742 (
            .O(N__25022),
            .I(N__25013));
    Odrv4 I__4741 (
            .O(N__25019),
            .I(SYNTHESIZED_WIRE_49_i_0_o3_0));
    Odrv4 I__4740 (
            .O(N__25016),
            .I(SYNTHESIZED_WIRE_49_i_0_o3_0));
    Odrv4 I__4739 (
            .O(N__25013),
            .I(SYNTHESIZED_WIRE_49_i_0_o3_0));
    InMux I__4738 (
            .O(N__25006),
            .I(N__25003));
    LocalMux I__4737 (
            .O(N__25003),
            .I(N__25000));
    Span4Mux_v I__4736 (
            .O(N__25000),
            .I(N__24997));
    Odrv4 I__4735 (
            .O(N__24997),
            .I(VPP_OK_c));
    IoInMux I__4734 (
            .O(N__24994),
            .I(N__24991));
    LocalMux I__4733 (
            .O(N__24991),
            .I(N__24988));
    IoSpan4Mux I__4732 (
            .O(N__24988),
            .I(N__24985));
    Odrv4 I__4731 (
            .O(N__24985),
            .I(VDDQ_EN_c));
    InMux I__4730 (
            .O(N__24982),
            .I(N__24979));
    LocalMux I__4729 (
            .O(N__24979),
            .I(VCCIO_OK_c));
    InMux I__4728 (
            .O(N__24976),
            .I(N__24973));
    LocalMux I__4727 (
            .O(N__24973),
            .I(V5S_OK_c));
    CascadeMux I__4726 (
            .O(N__24970),
            .I(N__24967));
    InMux I__4725 (
            .O(N__24967),
            .I(N__24964));
    LocalMux I__4724 (
            .O(N__24964),
            .I(\b2v_inst31.un8_outputZ0Z_0 ));
    InMux I__4723 (
            .O(N__24961),
            .I(N__24958));
    LocalMux I__4722 (
            .O(N__24958),
            .I(V33S_OK_c));
    IoInMux I__4721 (
            .O(N__24955),
            .I(N__24951));
    IoInMux I__4720 (
            .O(N__24954),
            .I(N__24948));
    LocalMux I__4719 (
            .O(N__24951),
            .I(N__24943));
    LocalMux I__4718 (
            .O(N__24948),
            .I(N__24943));
    IoSpan4Mux I__4717 (
            .O(N__24943),
            .I(N__24940));
    Span4Mux_s1_h I__4716 (
            .O(N__24940),
            .I(N__24937));
    Span4Mux_h I__4715 (
            .O(N__24937),
            .I(N__24934));
    Odrv4 I__4714 (
            .O(N__24934),
            .I(VCCIN_EN_c));
    InMux I__4713 (
            .O(N__24931),
            .I(\b2v_inst36.un2_count_1_cry_1 ));
    InMux I__4712 (
            .O(N__24928),
            .I(\b2v_inst36.un2_count_1_cry_2 ));
    InMux I__4711 (
            .O(N__24925),
            .I(\b2v_inst36.un2_count_1_cry_3 ));
    CascadeMux I__4710 (
            .O(N__24922),
            .I(N__24919));
    InMux I__4709 (
            .O(N__24919),
            .I(N__24912));
    InMux I__4708 (
            .O(N__24918),
            .I(N__24912));
    InMux I__4707 (
            .O(N__24917),
            .I(N__24909));
    LocalMux I__4706 (
            .O(N__24912),
            .I(\b2v_inst36.countZ0Z_5 ));
    LocalMux I__4705 (
            .O(N__24909),
            .I(\b2v_inst36.countZ0Z_5 ));
    InMux I__4704 (
            .O(N__24904),
            .I(N__24898));
    InMux I__4703 (
            .O(N__24903),
            .I(N__24898));
    LocalMux I__4702 (
            .O(N__24898),
            .I(\b2v_inst36.un2_count_1_cry_4_THRU_CO ));
    InMux I__4701 (
            .O(N__24895),
            .I(\b2v_inst36.un2_count_1_cry_4 ));
    InMux I__4700 (
            .O(N__24892),
            .I(N__24889));
    LocalMux I__4699 (
            .O(N__24889),
            .I(\b2v_inst11.un1_clk_100khz_26_and_i_o2_1 ));
    InMux I__4698 (
            .O(N__24886),
            .I(N__24883));
    LocalMux I__4697 (
            .O(N__24883),
            .I(N__24880));
    Odrv12 I__4696 (
            .O(N__24880),
            .I(\b2v_inst11.dutycycle_RNINJ641_0Z0Z_5 ));
    CascadeMux I__4695 (
            .O(N__24877),
            .I(\b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_cascade_ ));
    InMux I__4694 (
            .O(N__24874),
            .I(N__24871));
    LocalMux I__4693 (
            .O(N__24871),
            .I(\b2v_inst11.N_183 ));
    InMux I__4692 (
            .O(N__24868),
            .I(N__24864));
    InMux I__4691 (
            .O(N__24867),
            .I(N__24861));
    LocalMux I__4690 (
            .O(N__24864),
            .I(N__24858));
    LocalMux I__4689 (
            .O(N__24861),
            .I(N__24855));
    Span12Mux_s4_h I__4688 (
            .O(N__24858),
            .I(N__24851));
    Span4Mux_h I__4687 (
            .O(N__24855),
            .I(N__24848));
    InMux I__4686 (
            .O(N__24854),
            .I(N__24845));
    Odrv12 I__4685 (
            .O(N__24851),
            .I(\b2v_inst11.func_state_RNI_3Z0Z_1 ));
    Odrv4 I__4684 (
            .O(N__24848),
            .I(\b2v_inst11.func_state_RNI_3Z0Z_1 ));
    LocalMux I__4683 (
            .O(N__24845),
            .I(\b2v_inst11.func_state_RNI_3Z0Z_1 ));
    CascadeMux I__4682 (
            .O(N__24838),
            .I(\b2v_inst11.N_183_cascade_ ));
    InMux I__4681 (
            .O(N__24835),
            .I(N__24832));
    LocalMux I__4680 (
            .O(N__24832),
            .I(N__24828));
    InMux I__4679 (
            .O(N__24831),
            .I(N__24825));
    Odrv4 I__4678 (
            .O(N__24828),
            .I(\b2v_inst11.N_114_f0_1 ));
    LocalMux I__4677 (
            .O(N__24825),
            .I(\b2v_inst11.N_114_f0_1 ));
    InMux I__4676 (
            .O(N__24820),
            .I(N__24813));
    InMux I__4675 (
            .O(N__24819),
            .I(N__24809));
    InMux I__4674 (
            .O(N__24818),
            .I(N__24802));
    InMux I__4673 (
            .O(N__24817),
            .I(N__24802));
    CascadeMux I__4672 (
            .O(N__24816),
            .I(N__24799));
    LocalMux I__4671 (
            .O(N__24813),
            .I(N__24796));
    CascadeMux I__4670 (
            .O(N__24812),
            .I(N__24792));
    LocalMux I__4669 (
            .O(N__24809),
            .I(N__24789));
    CascadeMux I__4668 (
            .O(N__24808),
            .I(N__24786));
    CascadeMux I__4667 (
            .O(N__24807),
            .I(N__24783));
    LocalMux I__4666 (
            .O(N__24802),
            .I(N__24776));
    InMux I__4665 (
            .O(N__24799),
            .I(N__24773));
    Span4Mux_v I__4664 (
            .O(N__24796),
            .I(N__24770));
    InMux I__4663 (
            .O(N__24795),
            .I(N__24767));
    InMux I__4662 (
            .O(N__24792),
            .I(N__24764));
    Span12Mux_s10_v I__4661 (
            .O(N__24789),
            .I(N__24761));
    InMux I__4660 (
            .O(N__24786),
            .I(N__24754));
    InMux I__4659 (
            .O(N__24783),
            .I(N__24754));
    InMux I__4658 (
            .O(N__24782),
            .I(N__24754));
    InMux I__4657 (
            .O(N__24781),
            .I(N__24749));
    InMux I__4656 (
            .O(N__24780),
            .I(N__24749));
    InMux I__4655 (
            .O(N__24779),
            .I(N__24746));
    Span4Mux_h I__4654 (
            .O(N__24776),
            .I(N__24741));
    LocalMux I__4653 (
            .O(N__24773),
            .I(N__24741));
    Odrv4 I__4652 (
            .O(N__24770),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__4651 (
            .O(N__24767),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__4650 (
            .O(N__24764),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    Odrv12 I__4649 (
            .O(N__24761),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__4648 (
            .O(N__24754),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__4647 (
            .O(N__24749),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__4646 (
            .O(N__24746),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    Odrv4 I__4645 (
            .O(N__24741),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    InMux I__4644 (
            .O(N__24724),
            .I(N__24717));
    InMux I__4643 (
            .O(N__24723),
            .I(N__24717));
    InMux I__4642 (
            .O(N__24722),
            .I(N__24713));
    LocalMux I__4641 (
            .O(N__24717),
            .I(N__24710));
    InMux I__4640 (
            .O(N__24716),
            .I(N__24707));
    LocalMux I__4639 (
            .O(N__24713),
            .I(N__24702));
    Span4Mux_s1_v I__4638 (
            .O(N__24710),
            .I(N__24702));
    LocalMux I__4637 (
            .O(N__24707),
            .I(\b2v_inst11.N_379 ));
    Odrv4 I__4636 (
            .O(N__24702),
            .I(\b2v_inst11.N_379 ));
    CascadeMux I__4635 (
            .O(N__24697),
            .I(\b2v_inst6.curr_state_RNI8OKQ2Z0Z_0_cascade_ ));
    CascadeMux I__4634 (
            .O(N__24694),
            .I(N__24691));
    InMux I__4633 (
            .O(N__24691),
            .I(N__24684));
    InMux I__4632 (
            .O(N__24690),
            .I(N__24684));
    CascadeMux I__4631 (
            .O(N__24689),
            .I(N__24681));
    LocalMux I__4630 (
            .O(N__24684),
            .I(N__24678));
    InMux I__4629 (
            .O(N__24681),
            .I(N__24672));
    Span4Mux_s1_v I__4628 (
            .O(N__24678),
            .I(N__24669));
    InMux I__4627 (
            .O(N__24677),
            .I(N__24664));
    InMux I__4626 (
            .O(N__24676),
            .I(N__24664));
    InMux I__4625 (
            .O(N__24675),
            .I(N__24661));
    LocalMux I__4624 (
            .O(N__24672),
            .I(\b2v_inst11.un1_clk_100khz_52_and_i_a2Z0Z_1 ));
    Odrv4 I__4623 (
            .O(N__24669),
            .I(\b2v_inst11.un1_clk_100khz_52_and_i_a2Z0Z_1 ));
    LocalMux I__4622 (
            .O(N__24664),
            .I(\b2v_inst11.un1_clk_100khz_52_and_i_a2Z0Z_1 ));
    LocalMux I__4621 (
            .O(N__24661),
            .I(\b2v_inst11.un1_clk_100khz_52_and_i_a2Z0Z_1 ));
    InMux I__4620 (
            .O(N__24652),
            .I(N__24648));
    InMux I__4619 (
            .O(N__24651),
            .I(N__24645));
    LocalMux I__4618 (
            .O(N__24648),
            .I(N__24642));
    LocalMux I__4617 (
            .O(N__24645),
            .I(N__24639));
    Span4Mux_h I__4616 (
            .O(N__24642),
            .I(N__24636));
    Span4Mux_h I__4615 (
            .O(N__24639),
            .I(N__24633));
    Odrv4 I__4614 (
            .O(N__24636),
            .I(\b2v_inst11.func_state_RNIDINH9Z0Z_0 ));
    Odrv4 I__4613 (
            .O(N__24633),
            .I(\b2v_inst11.func_state_RNIDINH9Z0Z_0 ));
    CascadeMux I__4612 (
            .O(N__24628),
            .I(N__24625));
    InMux I__4611 (
            .O(N__24625),
            .I(N__24621));
    InMux I__4610 (
            .O(N__24624),
            .I(N__24618));
    LocalMux I__4609 (
            .O(N__24621),
            .I(N__24615));
    LocalMux I__4608 (
            .O(N__24618),
            .I(\b2v_inst11.func_stateZ0Z_1 ));
    Odrv4 I__4607 (
            .O(N__24615),
            .I(\b2v_inst11.func_stateZ0Z_1 ));
    InMux I__4606 (
            .O(N__24610),
            .I(N__24607));
    LocalMux I__4605 (
            .O(N__24607),
            .I(\b2v_inst6.curr_state_RNI8OKQ2Z0Z_0 ));
    CascadeMux I__4604 (
            .O(N__24604),
            .I(N__24601));
    InMux I__4603 (
            .O(N__24601),
            .I(N__24595));
    InMux I__4602 (
            .O(N__24600),
            .I(N__24595));
    LocalMux I__4601 (
            .O(N__24595),
            .I(\b2v_inst6.delayed_vccin_vccinaux_ok_0 ));
    CascadeMux I__4600 (
            .O(N__24592),
            .I(\b2v_inst11.func_state_cascade_ ));
    CascadeMux I__4599 (
            .O(N__24589),
            .I(\b2v_inst11.N_303_cascade_ ));
    InMux I__4598 (
            .O(N__24586),
            .I(N__24583));
    LocalMux I__4597 (
            .O(N__24583),
            .I(\b2v_inst11.dutycycle_eena_1 ));
    CascadeMux I__4596 (
            .O(N__24580),
            .I(N__24576));
    InMux I__4595 (
            .O(N__24579),
            .I(N__24573));
    InMux I__4594 (
            .O(N__24576),
            .I(N__24570));
    LocalMux I__4593 (
            .O(N__24573),
            .I(N__24567));
    LocalMux I__4592 (
            .O(N__24570),
            .I(N__24564));
    Span4Mux_h I__4591 (
            .O(N__24567),
            .I(N__24559));
    Span4Mux_h I__4590 (
            .O(N__24564),
            .I(N__24559));
    Odrv4 I__4589 (
            .O(N__24559),
            .I(\b2v_inst11.N_70 ));
    CascadeMux I__4588 (
            .O(N__24556),
            .I(\b2v_inst11.dutycycle_eena_1_cascade_ ));
    InMux I__4587 (
            .O(N__24553),
            .I(N__24547));
    InMux I__4586 (
            .O(N__24552),
            .I(N__24547));
    LocalMux I__4585 (
            .O(N__24547),
            .I(\b2v_inst11.dutycycleZ1Z_2 ));
    CascadeMux I__4584 (
            .O(N__24544),
            .I(N__24541));
    InMux I__4583 (
            .O(N__24541),
            .I(N__24538));
    LocalMux I__4582 (
            .O(N__24538),
            .I(N__24534));
    InMux I__4581 (
            .O(N__24537),
            .I(N__24531));
    Odrv4 I__4580 (
            .O(N__24534),
            .I(\b2v_inst11.dutycycle_eena_0 ));
    LocalMux I__4579 (
            .O(N__24531),
            .I(\b2v_inst11.dutycycle_eena_0 ));
    InMux I__4578 (
            .O(N__24526),
            .I(N__24522));
    InMux I__4577 (
            .O(N__24525),
            .I(N__24519));
    LocalMux I__4576 (
            .O(N__24522),
            .I(N__24516));
    LocalMux I__4575 (
            .O(N__24519),
            .I(N__24513));
    Span4Mux_v I__4574 (
            .O(N__24516),
            .I(N__24508));
    Span4Mux_h I__4573 (
            .O(N__24513),
            .I(N__24505));
    InMux I__4572 (
            .O(N__24512),
            .I(N__24500));
    InMux I__4571 (
            .O(N__24511),
            .I(N__24500));
    Odrv4 I__4570 (
            .O(N__24508),
            .I(\b2v_inst11.N_169 ));
    Odrv4 I__4569 (
            .O(N__24505),
            .I(\b2v_inst11.N_169 ));
    LocalMux I__4568 (
            .O(N__24500),
            .I(\b2v_inst11.N_169 ));
    InMux I__4567 (
            .O(N__24493),
            .I(N__24490));
    LocalMux I__4566 (
            .O(N__24490),
            .I(\b2v_inst11.N_375 ));
    CascadeMux I__4565 (
            .O(N__24487),
            .I(\b2v_inst11.un1_clk_100khz_52_and_i_a2_1_sxZ0_cascade_ ));
    InMux I__4564 (
            .O(N__24484),
            .I(N__24478));
    InMux I__4563 (
            .O(N__24483),
            .I(N__24473));
    InMux I__4562 (
            .O(N__24482),
            .I(N__24473));
    CascadeMux I__4561 (
            .O(N__24481),
            .I(N__24470));
    LocalMux I__4560 (
            .O(N__24478),
            .I(N__24465));
    LocalMux I__4559 (
            .O(N__24473),
            .I(N__24461));
    InMux I__4558 (
            .O(N__24470),
            .I(N__24456));
    InMux I__4557 (
            .O(N__24469),
            .I(N__24456));
    CascadeMux I__4556 (
            .O(N__24468),
            .I(N__24452));
    Span4Mux_h I__4555 (
            .O(N__24465),
            .I(N__24449));
    InMux I__4554 (
            .O(N__24464),
            .I(N__24446));
    Sp12to4 I__4553 (
            .O(N__24461),
            .I(N__24441));
    LocalMux I__4552 (
            .O(N__24456),
            .I(N__24441));
    InMux I__4551 (
            .O(N__24455),
            .I(N__24436));
    InMux I__4550 (
            .O(N__24452),
            .I(N__24436));
    Odrv4 I__4549 (
            .O(N__24449),
            .I(SYNTHESIZED_WIRE_47keep_fast));
    LocalMux I__4548 (
            .O(N__24446),
            .I(SYNTHESIZED_WIRE_47keep_fast));
    Odrv12 I__4547 (
            .O(N__24441),
            .I(SYNTHESIZED_WIRE_47keep_fast));
    LocalMux I__4546 (
            .O(N__24436),
            .I(SYNTHESIZED_WIRE_47keep_fast));
    InMux I__4545 (
            .O(N__24427),
            .I(N__24424));
    LocalMux I__4544 (
            .O(N__24424),
            .I(\b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_1 ));
    InMux I__4543 (
            .O(N__24421),
            .I(N__24418));
    LocalMux I__4542 (
            .O(N__24418),
            .I(N__24415));
    Odrv12 I__4541 (
            .O(N__24415),
            .I(\b2v_inst11.m15_e_3 ));
    InMux I__4540 (
            .O(N__24412),
            .I(N__24409));
    LocalMux I__4539 (
            .O(N__24409),
            .I(\b2v_inst11.un1_dutycycle_inv_4_0 ));
    InMux I__4538 (
            .O(N__24406),
            .I(N__24403));
    LocalMux I__4537 (
            .O(N__24403),
            .I(N__24400));
    Odrv4 I__4536 (
            .O(N__24400),
            .I(\b2v_inst11.g0_9_1 ));
    CascadeMux I__4535 (
            .O(N__24397),
            .I(\b2v_inst11.g1_0_1_cascade_ ));
    InMux I__4534 (
            .O(N__24394),
            .I(N__24390));
    InMux I__4533 (
            .O(N__24393),
            .I(N__24387));
    LocalMux I__4532 (
            .O(N__24390),
            .I(\b2v_inst11.un1_dutycycle_164_0 ));
    LocalMux I__4531 (
            .O(N__24387),
            .I(\b2v_inst11.un1_dutycycle_164_0 ));
    CascadeMux I__4530 (
            .O(N__24382),
            .I(N__24379));
    InMux I__4529 (
            .O(N__24379),
            .I(N__24375));
    CascadeMux I__4528 (
            .O(N__24378),
            .I(N__24372));
    LocalMux I__4527 (
            .O(N__24375),
            .I(N__24369));
    InMux I__4526 (
            .O(N__24372),
            .I(N__24366));
    Span4Mux_v I__4525 (
            .O(N__24369),
            .I(N__24361));
    LocalMux I__4524 (
            .O(N__24366),
            .I(N__24358));
    InMux I__4523 (
            .O(N__24365),
            .I(N__24353));
    InMux I__4522 (
            .O(N__24364),
            .I(N__24353));
    Span4Mux_h I__4521 (
            .O(N__24361),
            .I(N__24348));
    Span4Mux_s2_v I__4520 (
            .O(N__24358),
            .I(N__24348));
    LocalMux I__4519 (
            .O(N__24353),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_5 ));
    Odrv4 I__4518 (
            .O(N__24348),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_5 ));
    CascadeMux I__4517 (
            .O(N__24343),
            .I(N__24340));
    InMux I__4516 (
            .O(N__24340),
            .I(N__24337));
    LocalMux I__4515 (
            .O(N__24337),
            .I(N__24334));
    Span12Mux_s5_v I__4514 (
            .O(N__24334),
            .I(N__24331));
    Odrv12 I__4513 (
            .O(N__24331),
            .I(\b2v_inst11.mult1_un152_sum_i ));
    InMux I__4512 (
            .O(N__24328),
            .I(N__24325));
    LocalMux I__4511 (
            .O(N__24325),
            .I(N__24321));
    InMux I__4510 (
            .O(N__24324),
            .I(N__24318));
    Span4Mux_h I__4509 (
            .O(N__24321),
            .I(N__24308));
    LocalMux I__4508 (
            .O(N__24318),
            .I(N__24308));
    InMux I__4507 (
            .O(N__24317),
            .I(N__24305));
    InMux I__4506 (
            .O(N__24316),
            .I(N__24302));
    InMux I__4505 (
            .O(N__24315),
            .I(N__24298));
    InMux I__4504 (
            .O(N__24314),
            .I(N__24295));
    InMux I__4503 (
            .O(N__24313),
            .I(N__24292));
    Span4Mux_h I__4502 (
            .O(N__24308),
            .I(N__24286));
    LocalMux I__4501 (
            .O(N__24305),
            .I(N__24286));
    LocalMux I__4500 (
            .O(N__24302),
            .I(N__24283));
    InMux I__4499 (
            .O(N__24301),
            .I(N__24280));
    LocalMux I__4498 (
            .O(N__24298),
            .I(N__24274));
    LocalMux I__4497 (
            .O(N__24295),
            .I(N__24269));
    LocalMux I__4496 (
            .O(N__24292),
            .I(N__24269));
    InMux I__4495 (
            .O(N__24291),
            .I(N__24266));
    Span4Mux_v I__4494 (
            .O(N__24286),
            .I(N__24259));
    Span4Mux_h I__4493 (
            .O(N__24283),
            .I(N__24259));
    LocalMux I__4492 (
            .O(N__24280),
            .I(N__24259));
    InMux I__4491 (
            .O(N__24279),
            .I(N__24252));
    InMux I__4490 (
            .O(N__24278),
            .I(N__24252));
    InMux I__4489 (
            .O(N__24277),
            .I(N__24252));
    Span4Mux_v I__4488 (
            .O(N__24274),
            .I(N__24247));
    Span4Mux_h I__4487 (
            .O(N__24269),
            .I(N__24247));
    LocalMux I__4486 (
            .O(N__24266),
            .I(\b2v_inst11.N_3013_i ));
    Odrv4 I__4485 (
            .O(N__24259),
            .I(\b2v_inst11.N_3013_i ));
    LocalMux I__4484 (
            .O(N__24252),
            .I(\b2v_inst11.N_3013_i ));
    Odrv4 I__4483 (
            .O(N__24247),
            .I(\b2v_inst11.N_3013_i ));
    SRMux I__4482 (
            .O(N__24238),
            .I(N__24233));
    SRMux I__4481 (
            .O(N__24237),
            .I(N__24228));
    SRMux I__4480 (
            .O(N__24236),
            .I(N__24224));
    LocalMux I__4479 (
            .O(N__24233),
            .I(N__24221));
    SRMux I__4478 (
            .O(N__24232),
            .I(N__24218));
    SRMux I__4477 (
            .O(N__24231),
            .I(N__24215));
    LocalMux I__4476 (
            .O(N__24228),
            .I(N__24211));
    SRMux I__4475 (
            .O(N__24227),
            .I(N__24207));
    LocalMux I__4474 (
            .O(N__24224),
            .I(N__24204));
    Span4Mux_v I__4473 (
            .O(N__24221),
            .I(N__24197));
    LocalMux I__4472 (
            .O(N__24218),
            .I(N__24197));
    LocalMux I__4471 (
            .O(N__24215),
            .I(N__24197));
    SRMux I__4470 (
            .O(N__24214),
            .I(N__24194));
    Span4Mux_h I__4469 (
            .O(N__24211),
            .I(N__24191));
    SRMux I__4468 (
            .O(N__24210),
            .I(N__24188));
    LocalMux I__4467 (
            .O(N__24207),
            .I(N__24184));
    Span4Mux_v I__4466 (
            .O(N__24204),
            .I(N__24179));
    Span4Mux_v I__4465 (
            .O(N__24197),
            .I(N__24179));
    LocalMux I__4464 (
            .O(N__24194),
            .I(N__24176));
    Sp12to4 I__4463 (
            .O(N__24191),
            .I(N__24171));
    LocalMux I__4462 (
            .O(N__24188),
            .I(N__24171));
    SRMux I__4461 (
            .O(N__24187),
            .I(N__24168));
    Span4Mux_h I__4460 (
            .O(N__24184),
            .I(N__24165));
    Span4Mux_h I__4459 (
            .O(N__24179),
            .I(N__24157));
    Span4Mux_v I__4458 (
            .O(N__24176),
            .I(N__24154));
    Span12Mux_s6_v I__4457 (
            .O(N__24171),
            .I(N__24151));
    LocalMux I__4456 (
            .O(N__24168),
            .I(N__24148));
    Span4Mux_v I__4455 (
            .O(N__24165),
            .I(N__24145));
    SRMux I__4454 (
            .O(N__24164),
            .I(N__24142));
    SRMux I__4453 (
            .O(N__24163),
            .I(N__24139));
    SRMux I__4452 (
            .O(N__24162),
            .I(N__24136));
    SRMux I__4451 (
            .O(N__24161),
            .I(N__24133));
    SRMux I__4450 (
            .O(N__24160),
            .I(N__24130));
    Odrv4 I__4449 (
            .O(N__24157),
            .I(\b2v_inst11.N_221_iZ0 ));
    Odrv4 I__4448 (
            .O(N__24154),
            .I(\b2v_inst11.N_221_iZ0 ));
    Odrv12 I__4447 (
            .O(N__24151),
            .I(\b2v_inst11.N_221_iZ0 ));
    Odrv12 I__4446 (
            .O(N__24148),
            .I(\b2v_inst11.N_221_iZ0 ));
    Odrv4 I__4445 (
            .O(N__24145),
            .I(\b2v_inst11.N_221_iZ0 ));
    LocalMux I__4444 (
            .O(N__24142),
            .I(\b2v_inst11.N_221_iZ0 ));
    LocalMux I__4443 (
            .O(N__24139),
            .I(\b2v_inst11.N_221_iZ0 ));
    LocalMux I__4442 (
            .O(N__24136),
            .I(\b2v_inst11.N_221_iZ0 ));
    LocalMux I__4441 (
            .O(N__24133),
            .I(\b2v_inst11.N_221_iZ0 ));
    LocalMux I__4440 (
            .O(N__24130),
            .I(\b2v_inst11.N_221_iZ0 ));
    InMux I__4439 (
            .O(N__24109),
            .I(N__24106));
    LocalMux I__4438 (
            .O(N__24106),
            .I(N__24103));
    Span4Mux_v I__4437 (
            .O(N__24103),
            .I(N__24100));
    Odrv4 I__4436 (
            .O(N__24100),
            .I(\b2v_inst11.g0_1_1 ));
    CascadeMux I__4435 (
            .O(N__24097),
            .I(N__24093));
    InMux I__4434 (
            .O(N__24096),
            .I(N__24089));
    InMux I__4433 (
            .O(N__24093),
            .I(N__24086));
    InMux I__4432 (
            .O(N__24092),
            .I(N__24083));
    LocalMux I__4431 (
            .O(N__24089),
            .I(N__24079));
    LocalMux I__4430 (
            .O(N__24086),
            .I(N__24076));
    LocalMux I__4429 (
            .O(N__24083),
            .I(N__24073));
    InMux I__4428 (
            .O(N__24082),
            .I(N__24070));
    Span4Mux_s2_v I__4427 (
            .O(N__24079),
            .I(N__24067));
    Span4Mux_s2_v I__4426 (
            .O(N__24076),
            .I(N__24062));
    Span4Mux_s2_v I__4425 (
            .O(N__24073),
            .I(N__24062));
    LocalMux I__4424 (
            .O(N__24070),
            .I(N__24059));
    Span4Mux_v I__4423 (
            .O(N__24067),
            .I(N__24055));
    Span4Mux_v I__4422 (
            .O(N__24062),
            .I(N__24052));
    Span4Mux_s3_v I__4421 (
            .O(N__24059),
            .I(N__24049));
    InMux I__4420 (
            .O(N__24058),
            .I(N__24046));
    Odrv4 I__4419 (
            .O(N__24055),
            .I(\b2v_inst11.N_182 ));
    Odrv4 I__4418 (
            .O(N__24052),
            .I(\b2v_inst11.N_182 ));
    Odrv4 I__4417 (
            .O(N__24049),
            .I(\b2v_inst11.N_182 ));
    LocalMux I__4416 (
            .O(N__24046),
            .I(\b2v_inst11.N_182 ));
    CascadeMux I__4415 (
            .O(N__24037),
            .I(N__24034));
    InMux I__4414 (
            .O(N__24034),
            .I(N__24031));
    LocalMux I__4413 (
            .O(N__24031),
            .I(\b2v_inst11.func_state_RNIT4D71_0Z0Z_1 ));
    InMux I__4412 (
            .O(N__24028),
            .I(N__24022));
    InMux I__4411 (
            .O(N__24027),
            .I(N__24022));
    LocalMux I__4410 (
            .O(N__24022),
            .I(\b2v_inst11.dutycycle_0_5 ));
    InMux I__4409 (
            .O(N__24019),
            .I(N__24013));
    InMux I__4408 (
            .O(N__24018),
            .I(N__24013));
    LocalMux I__4407 (
            .O(N__24013),
            .I(N__24010));
    Span4Mux_h I__4406 (
            .O(N__24010),
            .I(N__24007));
    Odrv4 I__4405 (
            .O(N__24007),
            .I(\b2v_inst11.g1_4_0 ));
    CascadeMux I__4404 (
            .O(N__24004),
            .I(\b2v_inst11.func_state_RNIT4D71_0Z0Z_1_cascade_ ));
    CascadeMux I__4403 (
            .O(N__24001),
            .I(dutycycle_RNIIOE3D_0_5_cascade_));
    CascadeMux I__4402 (
            .O(N__23998),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_5_cascade_ ));
    CascadeMux I__4401 (
            .O(N__23995),
            .I(\b2v_inst11.un1_dutycycle_53_axb_3_1_cascade_ ));
    InMux I__4400 (
            .O(N__23992),
            .I(N__23989));
    LocalMux I__4399 (
            .O(N__23989),
            .I(N__23986));
    Span4Mux_h I__4398 (
            .O(N__23986),
            .I(N__23983));
    Span4Mux_v I__4397 (
            .O(N__23983),
            .I(N__23980));
    Odrv4 I__4396 (
            .O(N__23980),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_2 ));
    InMux I__4395 (
            .O(N__23977),
            .I(N__23974));
    LocalMux I__4394 (
            .O(N__23974),
            .I(\b2v_inst11.un1_i3_mux_1 ));
    InMux I__4393 (
            .O(N__23971),
            .I(N__23968));
    LocalMux I__4392 (
            .O(N__23968),
            .I(N__23965));
    Span4Mux_h I__4391 (
            .O(N__23965),
            .I(N__23962));
    Odrv4 I__4390 (
            .O(N__23962),
            .I(\b2v_inst11.g0_6_2 ));
    CascadeMux I__4389 (
            .O(N__23959),
            .I(\b2v_inst5.curr_stateZ0Z_1_cascade_ ));
    CascadeMux I__4388 (
            .O(N__23956),
            .I(curr_state_RNI5VS71_0_1_cascade_));
    InMux I__4387 (
            .O(N__23953),
            .I(N__23950));
    LocalMux I__4386 (
            .O(N__23950),
            .I(N__23946));
    InMux I__4385 (
            .O(N__23949),
            .I(N__23943));
    Span4Mux_s2_v I__4384 (
            .O(N__23946),
            .I(N__23938));
    LocalMux I__4383 (
            .O(N__23943),
            .I(N__23938));
    Span4Mux_v I__4382 (
            .O(N__23938),
            .I(N__23935));
    Odrv4 I__4381 (
            .O(N__23935),
            .I(\b2v_inst11.mult1_un145_sum ));
    CascadeMux I__4380 (
            .O(N__23932),
            .I(RSMRSTn_RNI8DFE_cascade_));
    InMux I__4379 (
            .O(N__23929),
            .I(N__23926));
    LocalMux I__4378 (
            .O(N__23926),
            .I(\b2v_inst11.count_0_11 ));
    InMux I__4377 (
            .O(N__23923),
            .I(N__23917));
    InMux I__4376 (
            .O(N__23922),
            .I(N__23917));
    LocalMux I__4375 (
            .O(N__23917),
            .I(N__23914));
    Odrv4 I__4374 (
            .O(N__23914),
            .I(\b2v_inst11.un1_count_cry_1_c_RNIIIQDZ0 ));
    InMux I__4373 (
            .O(N__23911),
            .I(N__23908));
    LocalMux I__4372 (
            .O(N__23908),
            .I(\b2v_inst11.count_0_2 ));
    InMux I__4371 (
            .O(N__23905),
            .I(N__23901));
    InMux I__4370 (
            .O(N__23904),
            .I(N__23898));
    LocalMux I__4369 (
            .O(N__23901),
            .I(\b2v_inst11.un1_count_cry_11_c_RNI36SZ0Z6 ));
    LocalMux I__4368 (
            .O(N__23898),
            .I(\b2v_inst11.un1_count_cry_11_c_RNI36SZ0Z6 ));
    InMux I__4367 (
            .O(N__23893),
            .I(N__23890));
    LocalMux I__4366 (
            .O(N__23890),
            .I(\b2v_inst11.count_0_12 ));
    CascadeMux I__4365 (
            .O(N__23887),
            .I(G_2727_cascade_));
    InMux I__4364 (
            .O(N__23884),
            .I(N__23881));
    LocalMux I__4363 (
            .O(N__23881),
            .I(\b2v_inst5.curr_state_2_1 ));
    CascadeMux I__4362 (
            .O(N__23878),
            .I(N_229_cascade_));
    InMux I__4361 (
            .O(N__23875),
            .I(N__23863));
    InMux I__4360 (
            .O(N__23874),
            .I(N__23863));
    InMux I__4359 (
            .O(N__23873),
            .I(N__23863));
    InMux I__4358 (
            .O(N__23872),
            .I(N__23863));
    LocalMux I__4357 (
            .O(N__23863),
            .I(\b2v_inst5.curr_stateZ0Z_1 ));
    InMux I__4356 (
            .O(N__23860),
            .I(\b2v_inst11.un1_count_cry_10 ));
    InMux I__4355 (
            .O(N__23857),
            .I(\b2v_inst11.un1_count_cry_11 ));
    InMux I__4354 (
            .O(N__23854),
            .I(\b2v_inst11.un1_count_cry_12 ));
    CascadeMux I__4353 (
            .O(N__23851),
            .I(N__23848));
    InMux I__4352 (
            .O(N__23848),
            .I(N__23842));
    InMux I__4351 (
            .O(N__23847),
            .I(N__23842));
    LocalMux I__4350 (
            .O(N__23842),
            .I(N__23839));
    Odrv4 I__4349 (
            .O(N__23839),
            .I(\b2v_inst11.un1_count_cry_13_c_RNI5AUZ0Z6 ));
    InMux I__4348 (
            .O(N__23836),
            .I(\b2v_inst11.un1_count_cry_13 ));
    InMux I__4347 (
            .O(N__23833),
            .I(\b2v_inst11.un1_count_cry_14 ));
    CascadeMux I__4346 (
            .O(N__23830),
            .I(N__23827));
    InMux I__4345 (
            .O(N__23827),
            .I(N__23821));
    InMux I__4344 (
            .O(N__23826),
            .I(N__23821));
    LocalMux I__4343 (
            .O(N__23821),
            .I(N__23818));
    Odrv4 I__4342 (
            .O(N__23818),
            .I(\b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6 ));
    CascadeMux I__4341 (
            .O(N__23815),
            .I(N__23811));
    InMux I__4340 (
            .O(N__23814),
            .I(N__23806));
    InMux I__4339 (
            .O(N__23811),
            .I(N__23806));
    LocalMux I__4338 (
            .O(N__23806),
            .I(\b2v_inst11.un1_count_cry_9_c_RNIQ23EZ0 ));
    InMux I__4337 (
            .O(N__23803),
            .I(N__23800));
    LocalMux I__4336 (
            .O(N__23800),
            .I(\b2v_inst11.count_0_10 ));
    InMux I__4335 (
            .O(N__23797),
            .I(N__23791));
    InMux I__4334 (
            .O(N__23796),
            .I(N__23791));
    LocalMux I__4333 (
            .O(N__23791),
            .I(\b2v_inst11.un1_count_cry_10_c_RNI24RZ0Z6 ));
    InMux I__4332 (
            .O(N__23788),
            .I(\b2v_inst11.un1_count_cry_1 ));
    InMux I__4331 (
            .O(N__23785),
            .I(\b2v_inst11.un1_count_cry_2 ));
    InMux I__4330 (
            .O(N__23782),
            .I(\b2v_inst11.un1_count_cry_3 ));
    InMux I__4329 (
            .O(N__23779),
            .I(\b2v_inst11.un1_count_cry_4 ));
    InMux I__4328 (
            .O(N__23776),
            .I(N__23770));
    InMux I__4327 (
            .O(N__23775),
            .I(N__23770));
    LocalMux I__4326 (
            .O(N__23770),
            .I(\b2v_inst11.un1_count_cry_5_c_RNIMQUDZ0 ));
    InMux I__4325 (
            .O(N__23767),
            .I(\b2v_inst11.un1_count_cry_5 ));
    InMux I__4324 (
            .O(N__23764),
            .I(N__23758));
    InMux I__4323 (
            .O(N__23763),
            .I(N__23758));
    LocalMux I__4322 (
            .O(N__23758),
            .I(\b2v_inst11.un1_count_cry_6_c_RNINSVDZ0 ));
    InMux I__4321 (
            .O(N__23755),
            .I(\b2v_inst11.un1_count_cry_6 ));
    InMux I__4320 (
            .O(N__23752),
            .I(\b2v_inst11.un1_count_cry_7 ));
    InMux I__4319 (
            .O(N__23749),
            .I(bfn_8_7_0_));
    InMux I__4318 (
            .O(N__23746),
            .I(\b2v_inst11.un1_count_cry_9 ));
    InMux I__4317 (
            .O(N__23743),
            .I(N__23740));
    LocalMux I__4316 (
            .O(N__23740),
            .I(\b2v_inst11.count_0_14 ));
    InMux I__4315 (
            .O(N__23737),
            .I(N__23734));
    LocalMux I__4314 (
            .O(N__23734),
            .I(\b2v_inst11.count_0_6 ));
    InMux I__4313 (
            .O(N__23731),
            .I(N__23728));
    LocalMux I__4312 (
            .O(N__23728),
            .I(\b2v_inst11.count_0_15 ));
    InMux I__4311 (
            .O(N__23725),
            .I(N__23722));
    LocalMux I__4310 (
            .O(N__23722),
            .I(\b2v_inst11.count_0_7 ));
    CascadeMux I__4309 (
            .O(N__23719),
            .I(N__23715));
    InMux I__4308 (
            .O(N__23718),
            .I(N__23710));
    InMux I__4307 (
            .O(N__23715),
            .I(N__23702));
    InMux I__4306 (
            .O(N__23714),
            .I(N__23702));
    InMux I__4305 (
            .O(N__23713),
            .I(N__23702));
    LocalMux I__4304 (
            .O(N__23710),
            .I(N__23699));
    InMux I__4303 (
            .O(N__23709),
            .I(N__23696));
    LocalMux I__4302 (
            .O(N__23702),
            .I(\b2v_inst11.mult1_un145_sum_s_8 ));
    Odrv4 I__4301 (
            .O(N__23699),
            .I(\b2v_inst11.mult1_un145_sum_s_8 ));
    LocalMux I__4300 (
            .O(N__23696),
            .I(\b2v_inst11.mult1_un145_sum_s_8 ));
    CascadeMux I__4299 (
            .O(N__23689),
            .I(N__23685));
    InMux I__4298 (
            .O(N__23688),
            .I(N__23677));
    InMux I__4297 (
            .O(N__23685),
            .I(N__23677));
    InMux I__4296 (
            .O(N__23684),
            .I(N__23677));
    LocalMux I__4295 (
            .O(N__23677),
            .I(\b2v_inst11.mult1_un145_sum_i_0_8 ));
    InMux I__4294 (
            .O(N__23674),
            .I(\b2v_inst11.mult1_un159_sum_cry_1 ));
    InMux I__4293 (
            .O(N__23671),
            .I(N__23668));
    LocalMux I__4292 (
            .O(N__23668),
            .I(\b2v_inst11.mult1_un152_sum_cry_3_s ));
    InMux I__4291 (
            .O(N__23665),
            .I(\b2v_inst11.mult1_un159_sum_cry_2 ));
    CascadeMux I__4290 (
            .O(N__23662),
            .I(N__23659));
    InMux I__4289 (
            .O(N__23659),
            .I(N__23656));
    LocalMux I__4288 (
            .O(N__23656),
            .I(\b2v_inst11.mult1_un152_sum_cry_4_s ));
    InMux I__4287 (
            .O(N__23653),
            .I(\b2v_inst11.mult1_un159_sum_cry_3 ));
    InMux I__4286 (
            .O(N__23650),
            .I(N__23647));
    LocalMux I__4285 (
            .O(N__23647),
            .I(\b2v_inst11.mult1_un152_sum_cry_5_s ));
    InMux I__4284 (
            .O(N__23644),
            .I(\b2v_inst11.mult1_un159_sum_cry_4 ));
    CascadeMux I__4283 (
            .O(N__23641),
            .I(N__23638));
    InMux I__4282 (
            .O(N__23638),
            .I(N__23635));
    LocalMux I__4281 (
            .O(N__23635),
            .I(\b2v_inst11.mult1_un152_sum_cry_6_s ));
    InMux I__4280 (
            .O(N__23632),
            .I(\b2v_inst11.mult1_un159_sum_cry_5 ));
    InMux I__4279 (
            .O(N__23629),
            .I(N__23626));
    LocalMux I__4278 (
            .O(N__23626),
            .I(\b2v_inst11.mult1_un159_sum_axb_7 ));
    InMux I__4277 (
            .O(N__23623),
            .I(\b2v_inst11.mult1_un159_sum_cry_6 ));
    CascadeMux I__4276 (
            .O(N__23620),
            .I(N__23616));
    InMux I__4275 (
            .O(N__23619),
            .I(N__23610));
    InMux I__4274 (
            .O(N__23616),
            .I(N__23603));
    InMux I__4273 (
            .O(N__23615),
            .I(N__23603));
    InMux I__4272 (
            .O(N__23614),
            .I(N__23603));
    InMux I__4271 (
            .O(N__23613),
            .I(N__23600));
    LocalMux I__4270 (
            .O(N__23610),
            .I(\b2v_inst11.mult1_un152_sum_s_8 ));
    LocalMux I__4269 (
            .O(N__23603),
            .I(\b2v_inst11.mult1_un152_sum_s_8 ));
    LocalMux I__4268 (
            .O(N__23600),
            .I(\b2v_inst11.mult1_un152_sum_s_8 ));
    CascadeMux I__4267 (
            .O(N__23593),
            .I(N__23589));
    InMux I__4266 (
            .O(N__23592),
            .I(N__23581));
    InMux I__4265 (
            .O(N__23589),
            .I(N__23581));
    InMux I__4264 (
            .O(N__23588),
            .I(N__23581));
    LocalMux I__4263 (
            .O(N__23581),
            .I(\b2v_inst11.mult1_un152_sum_i_0_8 ));
    CascadeMux I__4262 (
            .O(N__23578),
            .I(\b2v_inst36.countZ0Z_10_cascade_ ));
    InMux I__4261 (
            .O(N__23575),
            .I(N__23572));
    LocalMux I__4260 (
            .O(N__23572),
            .I(\b2v_inst36.count_1_10 ));
    CascadeMux I__4259 (
            .O(N__23569),
            .I(N__23566));
    InMux I__4258 (
            .O(N__23566),
            .I(N__23563));
    LocalMux I__4257 (
            .O(N__23563),
            .I(N__23560));
    Odrv4 I__4256 (
            .O(N__23560),
            .I(\b2v_inst11.mult1_un145_sum_i ));
    InMux I__4255 (
            .O(N__23557),
            .I(\b2v_inst11.mult1_un152_sum_cry_2 ));
    InMux I__4254 (
            .O(N__23554),
            .I(N__23551));
    LocalMux I__4253 (
            .O(N__23551),
            .I(\b2v_inst11.mult1_un145_sum_cry_3_s ));
    InMux I__4252 (
            .O(N__23548),
            .I(\b2v_inst11.mult1_un152_sum_cry_3 ));
    CascadeMux I__4251 (
            .O(N__23545),
            .I(N__23542));
    InMux I__4250 (
            .O(N__23542),
            .I(N__23539));
    LocalMux I__4249 (
            .O(N__23539),
            .I(\b2v_inst11.mult1_un145_sum_cry_4_s ));
    InMux I__4248 (
            .O(N__23536),
            .I(\b2v_inst11.mult1_un152_sum_cry_4 ));
    InMux I__4247 (
            .O(N__23533),
            .I(N__23530));
    LocalMux I__4246 (
            .O(N__23530),
            .I(\b2v_inst11.mult1_un145_sum_cry_5_s ));
    InMux I__4245 (
            .O(N__23527),
            .I(\b2v_inst11.mult1_un152_sum_cry_5 ));
    CascadeMux I__4244 (
            .O(N__23524),
            .I(N__23521));
    InMux I__4243 (
            .O(N__23521),
            .I(N__23518));
    LocalMux I__4242 (
            .O(N__23518),
            .I(N__23515));
    Odrv4 I__4241 (
            .O(N__23515),
            .I(\b2v_inst11.mult1_un145_sum_cry_6_s ));
    InMux I__4240 (
            .O(N__23512),
            .I(\b2v_inst11.mult1_un152_sum_cry_6 ));
    InMux I__4239 (
            .O(N__23509),
            .I(N__23506));
    LocalMux I__4238 (
            .O(N__23506),
            .I(\b2v_inst11.mult1_un152_sum_axb_8 ));
    InMux I__4237 (
            .O(N__23503),
            .I(\b2v_inst11.mult1_un152_sum_cry_7 ));
    CascadeMux I__4236 (
            .O(N__23500),
            .I(\b2v_inst36.count_rst_9_cascade_ ));
    CascadeMux I__4235 (
            .O(N__23497),
            .I(\b2v_inst36.countZ0Z_5_cascade_ ));
    InMux I__4234 (
            .O(N__23494),
            .I(N__23491));
    LocalMux I__4233 (
            .O(N__23491),
            .I(\b2v_inst36.count_1_5 ));
    InMux I__4232 (
            .O(N__23488),
            .I(N__23485));
    LocalMux I__4231 (
            .O(N__23485),
            .I(\b2v_inst36.count_rst_7 ));
    CascadeMux I__4230 (
            .O(N__23482),
            .I(\b2v_inst36.count_rst_6_cascade_ ));
    CascadeMux I__4229 (
            .O(N__23479),
            .I(\b2v_inst36.countZ0Z_8_cascade_ ));
    InMux I__4228 (
            .O(N__23476),
            .I(N__23473));
    LocalMux I__4227 (
            .O(N__23473),
            .I(\b2v_inst36.count_1_8 ));
    CascadeMux I__4226 (
            .O(N__23470),
            .I(\b2v_inst36.count_rst_4_cascade_ ));
    InMux I__4225 (
            .O(N__23467),
            .I(N__23463));
    InMux I__4224 (
            .O(N__23466),
            .I(N__23460));
    LocalMux I__4223 (
            .O(N__23463),
            .I(\b2v_inst11.func_state_RNI_0Z0Z_0 ));
    LocalMux I__4222 (
            .O(N__23460),
            .I(\b2v_inst11.func_state_RNI_0Z0Z_0 ));
    InMux I__4221 (
            .O(N__23455),
            .I(N__23452));
    LocalMux I__4220 (
            .O(N__23452),
            .I(\b2v_inst11.g1_1 ));
    InMux I__4219 (
            .O(N__23449),
            .I(N__23443));
    InMux I__4218 (
            .O(N__23448),
            .I(N__23443));
    LocalMux I__4217 (
            .O(N__23443),
            .I(\b2v_inst11.func_state_RNI673P9Z0Z_0 ));
    CascadeMux I__4216 (
            .O(N__23440),
            .I(N__23436));
    InMux I__4215 (
            .O(N__23439),
            .I(N__23431));
    InMux I__4214 (
            .O(N__23436),
            .I(N__23431));
    LocalMux I__4213 (
            .O(N__23431),
            .I(\b2v_inst11.func_stateZ1Z_0 ));
    CascadeMux I__4212 (
            .O(N__23428),
            .I(N__23424));
    CascadeMux I__4211 (
            .O(N__23427),
            .I(N__23419));
    InMux I__4210 (
            .O(N__23424),
            .I(N__23416));
    InMux I__4209 (
            .O(N__23423),
            .I(N__23409));
    InMux I__4208 (
            .O(N__23422),
            .I(N__23409));
    InMux I__4207 (
            .O(N__23419),
            .I(N__23406));
    LocalMux I__4206 (
            .O(N__23416),
            .I(N__23403));
    InMux I__4205 (
            .O(N__23415),
            .I(N__23398));
    InMux I__4204 (
            .O(N__23414),
            .I(N__23398));
    LocalMux I__4203 (
            .O(N__23409),
            .I(N__23395));
    LocalMux I__4202 (
            .O(N__23406),
            .I(\b2v_inst11.count_off_RNIZ0Z_9 ));
    Odrv4 I__4201 (
            .O(N__23403),
            .I(\b2v_inst11.count_off_RNIZ0Z_9 ));
    LocalMux I__4200 (
            .O(N__23398),
            .I(\b2v_inst11.count_off_RNIZ0Z_9 ));
    Odrv4 I__4199 (
            .O(N__23395),
            .I(\b2v_inst11.count_off_RNIZ0Z_9 ));
    CascadeMux I__4198 (
            .O(N__23386),
            .I(\b2v_inst11.N_335_cascade_ ));
    CascadeMux I__4197 (
            .O(N__23383),
            .I(N__23379));
    CascadeMux I__4196 (
            .O(N__23382),
            .I(N__23371));
    InMux I__4195 (
            .O(N__23379),
            .I(N__23368));
    InMux I__4194 (
            .O(N__23378),
            .I(N__23365));
    InMux I__4193 (
            .O(N__23377),
            .I(N__23360));
    InMux I__4192 (
            .O(N__23376),
            .I(N__23360));
    InMux I__4191 (
            .O(N__23375),
            .I(N__23355));
    InMux I__4190 (
            .O(N__23374),
            .I(N__23355));
    InMux I__4189 (
            .O(N__23371),
            .I(N__23352));
    LocalMux I__4188 (
            .O(N__23368),
            .I(N__23347));
    LocalMux I__4187 (
            .O(N__23365),
            .I(N__23347));
    LocalMux I__4186 (
            .O(N__23360),
            .I(N__23344));
    LocalMux I__4185 (
            .O(N__23355),
            .I(N__23333));
    LocalMux I__4184 (
            .O(N__23352),
            .I(N__23333));
    Span4Mux_s2_v I__4183 (
            .O(N__23347),
            .I(N__23333));
    Span4Mux_s2_v I__4182 (
            .O(N__23344),
            .I(N__23330));
    InMux I__4181 (
            .O(N__23343),
            .I(N__23327));
    InMux I__4180 (
            .O(N__23342),
            .I(N__23320));
    InMux I__4179 (
            .O(N__23341),
            .I(N__23320));
    InMux I__4178 (
            .O(N__23340),
            .I(N__23320));
    Span4Mux_h I__4177 (
            .O(N__23333),
            .I(N__23317));
    Odrv4 I__4176 (
            .O(N__23330),
            .I(\b2v_inst11.count_off_RNIQ1RAS1Z0Z_9 ));
    LocalMux I__4175 (
            .O(N__23327),
            .I(\b2v_inst11.count_off_RNIQ1RAS1Z0Z_9 ));
    LocalMux I__4174 (
            .O(N__23320),
            .I(\b2v_inst11.count_off_RNIQ1RAS1Z0Z_9 ));
    Odrv4 I__4173 (
            .O(N__23317),
            .I(\b2v_inst11.count_off_RNIQ1RAS1Z0Z_9 ));
    InMux I__4172 (
            .O(N__23308),
            .I(N__23305));
    LocalMux I__4171 (
            .O(N__23305),
            .I(\b2v_inst11.func_state_1_ss0_i_0_o2_0 ));
    CascadeMux I__4170 (
            .O(N__23302),
            .I(\b2v_inst36.count_rst_11_cascade_ ));
    CascadeMux I__4169 (
            .O(N__23299),
            .I(\b2v_inst36.countZ0Z_7_cascade_ ));
    InMux I__4168 (
            .O(N__23296),
            .I(N__23293));
    LocalMux I__4167 (
            .O(N__23293),
            .I(\b2v_inst36.count_1_7 ));
    InMux I__4166 (
            .O(N__23290),
            .I(N__23287));
    LocalMux I__4165 (
            .O(N__23287),
            .I(N__23281));
    CascadeMux I__4164 (
            .O(N__23286),
            .I(N__23278));
    CascadeMux I__4163 (
            .O(N__23285),
            .I(N__23275));
    InMux I__4162 (
            .O(N__23284),
            .I(N__23272));
    Span4Mux_h I__4161 (
            .O(N__23281),
            .I(N__23269));
    InMux I__4160 (
            .O(N__23278),
            .I(N__23264));
    InMux I__4159 (
            .O(N__23275),
            .I(N__23264));
    LocalMux I__4158 (
            .O(N__23272),
            .I(N__23261));
    Odrv4 I__4157 (
            .O(N__23269),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ));
    LocalMux I__4156 (
            .O(N__23264),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ));
    Odrv12 I__4155 (
            .O(N__23261),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ));
    CascadeMux I__4154 (
            .O(N__23254),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1_cascade_ ));
    InMux I__4153 (
            .O(N__23251),
            .I(N__23248));
    LocalMux I__4152 (
            .O(N__23248),
            .I(N__23245));
    Odrv12 I__4151 (
            .O(N__23245),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_4_sx ));
    InMux I__4150 (
            .O(N__23242),
            .I(N__23239));
    LocalMux I__4149 (
            .O(N__23239),
            .I(N__23235));
    InMux I__4148 (
            .O(N__23238),
            .I(N__23232));
    Sp12to4 I__4147 (
            .O(N__23235),
            .I(N__23226));
    LocalMux I__4146 (
            .O(N__23232),
            .I(N__23226));
    InMux I__4145 (
            .O(N__23231),
            .I(N__23223));
    Span12Mux_s3_v I__4144 (
            .O(N__23226),
            .I(N__23220));
    LocalMux I__4143 (
            .O(N__23223),
            .I(N__23217));
    Odrv12 I__4142 (
            .O(N__23220),
            .I(\b2v_inst11.func_state_RNI_0Z0Z_1 ));
    Odrv4 I__4141 (
            .O(N__23217),
            .I(\b2v_inst11.func_state_RNI_0Z0Z_1 ));
    InMux I__4140 (
            .O(N__23212),
            .I(N__23209));
    LocalMux I__4139 (
            .O(N__23209),
            .I(\b2v_inst11.func_state_1_m0_0_0_1 ));
    CascadeMux I__4138 (
            .O(N__23206),
            .I(N__23201));
    InMux I__4137 (
            .O(N__23205),
            .I(N__23196));
    InMux I__4136 (
            .O(N__23204),
            .I(N__23196));
    InMux I__4135 (
            .O(N__23201),
            .I(N__23193));
    LocalMux I__4134 (
            .O(N__23196),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_0 ));
    LocalMux I__4133 (
            .O(N__23193),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_0 ));
    InMux I__4132 (
            .O(N__23188),
            .I(N__23185));
    LocalMux I__4131 (
            .O(N__23185),
            .I(N__23180));
    CascadeMux I__4130 (
            .O(N__23184),
            .I(N__23177));
    InMux I__4129 (
            .O(N__23183),
            .I(N__23171));
    Span4Mux_s2_v I__4128 (
            .O(N__23180),
            .I(N__23168));
    InMux I__4127 (
            .O(N__23177),
            .I(N__23165));
    InMux I__4126 (
            .O(N__23176),
            .I(N__23162));
    InMux I__4125 (
            .O(N__23175),
            .I(N__23157));
    InMux I__4124 (
            .O(N__23174),
            .I(N__23157));
    LocalMux I__4123 (
            .O(N__23171),
            .I(N__23154));
    Odrv4 I__4122 (
            .O(N__23168),
            .I(\b2v_inst11.N_360 ));
    LocalMux I__4121 (
            .O(N__23165),
            .I(\b2v_inst11.N_360 ));
    LocalMux I__4120 (
            .O(N__23162),
            .I(\b2v_inst11.N_360 ));
    LocalMux I__4119 (
            .O(N__23157),
            .I(\b2v_inst11.N_360 ));
    Odrv4 I__4118 (
            .O(N__23154),
            .I(\b2v_inst11.N_360 ));
    InMux I__4117 (
            .O(N__23143),
            .I(N__23140));
    LocalMux I__4116 (
            .O(N__23140),
            .I(N__23137));
    Odrv12 I__4115 (
            .O(N__23137),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1 ));
    CascadeMux I__4114 (
            .O(N__23134),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_0_cascade_ ));
    CascadeMux I__4113 (
            .O(N__23131),
            .I(N__23128));
    InMux I__4112 (
            .O(N__23128),
            .I(N__23122));
    InMux I__4111 (
            .O(N__23127),
            .I(N__23122));
    LocalMux I__4110 (
            .O(N__23122),
            .I(N__23118));
    InMux I__4109 (
            .O(N__23121),
            .I(N__23115));
    Span4Mux_v I__4108 (
            .O(N__23118),
            .I(N__23103));
    LocalMux I__4107 (
            .O(N__23115),
            .I(N__23103));
    InMux I__4106 (
            .O(N__23114),
            .I(N__23100));
    InMux I__4105 (
            .O(N__23113),
            .I(N__23093));
    InMux I__4104 (
            .O(N__23112),
            .I(N__23093));
    InMux I__4103 (
            .O(N__23111),
            .I(N__23093));
    InMux I__4102 (
            .O(N__23110),
            .I(N__23090));
    InMux I__4101 (
            .O(N__23109),
            .I(N__23087));
    InMux I__4100 (
            .O(N__23108),
            .I(N__23084));
    Span4Mux_h I__4099 (
            .O(N__23103),
            .I(N__23077));
    LocalMux I__4098 (
            .O(N__23100),
            .I(N__23077));
    LocalMux I__4097 (
            .O(N__23093),
            .I(N__23077));
    LocalMux I__4096 (
            .O(N__23090),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    LocalMux I__4095 (
            .O(N__23087),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    LocalMux I__4094 (
            .O(N__23084),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    Odrv4 I__4093 (
            .O(N__23077),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    CascadeMux I__4092 (
            .O(N__23068),
            .I(\b2v_inst11.func_stateZ0Z_0_cascade_ ));
    CascadeMux I__4091 (
            .O(N__23065),
            .I(\b2v_inst11.N_3013_i_cascade_ ));
    InMux I__4090 (
            .O(N__23062),
            .I(N__23059));
    LocalMux I__4089 (
            .O(N__23059),
            .I(\b2v_inst11.N_330 ));
    CascadeMux I__4088 (
            .O(N__23056),
            .I(N__23050));
    CascadeMux I__4087 (
            .O(N__23055),
            .I(N__23047));
    InMux I__4086 (
            .O(N__23054),
            .I(N__23044));
    CascadeMux I__4085 (
            .O(N__23053),
            .I(N__23040));
    InMux I__4084 (
            .O(N__23050),
            .I(N__23037));
    InMux I__4083 (
            .O(N__23047),
            .I(N__23034));
    LocalMux I__4082 (
            .O(N__23044),
            .I(N__23031));
    InMux I__4081 (
            .O(N__23043),
            .I(N__23028));
    InMux I__4080 (
            .O(N__23040),
            .I(N__23025));
    LocalMux I__4079 (
            .O(N__23037),
            .I(N__23020));
    LocalMux I__4078 (
            .O(N__23034),
            .I(N__23020));
    Span4Mux_v I__4077 (
            .O(N__23031),
            .I(N__23017));
    LocalMux I__4076 (
            .O(N__23028),
            .I(N__23014));
    LocalMux I__4075 (
            .O(N__23025),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    Odrv4 I__4074 (
            .O(N__23020),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    Odrv4 I__4073 (
            .O(N__23017),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    Odrv12 I__4072 (
            .O(N__23014),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    CascadeMux I__4071 (
            .O(N__23005),
            .I(\b2v_inst11.dutycycle_1_0_0_cascade_ ));
    InMux I__4070 (
            .O(N__23002),
            .I(N__22999));
    LocalMux I__4069 (
            .O(N__22999),
            .I(N__22996));
    Span4Mux_h I__4068 (
            .O(N__22996),
            .I(N__22993));
    Odrv4 I__4067 (
            .O(N__22993),
            .I(\b2v_inst11.un1_dutycycle_94_cry_5_c_RNIZ0 ));
    InMux I__4066 (
            .O(N__22990),
            .I(N__22987));
    LocalMux I__4065 (
            .O(N__22987),
            .I(\b2v_inst11.g1 ));
    InMux I__4064 (
            .O(N__22984),
            .I(N__22978));
    InMux I__4063 (
            .O(N__22983),
            .I(N__22978));
    LocalMux I__4062 (
            .O(N__22978),
            .I(\b2v_inst11.dutycycle_0_6 ));
    CascadeMux I__4061 (
            .O(N__22975),
            .I(\b2v_inst11.g1_cascade_ ));
    InMux I__4060 (
            .O(N__22972),
            .I(N__22968));
    InMux I__4059 (
            .O(N__22971),
            .I(N__22965));
    LocalMux I__4058 (
            .O(N__22968),
            .I(\b2v_inst11.g1_0 ));
    LocalMux I__4057 (
            .O(N__22965),
            .I(\b2v_inst11.g1_0 ));
    InMux I__4056 (
            .O(N__22960),
            .I(N__22957));
    LocalMux I__4055 (
            .O(N__22957),
            .I(N__22954));
    Odrv4 I__4054 (
            .O(N__22954),
            .I(\b2v_inst11.dutycycle_eena ));
    InMux I__4053 (
            .O(N__22951),
            .I(N__22948));
    LocalMux I__4052 (
            .O(N__22948),
            .I(\b2v_inst11.dutycycle_1_0_0 ));
    CascadeMux I__4051 (
            .O(N__22945),
            .I(\b2v_inst11.dutycycle_eena_cascade_ ));
    InMux I__4050 (
            .O(N__22942),
            .I(N__22936));
    InMux I__4049 (
            .O(N__22941),
            .I(N__22936));
    LocalMux I__4048 (
            .O(N__22936),
            .I(\b2v_inst11.dutycycleZ1Z_0 ));
    CascadeMux I__4047 (
            .O(N__22933),
            .I(N__22930));
    InMux I__4046 (
            .O(N__22930),
            .I(N__22924));
    InMux I__4045 (
            .O(N__22929),
            .I(N__22924));
    LocalMux I__4044 (
            .O(N__22924),
            .I(N__22921));
    Span4Mux_s2_h I__4043 (
            .O(N__22921),
            .I(N__22918));
    Span4Mux_h I__4042 (
            .O(N__22918),
            .I(N__22915));
    Odrv4 I__4041 (
            .O(N__22915),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3 ));
    InMux I__4040 (
            .O(N__22912),
            .I(N__22909));
    LocalMux I__4039 (
            .O(N__22909),
            .I(\b2v_inst11.un1_clk_100khz_2_i_o3_out ));
    InMux I__4038 (
            .O(N__22906),
            .I(N__22903));
    LocalMux I__4037 (
            .O(N__22903),
            .I(\b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8 ));
    InMux I__4036 (
            .O(N__22900),
            .I(N__22897));
    LocalMux I__4035 (
            .O(N__22897),
            .I(\b2v_inst11.dutycycle_1_0_1 ));
    InMux I__4034 (
            .O(N__22894),
            .I(N__22888));
    InMux I__4033 (
            .O(N__22893),
            .I(N__22888));
    LocalMux I__4032 (
            .O(N__22888),
            .I(\b2v_inst11.dutycycleZ1Z_1 ));
    CascadeMux I__4031 (
            .O(N__22885),
            .I(\b2v_inst11.dutycycle_1_0_1_cascade_ ));
    InMux I__4030 (
            .O(N__22882),
            .I(N__22879));
    LocalMux I__4029 (
            .O(N__22879),
            .I(N__22876));
    Span4Mux_s3_v I__4028 (
            .O(N__22876),
            .I(N__22872));
    InMux I__4027 (
            .O(N__22875),
            .I(N__22869));
    Span4Mux_h I__4026 (
            .O(N__22872),
            .I(N__22866));
    LocalMux I__4025 (
            .O(N__22869),
            .I(N__22863));
    Span4Mux_h I__4024 (
            .O(N__22866),
            .I(N__22860));
    Span4Mux_h I__4023 (
            .O(N__22863),
            .I(N__22857));
    Odrv4 I__4022 (
            .O(N__22860),
            .I(\b2v_inst11.func_state_RNI_1Z0Z_0 ));
    Odrv4 I__4021 (
            .O(N__22857),
            .I(\b2v_inst11.func_state_RNI_1Z0Z_0 ));
    CascadeMux I__4020 (
            .O(N__22852),
            .I(\b2v_inst11.func_state_RNI_0Z0Z_1_cascade_ ));
    CascadeMux I__4019 (
            .O(N__22849),
            .I(\b2v_inst11.un1_func_state25_4_i_a2_1_cascade_ ));
    InMux I__4018 (
            .O(N__22846),
            .I(N__22843));
    LocalMux I__4017 (
            .O(N__22843),
            .I(N__22840));
    Span4Mux_s2_h I__4016 (
            .O(N__22840),
            .I(N__22837));
    Span4Mux_h I__4015 (
            .O(N__22837),
            .I(N__22834));
    Odrv4 I__4014 (
            .O(N__22834),
            .I(\b2v_inst11.N_321 ));
    InMux I__4013 (
            .O(N__22831),
            .I(N__22828));
    LocalMux I__4012 (
            .O(N__22828),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_3 ));
    InMux I__4011 (
            .O(N__22825),
            .I(N__22819));
    InMux I__4010 (
            .O(N__22824),
            .I(N__22819));
    LocalMux I__4009 (
            .O(N__22819),
            .I(N__22816));
    Odrv4 I__4008 (
            .O(N__22816),
            .I(\b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8 ));
    CascadeMux I__4007 (
            .O(N__22813),
            .I(N__22810));
    InMux I__4006 (
            .O(N__22810),
            .I(N__22804));
    InMux I__4005 (
            .O(N__22809),
            .I(N__22804));
    LocalMux I__4004 (
            .O(N__22804),
            .I(\b2v_inst11.dutycycle_e_1_3 ));
    CascadeMux I__4003 (
            .O(N__22801),
            .I(N__22797));
    InMux I__4002 (
            .O(N__22800),
            .I(N__22792));
    InMux I__4001 (
            .O(N__22797),
            .I(N__22792));
    LocalMux I__4000 (
            .O(N__22792),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    CascadeMux I__3999 (
            .O(N__22789),
            .I(\b2v_inst11.dutycycleZ0Z_6_cascade_ ));
    InMux I__3998 (
            .O(N__22786),
            .I(N__22780));
    InMux I__3997 (
            .O(N__22785),
            .I(N__22768));
    InMux I__3996 (
            .O(N__22784),
            .I(N__22765));
    CascadeMux I__3995 (
            .O(N__22783),
            .I(N__22758));
    LocalMux I__3994 (
            .O(N__22780),
            .I(N__22755));
    InMux I__3993 (
            .O(N__22779),
            .I(N__22750));
    InMux I__3992 (
            .O(N__22778),
            .I(N__22750));
    InMux I__3991 (
            .O(N__22777),
            .I(N__22743));
    InMux I__3990 (
            .O(N__22776),
            .I(N__22743));
    InMux I__3989 (
            .O(N__22775),
            .I(N__22743));
    InMux I__3988 (
            .O(N__22774),
            .I(N__22738));
    InMux I__3987 (
            .O(N__22773),
            .I(N__22738));
    InMux I__3986 (
            .O(N__22772),
            .I(N__22735));
    CascadeMux I__3985 (
            .O(N__22771),
            .I(N__22730));
    LocalMux I__3984 (
            .O(N__22768),
            .I(N__22722));
    LocalMux I__3983 (
            .O(N__22765),
            .I(N__22719));
    InMux I__3982 (
            .O(N__22764),
            .I(N__22716));
    InMux I__3981 (
            .O(N__22763),
            .I(N__22711));
    InMux I__3980 (
            .O(N__22762),
            .I(N__22711));
    InMux I__3979 (
            .O(N__22761),
            .I(N__22708));
    InMux I__3978 (
            .O(N__22758),
            .I(N__22705));
    Span4Mux_h I__3977 (
            .O(N__22755),
            .I(N__22702));
    LocalMux I__3976 (
            .O(N__22750),
            .I(N__22699));
    LocalMux I__3975 (
            .O(N__22743),
            .I(N__22692));
    LocalMux I__3974 (
            .O(N__22738),
            .I(N__22692));
    LocalMux I__3973 (
            .O(N__22735),
            .I(N__22692));
    InMux I__3972 (
            .O(N__22734),
            .I(N__22681));
    InMux I__3971 (
            .O(N__22733),
            .I(N__22681));
    InMux I__3970 (
            .O(N__22730),
            .I(N__22681));
    InMux I__3969 (
            .O(N__22729),
            .I(N__22681));
    InMux I__3968 (
            .O(N__22728),
            .I(N__22681));
    InMux I__3967 (
            .O(N__22727),
            .I(N__22674));
    InMux I__3966 (
            .O(N__22726),
            .I(N__22674));
    InMux I__3965 (
            .O(N__22725),
            .I(N__22674));
    Span4Mux_h I__3964 (
            .O(N__22722),
            .I(N__22669));
    Span4Mux_h I__3963 (
            .O(N__22719),
            .I(N__22669));
    LocalMux I__3962 (
            .O(N__22716),
            .I(N__22664));
    LocalMux I__3961 (
            .O(N__22711),
            .I(N__22664));
    LocalMux I__3960 (
            .O(N__22708),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__3959 (
            .O(N__22705),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    Odrv4 I__3958 (
            .O(N__22702),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    Odrv4 I__3957 (
            .O(N__22699),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    Odrv4 I__3956 (
            .O(N__22692),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__3955 (
            .O(N__22681),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__3954 (
            .O(N__22674),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    Odrv4 I__3953 (
            .O(N__22669),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    Odrv12 I__3952 (
            .O(N__22664),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    InMux I__3951 (
            .O(N__22645),
            .I(N__22642));
    LocalMux I__3950 (
            .O(N__22642),
            .I(N__22639));
    Odrv4 I__3949 (
            .O(N__22639),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_3 ));
    CascadeMux I__3948 (
            .O(N__22636),
            .I(\b2v_inst11.func_state_RNINJ641_0Z0Z_1_cascade_ ));
    CascadeMux I__3947 (
            .O(N__22633),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1_cascade_ ));
    InMux I__3946 (
            .O(N__22630),
            .I(N__22627));
    LocalMux I__3945 (
            .O(N__22627),
            .I(\b2v_inst11.g0_2_3 ));
    InMux I__3944 (
            .O(N__22624),
            .I(N__22621));
    LocalMux I__3943 (
            .O(N__22621),
            .I(N__22618));
    Odrv4 I__3942 (
            .O(N__22618),
            .I(\b2v_inst11.g0_2_2 ));
    CascadeMux I__3941 (
            .O(N__22615),
            .I(N__22612));
    InMux I__3940 (
            .O(N__22612),
            .I(N__22609));
    LocalMux I__3939 (
            .O(N__22609),
            .I(N__22606));
    Odrv4 I__3938 (
            .O(N__22606),
            .I(\b2v_inst11.g0_1_1_0 ));
    CascadeMux I__3937 (
            .O(N__22603),
            .I(N__22600));
    InMux I__3936 (
            .O(N__22600),
            .I(N__22597));
    LocalMux I__3935 (
            .O(N__22597),
            .I(N__22594));
    Span4Mux_s3_v I__3934 (
            .O(N__22594),
            .I(N__22589));
    InMux I__3933 (
            .O(N__22593),
            .I(N__22581));
    InMux I__3932 (
            .O(N__22592),
            .I(N__22578));
    Span4Mux_h I__3931 (
            .O(N__22589),
            .I(N__22574));
    InMux I__3930 (
            .O(N__22588),
            .I(N__22567));
    InMux I__3929 (
            .O(N__22587),
            .I(N__22567));
    InMux I__3928 (
            .O(N__22586),
            .I(N__22567));
    InMux I__3927 (
            .O(N__22585),
            .I(N__22562));
    InMux I__3926 (
            .O(N__22584),
            .I(N__22562));
    LocalMux I__3925 (
            .O(N__22581),
            .I(N__22557));
    LocalMux I__3924 (
            .O(N__22578),
            .I(N__22557));
    CascadeMux I__3923 (
            .O(N__22577),
            .I(N__22554));
    Span4Mux_v I__3922 (
            .O(N__22574),
            .I(N__22550));
    LocalMux I__3921 (
            .O(N__22567),
            .I(N__22547));
    LocalMux I__3920 (
            .O(N__22562),
            .I(N__22542));
    Span4Mux_h I__3919 (
            .O(N__22557),
            .I(N__22542));
    InMux I__3918 (
            .O(N__22554),
            .I(N__22537));
    InMux I__3917 (
            .O(N__22553),
            .I(N__22537));
    Odrv4 I__3916 (
            .O(N__22550),
            .I(\b2v_inst11.func_state_RNIJU083Z0Z_0 ));
    Odrv12 I__3915 (
            .O(N__22547),
            .I(\b2v_inst11.func_state_RNIJU083Z0Z_0 ));
    Odrv4 I__3914 (
            .O(N__22542),
            .I(\b2v_inst11.func_state_RNIJU083Z0Z_0 ));
    LocalMux I__3913 (
            .O(N__22537),
            .I(\b2v_inst11.func_state_RNIJU083Z0Z_0 ));
    CascadeMux I__3912 (
            .O(N__22528),
            .I(\b2v_inst11.un1_clk_100khz_43_and_i_o2_0_0_1_cascade_ ));
    InMux I__3911 (
            .O(N__22525),
            .I(N__22522));
    LocalMux I__3910 (
            .O(N__22522),
            .I(N__22519));
    Span4Mux_h I__3909 (
            .O(N__22519),
            .I(N__22516));
    Odrv4 I__3908 (
            .O(N__22516),
            .I(\b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJTZ0Z69 ));
    InMux I__3907 (
            .O(N__22513),
            .I(N__22510));
    LocalMux I__3906 (
            .O(N__22510),
            .I(\b2v_inst11.dutycycle_RNI4I3C2Z0Z_10 ));
    CascadeMux I__3905 (
            .O(N__22507),
            .I(\b2v_inst11.dutycycle_RNI4I3C2Z0Z_10_cascade_ ));
    InMux I__3904 (
            .O(N__22504),
            .I(N__22501));
    LocalMux I__3903 (
            .O(N__22501),
            .I(\b2v_inst11.dutycycle_RNIAI7C4Z0Z_10 ));
    CascadeMux I__3902 (
            .O(N__22498),
            .I(N__22494));
    InMux I__3901 (
            .O(N__22497),
            .I(N__22486));
    InMux I__3900 (
            .O(N__22494),
            .I(N__22486));
    InMux I__3899 (
            .O(N__22493),
            .I(N__22486));
    LocalMux I__3898 (
            .O(N__22486),
            .I(\b2v_inst11.dutycycleZ1Z_10 ));
    CascadeMux I__3897 (
            .O(N__22483),
            .I(N__22480));
    InMux I__3896 (
            .O(N__22480),
            .I(N__22477));
    LocalMux I__3895 (
            .O(N__22477),
            .I(N__22474));
    Span4Mux_h I__3894 (
            .O(N__22474),
            .I(N__22471));
    Odrv4 I__3893 (
            .O(N__22471),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_5 ));
    CascadeMux I__3892 (
            .O(N__22468),
            .I(\b2v_inst11.d_i3_mux_cascade_ ));
    InMux I__3891 (
            .O(N__22465),
            .I(N__22462));
    LocalMux I__3890 (
            .O(N__22462),
            .I(N__22459));
    Span4Mux_h I__3889 (
            .O(N__22459),
            .I(N__22456));
    Odrv4 I__3888 (
            .O(N__22456),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_5 ));
    CascadeMux I__3887 (
            .O(N__22453),
            .I(N__22450));
    InMux I__3886 (
            .O(N__22450),
            .I(N__22447));
    LocalMux I__3885 (
            .O(N__22447),
            .I(N__22443));
    InMux I__3884 (
            .O(N__22446),
            .I(N__22440));
    Span4Mux_h I__3883 (
            .O(N__22443),
            .I(N__22437));
    LocalMux I__3882 (
            .O(N__22440),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_3 ));
    Odrv4 I__3881 (
            .O(N__22437),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_3 ));
    InMux I__3880 (
            .O(N__22432),
            .I(N__22429));
    LocalMux I__3879 (
            .O(N__22429),
            .I(\b2v_inst11.curr_state_0_0 ));
    InMux I__3878 (
            .O(N__22426),
            .I(N__22423));
    LocalMux I__3877 (
            .O(N__22423),
            .I(\b2v_inst11.curr_state_3_0 ));
    CascadeMux I__3876 (
            .O(N__22420),
            .I(\b2v_inst11.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__3875 (
            .O(N__22417),
            .I(\b2v_inst11.count_0_sqmuxa_i_cascade_ ));
    InMux I__3874 (
            .O(N__22414),
            .I(N__22411));
    LocalMux I__3873 (
            .O(N__22411),
            .I(N__22408));
    Span4Mux_v I__3872 (
            .O(N__22408),
            .I(N__22405));
    Odrv4 I__3871 (
            .O(N__22405),
            .I(\b2v_inst11.N_349 ));
    CascadeMux I__3870 (
            .O(N__22402),
            .I(N__22397));
    InMux I__3869 (
            .O(N__22401),
            .I(N__22393));
    InMux I__3868 (
            .O(N__22400),
            .I(N__22386));
    InMux I__3867 (
            .O(N__22397),
            .I(N__22386));
    InMux I__3866 (
            .O(N__22396),
            .I(N__22386));
    LocalMux I__3865 (
            .O(N__22393),
            .I(N__22383));
    LocalMux I__3864 (
            .O(N__22386),
            .I(N__22380));
    Span4Mux_h I__3863 (
            .O(N__22383),
            .I(N__22377));
    Span4Mux_v I__3862 (
            .O(N__22380),
            .I(N__22374));
    Span4Mux_h I__3861 (
            .O(N__22377),
            .I(N__22371));
    Odrv4 I__3860 (
            .O(N__22374),
            .I(\b2v_inst11.un1_clk_100khz_32_and_i_o2_0_0_1 ));
    Odrv4 I__3859 (
            .O(N__22371),
            .I(\b2v_inst11.un1_clk_100khz_32_and_i_o2_0_0_1 ));
    CascadeMux I__3858 (
            .O(N__22366),
            .I(\b2v_inst11.dutycycle_RNIAI7C4Z0Z_10_cascade_ ));
    CascadeMux I__3857 (
            .O(N__22363),
            .I(N__22356));
    CascadeMux I__3856 (
            .O(N__22362),
            .I(N__22351));
    InMux I__3855 (
            .O(N__22361),
            .I(N__22342));
    InMux I__3854 (
            .O(N__22360),
            .I(N__22337));
    InMux I__3853 (
            .O(N__22359),
            .I(N__22337));
    InMux I__3852 (
            .O(N__22356),
            .I(N__22334));
    InMux I__3851 (
            .O(N__22355),
            .I(N__22331));
    InMux I__3850 (
            .O(N__22354),
            .I(N__22324));
    InMux I__3849 (
            .O(N__22351),
            .I(N__22324));
    InMux I__3848 (
            .O(N__22350),
            .I(N__22324));
    InMux I__3847 (
            .O(N__22349),
            .I(N__22321));
    InMux I__3846 (
            .O(N__22348),
            .I(N__22318));
    InMux I__3845 (
            .O(N__22347),
            .I(N__22311));
    InMux I__3844 (
            .O(N__22346),
            .I(N__22311));
    InMux I__3843 (
            .O(N__22345),
            .I(N__22311));
    LocalMux I__3842 (
            .O(N__22342),
            .I(N__22305));
    LocalMux I__3841 (
            .O(N__22337),
            .I(N__22302));
    LocalMux I__3840 (
            .O(N__22334),
            .I(N__22295));
    LocalMux I__3839 (
            .O(N__22331),
            .I(N__22295));
    LocalMux I__3838 (
            .O(N__22324),
            .I(N__22295));
    LocalMux I__3837 (
            .O(N__22321),
            .I(N__22288));
    LocalMux I__3836 (
            .O(N__22318),
            .I(N__22288));
    LocalMux I__3835 (
            .O(N__22311),
            .I(N__22288));
    InMux I__3834 (
            .O(N__22310),
            .I(N__22284));
    InMux I__3833 (
            .O(N__22309),
            .I(N__22279));
    InMux I__3832 (
            .O(N__22308),
            .I(N__22279));
    Span4Mux_h I__3831 (
            .O(N__22305),
            .I(N__22276));
    Span4Mux_h I__3830 (
            .O(N__22302),
            .I(N__22269));
    Span4Mux_v I__3829 (
            .O(N__22295),
            .I(N__22269));
    Span4Mux_v I__3828 (
            .O(N__22288),
            .I(N__22269));
    InMux I__3827 (
            .O(N__22287),
            .I(N__22266));
    LocalMux I__3826 (
            .O(N__22284),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    LocalMux I__3825 (
            .O(N__22279),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    Odrv4 I__3824 (
            .O(N__22276),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    Odrv4 I__3823 (
            .O(N__22269),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    LocalMux I__3822 (
            .O(N__22266),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    InMux I__3821 (
            .O(N__22255),
            .I(N__22250));
    InMux I__3820 (
            .O(N__22254),
            .I(N__22245));
    InMux I__3819 (
            .O(N__22253),
            .I(N__22245));
    LocalMux I__3818 (
            .O(N__22250),
            .I(N__22233));
    LocalMux I__3817 (
            .O(N__22245),
            .I(N__22233));
    InMux I__3816 (
            .O(N__22244),
            .I(N__22228));
    InMux I__3815 (
            .O(N__22243),
            .I(N__22228));
    InMux I__3814 (
            .O(N__22242),
            .I(N__22224));
    InMux I__3813 (
            .O(N__22241),
            .I(N__22221));
    InMux I__3812 (
            .O(N__22240),
            .I(N__22216));
    InMux I__3811 (
            .O(N__22239),
            .I(N__22216));
    InMux I__3810 (
            .O(N__22238),
            .I(N__22213));
    Span4Mux_v I__3809 (
            .O(N__22233),
            .I(N__22210));
    LocalMux I__3808 (
            .O(N__22228),
            .I(N__22207));
    InMux I__3807 (
            .O(N__22227),
            .I(N__22204));
    LocalMux I__3806 (
            .O(N__22224),
            .I(N__22199));
    LocalMux I__3805 (
            .O(N__22221),
            .I(N__22199));
    LocalMux I__3804 (
            .O(N__22216),
            .I(N__22194));
    LocalMux I__3803 (
            .O(N__22213),
            .I(N__22194));
    Span4Mux_v I__3802 (
            .O(N__22210),
            .I(N__22191));
    Span4Mux_v I__3801 (
            .O(N__22207),
            .I(N__22188));
    LocalMux I__3800 (
            .O(N__22204),
            .I(N__22181));
    Span4Mux_v I__3799 (
            .O(N__22199),
            .I(N__22181));
    Span4Mux_h I__3798 (
            .O(N__22194),
            .I(N__22181));
    Odrv4 I__3797 (
            .O(N__22191),
            .I(\b2v_inst11.N_418 ));
    Odrv4 I__3796 (
            .O(N__22188),
            .I(\b2v_inst11.N_418 ));
    Odrv4 I__3795 (
            .O(N__22181),
            .I(\b2v_inst11.N_418 ));
    CascadeMux I__3794 (
            .O(N__22174),
            .I(N__22171));
    InMux I__3793 (
            .O(N__22171),
            .I(N__22168));
    LocalMux I__3792 (
            .O(N__22168),
            .I(\b2v_inst11.mult1_un61_sum_i_8 ));
    InMux I__3791 (
            .O(N__22165),
            .I(N__22162));
    LocalMux I__3790 (
            .O(N__22162),
            .I(\b2v_inst11.N_5661_i ));
    InMux I__3789 (
            .O(N__22159),
            .I(bfn_7_7_0_));
    InMux I__3788 (
            .O(N__22156),
            .I(N__22153));
    LocalMux I__3787 (
            .O(N__22153),
            .I(N__22150));
    Odrv4 I__3786 (
            .O(N__22150),
            .I(\b2v_inst36.curr_state_RNI8TT2Z0Z_0 ));
    CascadeMux I__3785 (
            .O(N__22147),
            .I(\b2v_inst11.pwm_out_en_cascade_ ));
    IoInMux I__3784 (
            .O(N__22144),
            .I(N__22141));
    LocalMux I__3783 (
            .O(N__22141),
            .I(N__22138));
    Span4Mux_s0_v I__3782 (
            .O(N__22138),
            .I(N__22135));
    Span4Mux_v I__3781 (
            .O(N__22135),
            .I(N__22132));
    Span4Mux_v I__3780 (
            .O(N__22132),
            .I(N__22129));
    Odrv4 I__3779 (
            .O(N__22129),
            .I(PWRBTN_LED_c));
    InMux I__3778 (
            .O(N__22126),
            .I(N__22123));
    LocalMux I__3777 (
            .O(N__22123),
            .I(\b2v_inst11.pwm_out_1_sqmuxa_0 ));
    InMux I__3776 (
            .O(N__22120),
            .I(N__22117));
    LocalMux I__3775 (
            .O(N__22117),
            .I(\b2v_inst11.N_5653_i ));
    CascadeMux I__3774 (
            .O(N__22114),
            .I(N__22111));
    InMux I__3773 (
            .O(N__22111),
            .I(N__22108));
    LocalMux I__3772 (
            .O(N__22108),
            .I(\b2v_inst11.un85_clk_100khz_8 ));
    InMux I__3771 (
            .O(N__22105),
            .I(N__22102));
    LocalMux I__3770 (
            .O(N__22102),
            .I(\b2v_inst11.N_5654_i ));
    InMux I__3769 (
            .O(N__22099),
            .I(N__22096));
    LocalMux I__3768 (
            .O(N__22096),
            .I(N__22093));
    Span4Mux_v I__3767 (
            .O(N__22093),
            .I(N__22090));
    Odrv4 I__3766 (
            .O(N__22090),
            .I(\b2v_inst11.un85_clk_100khz_9 ));
    CascadeMux I__3765 (
            .O(N__22087),
            .I(N__22084));
    InMux I__3764 (
            .O(N__22084),
            .I(N__22081));
    LocalMux I__3763 (
            .O(N__22081),
            .I(\b2v_inst11.N_5655_i ));
    CascadeMux I__3762 (
            .O(N__22078),
            .I(N__22075));
    InMux I__3761 (
            .O(N__22075),
            .I(N__22072));
    LocalMux I__3760 (
            .O(N__22072),
            .I(\b2v_inst11.un85_clk_100khz_10 ));
    InMux I__3759 (
            .O(N__22069),
            .I(N__22066));
    LocalMux I__3758 (
            .O(N__22066),
            .I(\b2v_inst11.N_5656_i ));
    InMux I__3757 (
            .O(N__22063),
            .I(N__22060));
    LocalMux I__3756 (
            .O(N__22060),
            .I(N__22057));
    Span4Mux_v I__3755 (
            .O(N__22057),
            .I(N__22054));
    Odrv4 I__3754 (
            .O(N__22054),
            .I(\b2v_inst11.un85_clk_100khz_11 ));
    CascadeMux I__3753 (
            .O(N__22051),
            .I(N__22048));
    InMux I__3752 (
            .O(N__22048),
            .I(N__22045));
    LocalMux I__3751 (
            .O(N__22045),
            .I(\b2v_inst11.N_5657_i ));
    CascadeMux I__3750 (
            .O(N__22042),
            .I(N__22039));
    InMux I__3749 (
            .O(N__22039),
            .I(N__22036));
    LocalMux I__3748 (
            .O(N__22036),
            .I(N__22033));
    Odrv4 I__3747 (
            .O(N__22033),
            .I(\b2v_inst11.un85_clk_100khz_12 ));
    InMux I__3746 (
            .O(N__22030),
            .I(N__22027));
    LocalMux I__3745 (
            .O(N__22027),
            .I(\b2v_inst11.N_5658_i ));
    InMux I__3744 (
            .O(N__22024),
            .I(N__22021));
    LocalMux I__3743 (
            .O(N__22021),
            .I(\b2v_inst11.un85_clk_100khz_13 ));
    CascadeMux I__3742 (
            .O(N__22018),
            .I(N__22015));
    InMux I__3741 (
            .O(N__22015),
            .I(N__22012));
    LocalMux I__3740 (
            .O(N__22012),
            .I(\b2v_inst11.N_5659_i ));
    CascadeMux I__3739 (
            .O(N__22009),
            .I(N__22006));
    InMux I__3738 (
            .O(N__22006),
            .I(N__22003));
    LocalMux I__3737 (
            .O(N__22003),
            .I(\b2v_inst11.un85_clk_100khz_14 ));
    InMux I__3736 (
            .O(N__22000),
            .I(N__21997));
    LocalMux I__3735 (
            .O(N__21997),
            .I(\b2v_inst11.N_5660_i ));
    InMux I__3734 (
            .O(N__21994),
            .I(N__21991));
    LocalMux I__3733 (
            .O(N__21991),
            .I(\b2v_inst11.mult1_un131_sum_i ));
    CascadeMux I__3732 (
            .O(N__21988),
            .I(N__21985));
    InMux I__3731 (
            .O(N__21985),
            .I(N__21982));
    LocalMux I__3730 (
            .O(N__21982),
            .I(N__21979));
    Span4Mux_h I__3729 (
            .O(N__21979),
            .I(N__21976));
    Odrv4 I__3728 (
            .O(N__21976),
            .I(\b2v_inst11.un1_count_cry_0_i ));
    CascadeMux I__3727 (
            .O(N__21973),
            .I(N__21970));
    InMux I__3726 (
            .O(N__21970),
            .I(N__21967));
    LocalMux I__3725 (
            .O(N__21967),
            .I(\b2v_inst11.un85_clk_100khz_1 ));
    InMux I__3724 (
            .O(N__21964),
            .I(N__21961));
    LocalMux I__3723 (
            .O(N__21961),
            .I(\b2v_inst11.N_5647_i ));
    InMux I__3722 (
            .O(N__21958),
            .I(N__21955));
    LocalMux I__3721 (
            .O(N__21955),
            .I(\b2v_inst11.un85_clk_100khz_2 ));
    CascadeMux I__3720 (
            .O(N__21952),
            .I(N__21949));
    InMux I__3719 (
            .O(N__21949),
            .I(N__21946));
    LocalMux I__3718 (
            .O(N__21946),
            .I(\b2v_inst11.N_5648_i ));
    InMux I__3717 (
            .O(N__21943),
            .I(N__21940));
    LocalMux I__3716 (
            .O(N__21940),
            .I(\b2v_inst11.un85_clk_100khz_3 ));
    CascadeMux I__3715 (
            .O(N__21937),
            .I(N__21934));
    InMux I__3714 (
            .O(N__21934),
            .I(N__21931));
    LocalMux I__3713 (
            .O(N__21931),
            .I(N__21928));
    Odrv12 I__3712 (
            .O(N__21928),
            .I(\b2v_inst11.N_5649_i ));
    CascadeMux I__3711 (
            .O(N__21925),
            .I(N__21922));
    InMux I__3710 (
            .O(N__21922),
            .I(N__21919));
    LocalMux I__3709 (
            .O(N__21919),
            .I(N__21916));
    Odrv4 I__3708 (
            .O(N__21916),
            .I(\b2v_inst11.un85_clk_100khz_4 ));
    InMux I__3707 (
            .O(N__21913),
            .I(N__21910));
    LocalMux I__3706 (
            .O(N__21910),
            .I(\b2v_inst11.N_5650_i ));
    CascadeMux I__3705 (
            .O(N__21907),
            .I(N__21904));
    InMux I__3704 (
            .O(N__21904),
            .I(N__21901));
    LocalMux I__3703 (
            .O(N__21901),
            .I(\b2v_inst11.un85_clk_100khz_5 ));
    InMux I__3702 (
            .O(N__21898),
            .I(N__21895));
    LocalMux I__3701 (
            .O(N__21895),
            .I(\b2v_inst11.N_5651_i ));
    InMux I__3700 (
            .O(N__21892),
            .I(N__21889));
    LocalMux I__3699 (
            .O(N__21889),
            .I(\b2v_inst11.un85_clk_100khz_6 ));
    CascadeMux I__3698 (
            .O(N__21886),
            .I(N__21883));
    InMux I__3697 (
            .O(N__21883),
            .I(N__21880));
    LocalMux I__3696 (
            .O(N__21880),
            .I(\b2v_inst11.N_5652_i ));
    CascadeMux I__3695 (
            .O(N__21877),
            .I(N__21874));
    InMux I__3694 (
            .O(N__21874),
            .I(N__21871));
    LocalMux I__3693 (
            .O(N__21871),
            .I(\b2v_inst11.un85_clk_100khz_7 ));
    InMux I__3692 (
            .O(N__21868),
            .I(N__21865));
    LocalMux I__3691 (
            .O(N__21865),
            .I(\b2v_inst11.mult1_un138_sum_axb_8 ));
    InMux I__3690 (
            .O(N__21862),
            .I(\b2v_inst11.mult1_un138_sum_cry_7 ));
    CascadeMux I__3689 (
            .O(N__21859),
            .I(N__21856));
    InMux I__3688 (
            .O(N__21856),
            .I(N__21846));
    InMux I__3687 (
            .O(N__21855),
            .I(N__21846));
    InMux I__3686 (
            .O(N__21854),
            .I(N__21846));
    InMux I__3685 (
            .O(N__21853),
            .I(N__21843));
    LocalMux I__3684 (
            .O(N__21846),
            .I(\b2v_inst11.mult1_un138_sum_s_8 ));
    LocalMux I__3683 (
            .O(N__21843),
            .I(\b2v_inst11.mult1_un138_sum_s_8 ));
    CascadeMux I__3682 (
            .O(N__21838),
            .I(\b2v_inst11.mult1_un138_sum_s_8_cascade_ ));
    InMux I__3681 (
            .O(N__21835),
            .I(N__21832));
    LocalMux I__3680 (
            .O(N__21832),
            .I(N__21828));
    CascadeMux I__3679 (
            .O(N__21831),
            .I(N__21825));
    Span4Mux_v I__3678 (
            .O(N__21828),
            .I(N__21819));
    InMux I__3677 (
            .O(N__21825),
            .I(N__21812));
    InMux I__3676 (
            .O(N__21824),
            .I(N__21812));
    InMux I__3675 (
            .O(N__21823),
            .I(N__21812));
    InMux I__3674 (
            .O(N__21822),
            .I(N__21809));
    Odrv4 I__3673 (
            .O(N__21819),
            .I(\b2v_inst11.mult1_un82_sum_s_8 ));
    LocalMux I__3672 (
            .O(N__21812),
            .I(\b2v_inst11.mult1_un82_sum_s_8 ));
    LocalMux I__3671 (
            .O(N__21809),
            .I(\b2v_inst11.mult1_un82_sum_s_8 ));
    CascadeMux I__3670 (
            .O(N__21802),
            .I(N__21798));
    InMux I__3669 (
            .O(N__21801),
            .I(N__21793));
    InMux I__3668 (
            .O(N__21798),
            .I(N__21788));
    InMux I__3667 (
            .O(N__21797),
            .I(N__21788));
    InMux I__3666 (
            .O(N__21796),
            .I(N__21785));
    LocalMux I__3665 (
            .O(N__21793),
            .I(\b2v_inst11.mult1_un131_sum_s_8 ));
    LocalMux I__3664 (
            .O(N__21788),
            .I(\b2v_inst11.mult1_un131_sum_s_8 ));
    LocalMux I__3663 (
            .O(N__21785),
            .I(\b2v_inst11.mult1_un131_sum_s_8 ));
    InMux I__3662 (
            .O(N__21778),
            .I(N__21775));
    LocalMux I__3661 (
            .O(N__21775),
            .I(N__21771));
    InMux I__3660 (
            .O(N__21774),
            .I(N__21768));
    Span4Mux_s2_v I__3659 (
            .O(N__21771),
            .I(N__21763));
    LocalMux I__3658 (
            .O(N__21768),
            .I(N__21763));
    Span4Mux_v I__3657 (
            .O(N__21763),
            .I(N__21760));
    Odrv4 I__3656 (
            .O(N__21760),
            .I(\b2v_inst11.mult1_un138_sum ));
    CascadeMux I__3655 (
            .O(N__21757),
            .I(N__21754));
    InMux I__3654 (
            .O(N__21754),
            .I(N__21751));
    LocalMux I__3653 (
            .O(N__21751),
            .I(N__21748));
    Odrv4 I__3652 (
            .O(N__21748),
            .I(\b2v_inst11.mult1_un138_sum_i ));
    InMux I__3651 (
            .O(N__21745),
            .I(N__21741));
    InMux I__3650 (
            .O(N__21744),
            .I(N__21738));
    LocalMux I__3649 (
            .O(N__21741),
            .I(N__21735));
    LocalMux I__3648 (
            .O(N__21738),
            .I(N__21732));
    Span4Mux_h I__3647 (
            .O(N__21735),
            .I(N__21729));
    Span4Mux_h I__3646 (
            .O(N__21732),
            .I(N__21726));
    Odrv4 I__3645 (
            .O(N__21729),
            .I(\b2v_inst11.mult1_un131_sum ));
    Odrv4 I__3644 (
            .O(N__21726),
            .I(\b2v_inst11.mult1_un131_sum ));
    InMux I__3643 (
            .O(N__21721),
            .I(\b2v_inst11.mult1_un145_sum_cry_7 ));
    CascadeMux I__3642 (
            .O(N__21718),
            .I(N__21714));
    InMux I__3641 (
            .O(N__21717),
            .I(N__21706));
    InMux I__3640 (
            .O(N__21714),
            .I(N__21706));
    InMux I__3639 (
            .O(N__21713),
            .I(N__21706));
    LocalMux I__3638 (
            .O(N__21706),
            .I(\b2v_inst11.mult1_un138_sum_i_0_8 ));
    InMux I__3637 (
            .O(N__21703),
            .I(N__21700));
    LocalMux I__3636 (
            .O(N__21700),
            .I(\b2v_inst11.mult1_un138_sum_cry_3_s ));
    InMux I__3635 (
            .O(N__21697),
            .I(\b2v_inst11.mult1_un138_sum_cry_2 ));
    CascadeMux I__3634 (
            .O(N__21694),
            .I(N__21691));
    InMux I__3633 (
            .O(N__21691),
            .I(N__21688));
    LocalMux I__3632 (
            .O(N__21688),
            .I(\b2v_inst11.mult1_un131_sum_cry_3_s ));
    CascadeMux I__3631 (
            .O(N__21685),
            .I(N__21682));
    InMux I__3630 (
            .O(N__21682),
            .I(N__21679));
    LocalMux I__3629 (
            .O(N__21679),
            .I(\b2v_inst11.mult1_un138_sum_cry_4_s ));
    InMux I__3628 (
            .O(N__21676),
            .I(\b2v_inst11.mult1_un138_sum_cry_3 ));
    CascadeMux I__3627 (
            .O(N__21673),
            .I(N__21670));
    InMux I__3626 (
            .O(N__21670),
            .I(N__21667));
    LocalMux I__3625 (
            .O(N__21667),
            .I(N__21664));
    Odrv4 I__3624 (
            .O(N__21664),
            .I(\b2v_inst11.mult1_un131_sum_cry_4_s ));
    InMux I__3623 (
            .O(N__21661),
            .I(N__21658));
    LocalMux I__3622 (
            .O(N__21658),
            .I(\b2v_inst11.mult1_un138_sum_cry_5_s ));
    InMux I__3621 (
            .O(N__21655),
            .I(\b2v_inst11.mult1_un138_sum_cry_4 ));
    InMux I__3620 (
            .O(N__21652),
            .I(N__21649));
    LocalMux I__3619 (
            .O(N__21649),
            .I(\b2v_inst11.mult1_un131_sum_cry_5_s ));
    CascadeMux I__3618 (
            .O(N__21646),
            .I(N__21643));
    InMux I__3617 (
            .O(N__21643),
            .I(N__21640));
    LocalMux I__3616 (
            .O(N__21640),
            .I(\b2v_inst11.mult1_un138_sum_cry_6_s ));
    InMux I__3615 (
            .O(N__21637),
            .I(\b2v_inst11.mult1_un138_sum_cry_5 ));
    InMux I__3614 (
            .O(N__21634),
            .I(N__21631));
    LocalMux I__3613 (
            .O(N__21631),
            .I(\b2v_inst11.mult1_un131_sum_cry_6_s ));
    CascadeMux I__3612 (
            .O(N__21628),
            .I(N__21624));
    CascadeMux I__3611 (
            .O(N__21627),
            .I(N__21620));
    InMux I__3610 (
            .O(N__21624),
            .I(N__21613));
    InMux I__3609 (
            .O(N__21623),
            .I(N__21613));
    InMux I__3608 (
            .O(N__21620),
            .I(N__21613));
    LocalMux I__3607 (
            .O(N__21613),
            .I(\b2v_inst11.mult1_un131_sum_i_0_8 ));
    InMux I__3606 (
            .O(N__21610),
            .I(N__21607));
    LocalMux I__3605 (
            .O(N__21607),
            .I(\b2v_inst11.mult1_un145_sum_axb_8 ));
    InMux I__3604 (
            .O(N__21604),
            .I(\b2v_inst11.mult1_un138_sum_cry_6 ));
    InMux I__3603 (
            .O(N__21601),
            .I(N__21592));
    InMux I__3602 (
            .O(N__21600),
            .I(N__21592));
    InMux I__3601 (
            .O(N__21599),
            .I(N__21586));
    InMux I__3600 (
            .O(N__21598),
            .I(N__21586));
    InMux I__3599 (
            .O(N__21597),
            .I(N__21583));
    LocalMux I__3598 (
            .O(N__21592),
            .I(N__21580));
    InMux I__3597 (
            .O(N__21591),
            .I(N__21577));
    LocalMux I__3596 (
            .O(N__21586),
            .I(N__21574));
    LocalMux I__3595 (
            .O(N__21583),
            .I(N__21571));
    Span4Mux_h I__3594 (
            .O(N__21580),
            .I(N__21568));
    LocalMux I__3593 (
            .O(N__21577),
            .I(N__21563));
    Span4Mux_v I__3592 (
            .O(N__21574),
            .I(N__21563));
    Span4Mux_s3_h I__3591 (
            .O(N__21571),
            .I(N__21560));
    Odrv4 I__3590 (
            .O(N__21568),
            .I(\b2v_inst11.func_state_RNI_1Z0Z_1 ));
    Odrv4 I__3589 (
            .O(N__21563),
            .I(\b2v_inst11.func_state_RNI_1Z0Z_1 ));
    Odrv4 I__3588 (
            .O(N__21560),
            .I(\b2v_inst11.func_state_RNI_1Z0Z_1 ));
    InMux I__3587 (
            .O(N__21553),
            .I(N__21550));
    LocalMux I__3586 (
            .O(N__21550),
            .I(\b2v_inst11.func_state_1_m2s2_i_1 ));
    InMux I__3585 (
            .O(N__21547),
            .I(N__21544));
    LocalMux I__3584 (
            .O(N__21544),
            .I(\b2v_inst11.N_73 ));
    InMux I__3583 (
            .O(N__21541),
            .I(N__21538));
    LocalMux I__3582 (
            .O(N__21538),
            .I(\b2v_inst11.func_state_1_m0_0 ));
    CascadeMux I__3581 (
            .O(N__21535),
            .I(\b2v_inst11.N_73_cascade_ ));
    InMux I__3580 (
            .O(N__21532),
            .I(N__21529));
    LocalMux I__3579 (
            .O(N__21529),
            .I(\b2v_inst11.count_off_RNIQCBN4Z0Z_9 ));
    InMux I__3578 (
            .O(N__21526),
            .I(N__21523));
    LocalMux I__3577 (
            .O(N__21523),
            .I(\b2v_inst11.func_state_1_m0_1 ));
    InMux I__3576 (
            .O(N__21520),
            .I(\b2v_inst11.mult1_un145_sum_cry_2 ));
    InMux I__3575 (
            .O(N__21517),
            .I(\b2v_inst11.mult1_un145_sum_cry_3 ));
    InMux I__3574 (
            .O(N__21514),
            .I(\b2v_inst11.mult1_un145_sum_cry_4 ));
    InMux I__3573 (
            .O(N__21511),
            .I(\b2v_inst11.mult1_un145_sum_cry_5 ));
    InMux I__3572 (
            .O(N__21508),
            .I(\b2v_inst11.mult1_un145_sum_cry_6 ));
    InMux I__3571 (
            .O(N__21505),
            .I(N__21502));
    LocalMux I__3570 (
            .O(N__21502),
            .I(N__21499));
    Span4Mux_h I__3569 (
            .O(N__21499),
            .I(N__21496));
    Odrv4 I__3568 (
            .O(N__21496),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_307_N ));
    InMux I__3567 (
            .O(N__21493),
            .I(N__21489));
    InMux I__3566 (
            .O(N__21492),
            .I(N__21486));
    LocalMux I__3565 (
            .O(N__21489),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_5 ));
    LocalMux I__3564 (
            .O(N__21486),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_5 ));
    CascadeMux I__3563 (
            .O(N__21481),
            .I(\b2v_inst11.N_4_cascade_ ));
    CascadeMux I__3562 (
            .O(N__21478),
            .I(\b2v_inst11.func_state_RNI_0Z0Z_0_cascade_ ));
    InMux I__3561 (
            .O(N__21475),
            .I(N__21472));
    LocalMux I__3560 (
            .O(N__21472),
            .I(\b2v_inst11.func_state_RNINJ641_0Z0Z_0 ));
    CascadeMux I__3559 (
            .O(N__21469),
            .I(\b2v_inst11.func_state_RNINJ641_0Z0Z_0_cascade_ ));
    CascadeMux I__3558 (
            .O(N__21466),
            .I(\b2v_inst11.count_off_RNIQCBN4Z0Z_9_cascade_ ));
    InMux I__3557 (
            .O(N__21463),
            .I(N__21460));
    LocalMux I__3556 (
            .O(N__21460),
            .I(\b2v_inst11.N_333 ));
    CascadeMux I__3555 (
            .O(N__21457),
            .I(N__21454));
    InMux I__3554 (
            .O(N__21454),
            .I(N__21448));
    InMux I__3553 (
            .O(N__21453),
            .I(N__21448));
    LocalMux I__3552 (
            .O(N__21448),
            .I(\b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNPZ0Z5 ));
    InMux I__3551 (
            .O(N__21445),
            .I(\b2v_inst11.un1_dutycycle_94_cry_10 ));
    InMux I__3550 (
            .O(N__21442),
            .I(N__21437));
    CascadeMux I__3549 (
            .O(N__21441),
            .I(N__21430));
    InMux I__3548 (
            .O(N__21440),
            .I(N__21427));
    LocalMux I__3547 (
            .O(N__21437),
            .I(N__21424));
    InMux I__3546 (
            .O(N__21436),
            .I(N__21421));
    InMux I__3545 (
            .O(N__21435),
            .I(N__21418));
    InMux I__3544 (
            .O(N__21434),
            .I(N__21410));
    InMux I__3543 (
            .O(N__21433),
            .I(N__21410));
    InMux I__3542 (
            .O(N__21430),
            .I(N__21406));
    LocalMux I__3541 (
            .O(N__21427),
            .I(N__21399));
    Span4Mux_v I__3540 (
            .O(N__21424),
            .I(N__21399));
    LocalMux I__3539 (
            .O(N__21421),
            .I(N__21399));
    LocalMux I__3538 (
            .O(N__21418),
            .I(N__21396));
    InMux I__3537 (
            .O(N__21417),
            .I(N__21389));
    InMux I__3536 (
            .O(N__21416),
            .I(N__21389));
    InMux I__3535 (
            .O(N__21415),
            .I(N__21386));
    LocalMux I__3534 (
            .O(N__21410),
            .I(N__21383));
    InMux I__3533 (
            .O(N__21409),
            .I(N__21380));
    LocalMux I__3532 (
            .O(N__21406),
            .I(N__21373));
    Span4Mux_v I__3531 (
            .O(N__21399),
            .I(N__21373));
    Span4Mux_s3_v I__3530 (
            .O(N__21396),
            .I(N__21373));
    InMux I__3529 (
            .O(N__21395),
            .I(N__21368));
    InMux I__3528 (
            .O(N__21394),
            .I(N__21368));
    LocalMux I__3527 (
            .O(N__21389),
            .I(\b2v_inst11.dutycycleZ0Z_10 ));
    LocalMux I__3526 (
            .O(N__21386),
            .I(\b2v_inst11.dutycycleZ0Z_10 ));
    Odrv4 I__3525 (
            .O(N__21383),
            .I(\b2v_inst11.dutycycleZ0Z_10 ));
    LocalMux I__3524 (
            .O(N__21380),
            .I(\b2v_inst11.dutycycleZ0Z_10 ));
    Odrv4 I__3523 (
            .O(N__21373),
            .I(\b2v_inst11.dutycycleZ0Z_10 ));
    LocalMux I__3522 (
            .O(N__21368),
            .I(\b2v_inst11.dutycycleZ0Z_10 ));
    InMux I__3521 (
            .O(N__21355),
            .I(N__21349));
    InMux I__3520 (
            .O(N__21354),
            .I(N__21349));
    LocalMux I__3519 (
            .O(N__21349),
            .I(N__21346));
    Span4Mux_h I__3518 (
            .O(N__21346),
            .I(N__21343));
    Odrv4 I__3517 (
            .O(N__21343),
            .I(\b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQZ0Z5 ));
    InMux I__3516 (
            .O(N__21340),
            .I(\b2v_inst11.un1_dutycycle_94_cry_11 ));
    CascadeMux I__3515 (
            .O(N__21337),
            .I(N__21332));
    InMux I__3514 (
            .O(N__21336),
            .I(N__21329));
    InMux I__3513 (
            .O(N__21335),
            .I(N__21326));
    InMux I__3512 (
            .O(N__21332),
            .I(N__21321));
    LocalMux I__3511 (
            .O(N__21329),
            .I(N__21318));
    LocalMux I__3510 (
            .O(N__21326),
            .I(N__21315));
    InMux I__3509 (
            .O(N__21325),
            .I(N__21310));
    InMux I__3508 (
            .O(N__21324),
            .I(N__21307));
    LocalMux I__3507 (
            .O(N__21321),
            .I(N__21303));
    Span4Mux_h I__3506 (
            .O(N__21318),
            .I(N__21300));
    Span4Mux_v I__3505 (
            .O(N__21315),
            .I(N__21297));
    InMux I__3504 (
            .O(N__21314),
            .I(N__21294));
    InMux I__3503 (
            .O(N__21313),
            .I(N__21291));
    LocalMux I__3502 (
            .O(N__21310),
            .I(N__21286));
    LocalMux I__3501 (
            .O(N__21307),
            .I(N__21286));
    InMux I__3500 (
            .O(N__21306),
            .I(N__21283));
    Span12Mux_s8_h I__3499 (
            .O(N__21303),
            .I(N__21280));
    Odrv4 I__3498 (
            .O(N__21300),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    Odrv4 I__3497 (
            .O(N__21297),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    LocalMux I__3496 (
            .O(N__21294),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    LocalMux I__3495 (
            .O(N__21291),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    Odrv4 I__3494 (
            .O(N__21286),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    LocalMux I__3493 (
            .O(N__21283),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    Odrv12 I__3492 (
            .O(N__21280),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    InMux I__3491 (
            .O(N__21265),
            .I(N__21259));
    InMux I__3490 (
            .O(N__21264),
            .I(N__21259));
    LocalMux I__3489 (
            .O(N__21259),
            .I(N__21256));
    Span4Mux_h I__3488 (
            .O(N__21256),
            .I(N__21253));
    Odrv4 I__3487 (
            .O(N__21253),
            .I(\b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5 ));
    InMux I__3486 (
            .O(N__21250),
            .I(\b2v_inst11.un1_dutycycle_94_cry_12 ));
    InMux I__3485 (
            .O(N__21247),
            .I(N__21241));
    InMux I__3484 (
            .O(N__21246),
            .I(N__21235));
    InMux I__3483 (
            .O(N__21245),
            .I(N__21235));
    InMux I__3482 (
            .O(N__21244),
            .I(N__21232));
    LocalMux I__3481 (
            .O(N__21241),
            .I(N__21228));
    CascadeMux I__3480 (
            .O(N__21240),
            .I(N__21225));
    LocalMux I__3479 (
            .O(N__21235),
            .I(N__21220));
    LocalMux I__3478 (
            .O(N__21232),
            .I(N__21217));
    InMux I__3477 (
            .O(N__21231),
            .I(N__21214));
    Span4Mux_v I__3476 (
            .O(N__21228),
            .I(N__21211));
    InMux I__3475 (
            .O(N__21225),
            .I(N__21206));
    InMux I__3474 (
            .O(N__21224),
            .I(N__21206));
    InMux I__3473 (
            .O(N__21223),
            .I(N__21203));
    Span4Mux_h I__3472 (
            .O(N__21220),
            .I(N__21200));
    Odrv12 I__3471 (
            .O(N__21217),
            .I(\b2v_inst11.dutycycleZ0Z_13 ));
    LocalMux I__3470 (
            .O(N__21214),
            .I(\b2v_inst11.dutycycleZ0Z_13 ));
    Odrv4 I__3469 (
            .O(N__21211),
            .I(\b2v_inst11.dutycycleZ0Z_13 ));
    LocalMux I__3468 (
            .O(N__21206),
            .I(\b2v_inst11.dutycycleZ0Z_13 ));
    LocalMux I__3467 (
            .O(N__21203),
            .I(\b2v_inst11.dutycycleZ0Z_13 ));
    Odrv4 I__3466 (
            .O(N__21200),
            .I(\b2v_inst11.dutycycleZ0Z_13 ));
    CascadeMux I__3465 (
            .O(N__21187),
            .I(N__21183));
    CascadeMux I__3464 (
            .O(N__21186),
            .I(N__21180));
    InMux I__3463 (
            .O(N__21183),
            .I(N__21177));
    InMux I__3462 (
            .O(N__21180),
            .I(N__21174));
    LocalMux I__3461 (
            .O(N__21177),
            .I(N__21169));
    LocalMux I__3460 (
            .O(N__21174),
            .I(N__21169));
    Odrv12 I__3459 (
            .O(N__21169),
            .I(\b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5 ));
    InMux I__3458 (
            .O(N__21166),
            .I(\b2v_inst11.un1_dutycycle_94_cry_13 ));
    InMux I__3457 (
            .O(N__21163),
            .I(N__21160));
    LocalMux I__3456 (
            .O(N__21160),
            .I(N__21157));
    Span4Mux_s3_v I__3455 (
            .O(N__21157),
            .I(N__21150));
    InMux I__3454 (
            .O(N__21156),
            .I(N__21144));
    InMux I__3453 (
            .O(N__21155),
            .I(N__21144));
    CascadeMux I__3452 (
            .O(N__21154),
            .I(N__21141));
    InMux I__3451 (
            .O(N__21153),
            .I(N__21137));
    Span4Mux_v I__3450 (
            .O(N__21150),
            .I(N__21134));
    InMux I__3449 (
            .O(N__21149),
            .I(N__21131));
    LocalMux I__3448 (
            .O(N__21144),
            .I(N__21128));
    InMux I__3447 (
            .O(N__21141),
            .I(N__21123));
    InMux I__3446 (
            .O(N__21140),
            .I(N__21123));
    LocalMux I__3445 (
            .O(N__21137),
            .I(N__21120));
    Odrv4 I__3444 (
            .O(N__21134),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    LocalMux I__3443 (
            .O(N__21131),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    Odrv4 I__3442 (
            .O(N__21128),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    LocalMux I__3441 (
            .O(N__21123),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    Odrv4 I__3440 (
            .O(N__21120),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    InMux I__3439 (
            .O(N__21109),
            .I(\b2v_inst11.un1_dutycycle_94_cry_14 ));
    CascadeMux I__3438 (
            .O(N__21106),
            .I(N__21102));
    InMux I__3437 (
            .O(N__21105),
            .I(N__21099));
    InMux I__3436 (
            .O(N__21102),
            .I(N__21096));
    LocalMux I__3435 (
            .O(N__21099),
            .I(N__21091));
    LocalMux I__3434 (
            .O(N__21096),
            .I(N__21091));
    Span12Mux_s5_h I__3433 (
            .O(N__21091),
            .I(N__21088));
    Odrv12 I__3432 (
            .O(N__21088),
            .I(\b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5 ));
    CascadeMux I__3431 (
            .O(N__21085),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_5_cascade_ ));
    InMux I__3430 (
            .O(N__21082),
            .I(N__21079));
    LocalMux I__3429 (
            .O(N__21079),
            .I(\b2v_inst11.N_156 ));
    CascadeMux I__3428 (
            .O(N__21076),
            .I(\b2v_inst11.N_156_cascade_ ));
    InMux I__3427 (
            .O(N__21073),
            .I(N__21070));
    LocalMux I__3426 (
            .O(N__21070),
            .I(\b2v_inst11.N_331 ));
    InMux I__3425 (
            .O(N__21067),
            .I(\b2v_inst11.un1_dutycycle_94_cry_2 ));
    InMux I__3424 (
            .O(N__21064),
            .I(N__21058));
    InMux I__3423 (
            .O(N__21063),
            .I(N__21058));
    LocalMux I__3422 (
            .O(N__21058),
            .I(N__21055));
    Odrv4 I__3421 (
            .O(N__21055),
            .I(\b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09 ));
    InMux I__3420 (
            .O(N__21052),
            .I(\b2v_inst11.un1_dutycycle_94_cry_3 ));
    InMux I__3419 (
            .O(N__21049),
            .I(\b2v_inst11.un1_dutycycle_94_cry_4 ));
    InMux I__3418 (
            .O(N__21046),
            .I(\b2v_inst11.un1_dutycycle_94_cry_5_cZ0 ));
    InMux I__3417 (
            .O(N__21043),
            .I(N__21040));
    LocalMux I__3416 (
            .O(N__21040),
            .I(\b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39 ));
    InMux I__3415 (
            .O(N__21037),
            .I(\b2v_inst11.un1_dutycycle_94_cry_6_cZ0 ));
    CascadeMux I__3414 (
            .O(N__21034),
            .I(N__21031));
    InMux I__3413 (
            .O(N__21031),
            .I(N__21028));
    LocalMux I__3412 (
            .O(N__21028),
            .I(N__21025));
    Span4Mux_h I__3411 (
            .O(N__21025),
            .I(N__21022));
    Odrv4 I__3410 (
            .O(N__21022),
            .I(\b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHPZ0Z49 ));
    InMux I__3409 (
            .O(N__21019),
            .I(bfn_6_14_0_));
    CascadeMux I__3408 (
            .O(N__21016),
            .I(N__21008));
    InMux I__3407 (
            .O(N__21015),
            .I(N__21005));
    InMux I__3406 (
            .O(N__21014),
            .I(N__21002));
    InMux I__3405 (
            .O(N__21013),
            .I(N__20999));
    InMux I__3404 (
            .O(N__21012),
            .I(N__20989));
    InMux I__3403 (
            .O(N__21011),
            .I(N__20989));
    InMux I__3402 (
            .O(N__21008),
            .I(N__20986));
    LocalMux I__3401 (
            .O(N__21005),
            .I(N__20983));
    LocalMux I__3400 (
            .O(N__21002),
            .I(N__20980));
    LocalMux I__3399 (
            .O(N__20999),
            .I(N__20977));
    InMux I__3398 (
            .O(N__20998),
            .I(N__20971));
    InMux I__3397 (
            .O(N__20997),
            .I(N__20971));
    InMux I__3396 (
            .O(N__20996),
            .I(N__20968));
    InMux I__3395 (
            .O(N__20995),
            .I(N__20963));
    InMux I__3394 (
            .O(N__20994),
            .I(N__20963));
    LocalMux I__3393 (
            .O(N__20989),
            .I(N__20960));
    LocalMux I__3392 (
            .O(N__20986),
            .I(N__20949));
    Span4Mux_v I__3391 (
            .O(N__20983),
            .I(N__20949));
    Span4Mux_h I__3390 (
            .O(N__20980),
            .I(N__20949));
    Span4Mux_h I__3389 (
            .O(N__20977),
            .I(N__20946));
    InMux I__3388 (
            .O(N__20976),
            .I(N__20943));
    LocalMux I__3387 (
            .O(N__20971),
            .I(N__20934));
    LocalMux I__3386 (
            .O(N__20968),
            .I(N__20934));
    LocalMux I__3385 (
            .O(N__20963),
            .I(N__20934));
    Span4Mux_h I__3384 (
            .O(N__20960),
            .I(N__20934));
    InMux I__3383 (
            .O(N__20959),
            .I(N__20925));
    InMux I__3382 (
            .O(N__20958),
            .I(N__20925));
    InMux I__3381 (
            .O(N__20957),
            .I(N__20925));
    InMux I__3380 (
            .O(N__20956),
            .I(N__20925));
    Odrv4 I__3379 (
            .O(N__20949),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    Odrv4 I__3378 (
            .O(N__20946),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    LocalMux I__3377 (
            .O(N__20943),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    Odrv4 I__3376 (
            .O(N__20934),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    LocalMux I__3375 (
            .O(N__20925),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    CascadeMux I__3374 (
            .O(N__20914),
            .I(N__20911));
    InMux I__3373 (
            .O(N__20911),
            .I(N__20905));
    InMux I__3372 (
            .O(N__20910),
            .I(N__20905));
    LocalMux I__3371 (
            .O(N__20905),
            .I(N__20902));
    Odrv4 I__3370 (
            .O(N__20902),
            .I(\b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59 ));
    InMux I__3369 (
            .O(N__20899),
            .I(\b2v_inst11.un1_dutycycle_94_cry_8_cZ0 ));
    InMux I__3368 (
            .O(N__20896),
            .I(\b2v_inst11.un1_dutycycle_94_cry_9_cZ0 ));
    CascadeMux I__3367 (
            .O(N__20893),
            .I(N__20887));
    InMux I__3366 (
            .O(N__20892),
            .I(N__20884));
    InMux I__3365 (
            .O(N__20891),
            .I(N__20881));
    InMux I__3364 (
            .O(N__20890),
            .I(N__20877));
    InMux I__3363 (
            .O(N__20887),
            .I(N__20871));
    LocalMux I__3362 (
            .O(N__20884),
            .I(N__20866));
    LocalMux I__3361 (
            .O(N__20881),
            .I(N__20866));
    InMux I__3360 (
            .O(N__20880),
            .I(N__20863));
    LocalMux I__3359 (
            .O(N__20877),
            .I(N__20860));
    InMux I__3358 (
            .O(N__20876),
            .I(N__20853));
    InMux I__3357 (
            .O(N__20875),
            .I(N__20853));
    InMux I__3356 (
            .O(N__20874),
            .I(N__20853));
    LocalMux I__3355 (
            .O(N__20871),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    Odrv12 I__3354 (
            .O(N__20866),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    LocalMux I__3353 (
            .O(N__20863),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    Odrv4 I__3352 (
            .O(N__20860),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    LocalMux I__3351 (
            .O(N__20853),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    CascadeMux I__3350 (
            .O(N__20842),
            .I(\b2v_inst11.dutycycle_RNI74A23Z0Z_7_cascade_ ));
    InMux I__3349 (
            .O(N__20839),
            .I(N__20836));
    LocalMux I__3348 (
            .O(N__20836),
            .I(\b2v_inst11.dutycycle_e_1_7 ));
    InMux I__3347 (
            .O(N__20833),
            .I(N__20830));
    LocalMux I__3346 (
            .O(N__20830),
            .I(\b2v_inst11.dutycycle_RNI74A23Z0Z_7 ));
    CascadeMux I__3345 (
            .O(N__20827),
            .I(\b2v_inst11.dutycycle_e_1_7_cascade_ ));
    InMux I__3344 (
            .O(N__20824),
            .I(N__20821));
    LocalMux I__3343 (
            .O(N__20821),
            .I(N__20818));
    Span4Mux_h I__3342 (
            .O(N__20818),
            .I(N__20815));
    Odrv4 I__3341 (
            .O(N__20815),
            .I(\b2v_inst11.dutycycle_RNI01TT1Z0Z_7 ));
    CascadeMux I__3340 (
            .O(N__20812),
            .I(\b2v_inst11.dutycycle_RNI25OT3Z0Z_7_cascade_ ));
    CascadeMux I__3339 (
            .O(N__20809),
            .I(N__20806));
    InMux I__3338 (
            .O(N__20806),
            .I(N__20803));
    LocalMux I__3337 (
            .O(N__20803),
            .I(\b2v_inst11.func_state_RNIGALV4Z0Z_0 ));
    InMux I__3336 (
            .O(N__20800),
            .I(N__20788));
    InMux I__3335 (
            .O(N__20799),
            .I(N__20788));
    InMux I__3334 (
            .O(N__20798),
            .I(N__20788));
    InMux I__3333 (
            .O(N__20797),
            .I(N__20788));
    LocalMux I__3332 (
            .O(N__20788),
            .I(\b2v_inst11.dutycycleZ1Z_7 ));
    InMux I__3331 (
            .O(N__20785),
            .I(N__20782));
    LocalMux I__3330 (
            .O(N__20782),
            .I(\b2v_inst11.dutycycle_RNIGSFQZ0Z_7 ));
    InMux I__3329 (
            .O(N__20779),
            .I(\b2v_inst11.un1_dutycycle_94_cry_0_cZ0 ));
    InMux I__3328 (
            .O(N__20776),
            .I(N__20773));
    LocalMux I__3327 (
            .O(N__20773),
            .I(N__20770));
    Span4Mux_h I__3326 (
            .O(N__20770),
            .I(N__20767));
    Odrv4 I__3325 (
            .O(N__20767),
            .I(\b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDUZ0Z8 ));
    InMux I__3324 (
            .O(N__20764),
            .I(\b2v_inst11.un1_dutycycle_94_cry_1 ));
    CascadeMux I__3323 (
            .O(N__20761),
            .I(\b2v_inst11.dutycycleZ0Z_8_cascade_ ));
    CascadeMux I__3322 (
            .O(N__20758),
            .I(\b2v_inst11.dutycycle_RNIAI7C4Z0Z_4_cascade_ ));
    CascadeMux I__3321 (
            .O(N__20755),
            .I(N__20752));
    InMux I__3320 (
            .O(N__20752),
            .I(N__20749));
    LocalMux I__3319 (
            .O(N__20749),
            .I(\b2v_inst11.dutycycle_eena_2_0_1 ));
    CascadeMux I__3318 (
            .O(N__20746),
            .I(\b2v_inst11.func_state_RNI3JFN6Z0Z_0_cascade_ ));
    InMux I__3317 (
            .O(N__20743),
            .I(N__20737));
    InMux I__3316 (
            .O(N__20742),
            .I(N__20737));
    LocalMux I__3315 (
            .O(N__20737),
            .I(\b2v_inst11.dutycycle_RNI3JFN6Z0Z_4 ));
    CascadeMux I__3314 (
            .O(N__20734),
            .I(N__20730));
    CascadeMux I__3313 (
            .O(N__20733),
            .I(N__20727));
    InMux I__3312 (
            .O(N__20730),
            .I(N__20722));
    InMux I__3311 (
            .O(N__20727),
            .I(N__20722));
    LocalMux I__3310 (
            .O(N__20722),
            .I(\b2v_inst11.dutycycleZ1Z_4 ));
    InMux I__3309 (
            .O(N__20719),
            .I(N__20713));
    InMux I__3308 (
            .O(N__20718),
            .I(N__20713));
    LocalMux I__3307 (
            .O(N__20713),
            .I(\b2v_inst11.dutycycleZ1Z_9 ));
    InMux I__3306 (
            .O(N__20710),
            .I(N__20707));
    LocalMux I__3305 (
            .O(N__20707),
            .I(\b2v_inst11.func_state_RNI3JFN6Z0Z_0 ));
    CascadeMux I__3304 (
            .O(N__20704),
            .I(\b2v_inst11.dutycycle_RNI0KJ31Z0Z_7_cascade_ ));
    InMux I__3303 (
            .O(N__20701),
            .I(N__20695));
    InMux I__3302 (
            .O(N__20700),
            .I(N__20695));
    LocalMux I__3301 (
            .O(N__20695),
            .I(\b2v_inst11.dutycycleZ0Z_14 ));
    InMux I__3300 (
            .O(N__20692),
            .I(N__20688));
    InMux I__3299 (
            .O(N__20691),
            .I(N__20685));
    LocalMux I__3298 (
            .O(N__20688),
            .I(N__20680));
    LocalMux I__3297 (
            .O(N__20685),
            .I(N__20680));
    Odrv4 I__3296 (
            .O(N__20680),
            .I(\b2v_inst11.dutycycle_en_11 ));
    CascadeMux I__3295 (
            .O(N__20677),
            .I(\b2v_inst11.dutycycleZ0Z_13_cascade_ ));
    InMux I__3294 (
            .O(N__20674),
            .I(N__20671));
    LocalMux I__3293 (
            .O(N__20671),
            .I(\b2v_inst11.un2_count_clk_17_0_a2_1_4 ));
    InMux I__3292 (
            .O(N__20668),
            .I(N__20665));
    LocalMux I__3291 (
            .O(N__20665),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_4 ));
    CascadeMux I__3290 (
            .O(N__20662),
            .I(\b2v_inst11.un1_dutycycle_53_50_a4_0_cascade_ ));
    InMux I__3289 (
            .O(N__20659),
            .I(N__20655));
    InMux I__3288 (
            .O(N__20658),
            .I(N__20652));
    LocalMux I__3287 (
            .O(N__20655),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_10 ));
    LocalMux I__3286 (
            .O(N__20652),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_10 ));
    InMux I__3285 (
            .O(N__20647),
            .I(N__20644));
    LocalMux I__3284 (
            .O(N__20644),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_7 ));
    InMux I__3283 (
            .O(N__20641),
            .I(N__20638));
    LocalMux I__3282 (
            .O(N__20638),
            .I(N__20635));
    Sp12to4 I__3281 (
            .O(N__20635),
            .I(N__20632));
    Odrv12 I__3280 (
            .O(N__20632),
            .I(VCCST_OK_c));
    InMux I__3279 (
            .O(N__20629),
            .I(N__20619));
    InMux I__3278 (
            .O(N__20628),
            .I(N__20619));
    InMux I__3277 (
            .O(N__20627),
            .I(N__20619));
    InMux I__3276 (
            .O(N__20626),
            .I(N__20616));
    LocalMux I__3275 (
            .O(N__20619),
            .I(N__20613));
    LocalMux I__3274 (
            .O(N__20616),
            .I(N__20610));
    Odrv12 I__3273 (
            .O(N__20613),
            .I(VDDQ_OK_c));
    Odrv12 I__3272 (
            .O(N__20610),
            .I(VDDQ_OK_c));
    IoInMux I__3271 (
            .O(N__20605),
            .I(N__20602));
    LocalMux I__3270 (
            .O(N__20602),
            .I(N__20599));
    Odrv12 I__3269 (
            .O(N__20599),
            .I(VCCIO_EN_c));
    InMux I__3268 (
            .O(N__20596),
            .I(N__20593));
    LocalMux I__3267 (
            .O(N__20593),
            .I(N__20589));
    InMux I__3266 (
            .O(N__20592),
            .I(N__20586));
    Odrv4 I__3265 (
            .O(N__20589),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_3 ));
    LocalMux I__3264 (
            .O(N__20586),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_3 ));
    CascadeMux I__3263 (
            .O(N__20581),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_3_cascade_ ));
    InMux I__3262 (
            .O(N__20578),
            .I(N__20575));
    LocalMux I__3261 (
            .O(N__20575),
            .I(\b2v_inst11.un1_dutycycle_53_axb_7_1 ));
    CascadeMux I__3260 (
            .O(N__20572),
            .I(N__20569));
    InMux I__3259 (
            .O(N__20569),
            .I(N__20566));
    LocalMux I__3258 (
            .O(N__20566),
            .I(N__20563));
    Odrv4 I__3257 (
            .O(N__20563),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_9 ));
    InMux I__3256 (
            .O(N__20560),
            .I(N__20557));
    LocalMux I__3255 (
            .O(N__20557),
            .I(\b2v_inst16.curr_state_1_0 ));
    InMux I__3254 (
            .O(N__20554),
            .I(N__20551));
    LocalMux I__3253 (
            .O(N__20551),
            .I(\b2v_inst16.curr_stateZ0Z_0 ));
    CascadeMux I__3252 (
            .O(N__20548),
            .I(N__20545));
    InMux I__3251 (
            .O(N__20545),
            .I(N__20537));
    InMux I__3250 (
            .O(N__20544),
            .I(N__20526));
    InMux I__3249 (
            .O(N__20543),
            .I(N__20526));
    InMux I__3248 (
            .O(N__20542),
            .I(N__20526));
    InMux I__3247 (
            .O(N__20541),
            .I(N__20526));
    InMux I__3246 (
            .O(N__20540),
            .I(N__20526));
    LocalMux I__3245 (
            .O(N__20537),
            .I(\b2v_inst16.curr_stateZ0Z_1 ));
    LocalMux I__3244 (
            .O(N__20526),
            .I(\b2v_inst16.curr_stateZ0Z_1 ));
    CascadeMux I__3243 (
            .O(N__20521),
            .I(N__20518));
    InMux I__3242 (
            .O(N__20518),
            .I(N__20515));
    LocalMux I__3241 (
            .O(N__20515),
            .I(N__20512));
    Odrv4 I__3240 (
            .O(N__20512),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_0 ));
    InMux I__3239 (
            .O(N__20509),
            .I(N__20506));
    LocalMux I__3238 (
            .O(N__20506),
            .I(N__20503));
    Span4Mux_h I__3237 (
            .O(N__20503),
            .I(N__20500));
    Span4Mux_h I__3236 (
            .O(N__20500),
            .I(N__20497));
    Odrv4 I__3235 (
            .O(N__20497),
            .I(\b2v_inst200.count_RNIC03N_3Z0Z_0 ));
    IoInMux I__3234 (
            .O(N__20494),
            .I(N__20490));
    IoInMux I__3233 (
            .O(N__20493),
            .I(N__20487));
    LocalMux I__3232 (
            .O(N__20490),
            .I(N__20484));
    LocalMux I__3231 (
            .O(N__20487),
            .I(N__20481));
    Span4Mux_s1_h I__3230 (
            .O(N__20484),
            .I(N__20478));
    IoSpan4Mux I__3229 (
            .O(N__20481),
            .I(N__20475));
    Span4Mux_v I__3228 (
            .O(N__20478),
            .I(N__20470));
    Span4Mux_s1_h I__3227 (
            .O(N__20475),
            .I(N__20470));
    Span4Mux_h I__3226 (
            .O(N__20470),
            .I(N__20467));
    Odrv4 I__3225 (
            .O(N__20467),
            .I(V105A_EN_c));
    CascadeMux I__3224 (
            .O(N__20464),
            .I(N__20461));
    InMux I__3223 (
            .O(N__20461),
            .I(N__20458));
    LocalMux I__3222 (
            .O(N__20458),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_5 ));
    InMux I__3221 (
            .O(N__20455),
            .I(N__20452));
    LocalMux I__3220 (
            .O(N__20452),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_10 ));
    InMux I__3219 (
            .O(N__20449),
            .I(N__20446));
    LocalMux I__3218 (
            .O(N__20446),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_5 ));
    CascadeMux I__3217 (
            .O(N__20443),
            .I(N__20439));
    InMux I__3216 (
            .O(N__20442),
            .I(N__20436));
    InMux I__3215 (
            .O(N__20439),
            .I(N__20433));
    LocalMux I__3214 (
            .O(N__20436),
            .I(N__20430));
    LocalMux I__3213 (
            .O(N__20433),
            .I(N__20427));
    Odrv4 I__3212 (
            .O(N__20430),
            .I(\b2v_inst11.mult1_un54_sum ));
    Odrv4 I__3211 (
            .O(N__20427),
            .I(\b2v_inst11.mult1_un54_sum ));
    InMux I__3210 (
            .O(N__20422),
            .I(N__20419));
    LocalMux I__3209 (
            .O(N__20419),
            .I(\b2v_inst11.mult1_un54_sum_i ));
    InMux I__3208 (
            .O(N__20416),
            .I(N__20412));
    InMux I__3207 (
            .O(N__20415),
            .I(N__20409));
    LocalMux I__3206 (
            .O(N__20412),
            .I(N__20406));
    LocalMux I__3205 (
            .O(N__20409),
            .I(N__20403));
    Odrv4 I__3204 (
            .O(N__20406),
            .I(\b2v_inst11.mult1_un61_sum ));
    Odrv4 I__3203 (
            .O(N__20403),
            .I(\b2v_inst11.mult1_un61_sum ));
    CascadeMux I__3202 (
            .O(N__20398),
            .I(N__20395));
    InMux I__3201 (
            .O(N__20395),
            .I(N__20392));
    LocalMux I__3200 (
            .O(N__20392),
            .I(\b2v_inst11.mult1_un61_sum_i ));
    CascadeMux I__3199 (
            .O(N__20389),
            .I(N__20385));
    InMux I__3198 (
            .O(N__20388),
            .I(N__20380));
    InMux I__3197 (
            .O(N__20385),
            .I(N__20375));
    InMux I__3196 (
            .O(N__20384),
            .I(N__20375));
    InMux I__3195 (
            .O(N__20383),
            .I(N__20372));
    LocalMux I__3194 (
            .O(N__20380),
            .I(\b2v_inst11.mult1_un68_sum_s_8 ));
    LocalMux I__3193 (
            .O(N__20375),
            .I(\b2v_inst11.mult1_un68_sum_s_8 ));
    LocalMux I__3192 (
            .O(N__20372),
            .I(\b2v_inst11.mult1_un68_sum_s_8 ));
    CascadeMux I__3191 (
            .O(N__20365),
            .I(\b2v_inst16.curr_stateZ0Z_1_cascade_ ));
    CascadeMux I__3190 (
            .O(N__20362),
            .I(\b2v_inst16.curr_state_7_0_cascade_ ));
    InMux I__3189 (
            .O(N__20359),
            .I(N__20353));
    InMux I__3188 (
            .O(N__20358),
            .I(N__20353));
    LocalMux I__3187 (
            .O(N__20353),
            .I(N__20350));
    Span4Mux_h I__3186 (
            .O(N__20350),
            .I(N__20347));
    Span4Mux_v I__3185 (
            .O(N__20347),
            .I(N__20336));
    InMux I__3184 (
            .O(N__20346),
            .I(N__20331));
    InMux I__3183 (
            .O(N__20345),
            .I(N__20331));
    InMux I__3182 (
            .O(N__20344),
            .I(N__20326));
    InMux I__3181 (
            .O(N__20343),
            .I(N__20326));
    InMux I__3180 (
            .O(N__20342),
            .I(N__20319));
    InMux I__3179 (
            .O(N__20341),
            .I(N__20319));
    InMux I__3178 (
            .O(N__20340),
            .I(N__20319));
    InMux I__3177 (
            .O(N__20339),
            .I(N__20316));
    Odrv4 I__3176 (
            .O(N__20336),
            .I(\b2v_inst16.un13_clk_100khz_i ));
    LocalMux I__3175 (
            .O(N__20331),
            .I(\b2v_inst16.un13_clk_100khz_i ));
    LocalMux I__3174 (
            .O(N__20326),
            .I(\b2v_inst16.un13_clk_100khz_i ));
    LocalMux I__3173 (
            .O(N__20319),
            .I(\b2v_inst16.un13_clk_100khz_i ));
    LocalMux I__3172 (
            .O(N__20316),
            .I(\b2v_inst16.un13_clk_100khz_i ));
    CascadeMux I__3171 (
            .O(N__20305),
            .I(N__20302));
    InMux I__3170 (
            .O(N__20302),
            .I(N__20299));
    LocalMux I__3169 (
            .O(N__20299),
            .I(\b2v_inst16.curr_state_0_1 ));
    InMux I__3168 (
            .O(N__20296),
            .I(N__20293));
    LocalMux I__3167 (
            .O(N__20293),
            .I(\b2v_inst16.delayed_vddq_pwrgdZ0 ));
    IoInMux I__3166 (
            .O(N__20290),
            .I(N__20287));
    LocalMux I__3165 (
            .O(N__20287),
            .I(N__20284));
    Span4Mux_s2_h I__3164 (
            .O(N__20284),
            .I(N__20281));
    Span4Mux_h I__3163 (
            .O(N__20281),
            .I(N__20278));
    Odrv4 I__3162 (
            .O(N__20278),
            .I(b2v_inst16_un2_vpp_en_0_i));
    InMux I__3161 (
            .O(N__20275),
            .I(N__20268));
    CascadeMux I__3160 (
            .O(N__20274),
            .I(N__20265));
    InMux I__3159 (
            .O(N__20273),
            .I(N__20256));
    InMux I__3158 (
            .O(N__20272),
            .I(N__20256));
    InMux I__3157 (
            .O(N__20271),
            .I(N__20256));
    LocalMux I__3156 (
            .O(N__20268),
            .I(N__20253));
    InMux I__3155 (
            .O(N__20265),
            .I(N__20248));
    InMux I__3154 (
            .O(N__20264),
            .I(N__20248));
    InMux I__3153 (
            .O(N__20263),
            .I(N__20245));
    LocalMux I__3152 (
            .O(N__20256),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    Odrv4 I__3151 (
            .O(N__20253),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    LocalMux I__3150 (
            .O(N__20248),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    LocalMux I__3149 (
            .O(N__20245),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    InMux I__3148 (
            .O(N__20236),
            .I(N__20233));
    LocalMux I__3147 (
            .O(N__20233),
            .I(N__20229));
    InMux I__3146 (
            .O(N__20232),
            .I(N__20226));
    Span4Mux_s2_v I__3145 (
            .O(N__20229),
            .I(N__20221));
    LocalMux I__3144 (
            .O(N__20226),
            .I(N__20221));
    Odrv4 I__3143 (
            .O(N__20221),
            .I(\b2v_inst11.mult1_un124_sum ));
    InMux I__3142 (
            .O(N__20218),
            .I(N__20215));
    LocalMux I__3141 (
            .O(N__20215),
            .I(\b2v_inst11.mult1_un124_sum_i ));
    InMux I__3140 (
            .O(N__20212),
            .I(N__20209));
    LocalMux I__3139 (
            .O(N__20209),
            .I(N__20205));
    InMux I__3138 (
            .O(N__20208),
            .I(N__20202));
    Span4Mux_h I__3137 (
            .O(N__20205),
            .I(N__20197));
    LocalMux I__3136 (
            .O(N__20202),
            .I(N__20197));
    Span4Mux_v I__3135 (
            .O(N__20197),
            .I(N__20194));
    Odrv4 I__3134 (
            .O(N__20194),
            .I(\b2v_inst11.mult1_un89_sum ));
    CascadeMux I__3133 (
            .O(N__20191),
            .I(N__20188));
    InMux I__3132 (
            .O(N__20188),
            .I(N__20185));
    LocalMux I__3131 (
            .O(N__20185),
            .I(N__20182));
    Span4Mux_s3_v I__3130 (
            .O(N__20182),
            .I(N__20179));
    Odrv4 I__3129 (
            .O(N__20179),
            .I(\b2v_inst11.mult1_un89_sum_i ));
    CascadeMux I__3128 (
            .O(N__20176),
            .I(N__20172));
    InMux I__3127 (
            .O(N__20175),
            .I(N__20164));
    InMux I__3126 (
            .O(N__20172),
            .I(N__20164));
    InMux I__3125 (
            .O(N__20171),
            .I(N__20164));
    LocalMux I__3124 (
            .O(N__20164),
            .I(\b2v_inst11.mult1_un61_sum_i_0_8 ));
    InMux I__3123 (
            .O(N__20161),
            .I(N__20158));
    LocalMux I__3122 (
            .O(N__20158),
            .I(N__20154));
    CascadeMux I__3121 (
            .O(N__20157),
            .I(N__20150));
    Span4Mux_v I__3120 (
            .O(N__20154),
            .I(N__20145));
    InMux I__3119 (
            .O(N__20153),
            .I(N__20142));
    InMux I__3118 (
            .O(N__20150),
            .I(N__20137));
    InMux I__3117 (
            .O(N__20149),
            .I(N__20137));
    InMux I__3116 (
            .O(N__20148),
            .I(N__20134));
    Odrv4 I__3115 (
            .O(N__20145),
            .I(\b2v_inst11.mult1_un110_sum_s_8 ));
    LocalMux I__3114 (
            .O(N__20142),
            .I(\b2v_inst11.mult1_un110_sum_s_8 ));
    LocalMux I__3113 (
            .O(N__20137),
            .I(\b2v_inst11.mult1_un110_sum_s_8 ));
    LocalMux I__3112 (
            .O(N__20134),
            .I(\b2v_inst11.mult1_un110_sum_s_8 ));
    IoInMux I__3111 (
            .O(N__20125),
            .I(N__20122));
    LocalMux I__3110 (
            .O(N__20122),
            .I(N__20119));
    IoSpan4Mux I__3109 (
            .O(N__20119),
            .I(N__20115));
    InMux I__3108 (
            .O(N__20118),
            .I(N__20111));
    Span4Mux_s1_h I__3107 (
            .O(N__20115),
            .I(N__20108));
    InMux I__3106 (
            .O(N__20114),
            .I(N__20105));
    LocalMux I__3105 (
            .O(N__20111),
            .I(N__20102));
    Span4Mux_h I__3104 (
            .O(N__20108),
            .I(N__20097));
    LocalMux I__3103 (
            .O(N__20105),
            .I(N__20097));
    Span4Mux_v I__3102 (
            .O(N__20102),
            .I(N__20093));
    Span4Mux_v I__3101 (
            .O(N__20097),
            .I(N__20090));
    InMux I__3100 (
            .O(N__20096),
            .I(N__20087));
    Odrv4 I__3099 (
            .O(N__20093),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3098 (
            .O(N__20090),
            .I(CONSTANT_ONE_NET));
    LocalMux I__3097 (
            .O(N__20087),
            .I(CONSTANT_ONE_NET));
    InMux I__3096 (
            .O(N__20080),
            .I(N__20077));
    LocalMux I__3095 (
            .O(N__20077),
            .I(N__20073));
    CascadeMux I__3094 (
            .O(N__20076),
            .I(N__20070));
    Span4Mux_v I__3093 (
            .O(N__20073),
            .I(N__20065));
    InMux I__3092 (
            .O(N__20070),
            .I(N__20060));
    InMux I__3091 (
            .O(N__20069),
            .I(N__20060));
    InMux I__3090 (
            .O(N__20068),
            .I(N__20057));
    Odrv4 I__3089 (
            .O(N__20065),
            .I(\b2v_inst11.mult1_un75_sum_s_8 ));
    LocalMux I__3088 (
            .O(N__20060),
            .I(\b2v_inst11.mult1_un75_sum_s_8 ));
    LocalMux I__3087 (
            .O(N__20057),
            .I(\b2v_inst11.mult1_un75_sum_s_8 ));
    CascadeMux I__3086 (
            .O(N__20050),
            .I(N__20046));
    CascadeMux I__3085 (
            .O(N__20049),
            .I(N__20042));
    InMux I__3084 (
            .O(N__20046),
            .I(N__20039));
    InMux I__3083 (
            .O(N__20045),
            .I(N__20034));
    InMux I__3082 (
            .O(N__20042),
            .I(N__20031));
    LocalMux I__3081 (
            .O(N__20039),
            .I(N__20028));
    InMux I__3080 (
            .O(N__20038),
            .I(N__20025));
    InMux I__3079 (
            .O(N__20037),
            .I(N__20022));
    LocalMux I__3078 (
            .O(N__20034),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    LocalMux I__3077 (
            .O(N__20031),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    Odrv4 I__3076 (
            .O(N__20028),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    LocalMux I__3075 (
            .O(N__20025),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    LocalMux I__3074 (
            .O(N__20022),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    InMux I__3073 (
            .O(N__20011),
            .I(N__20008));
    LocalMux I__3072 (
            .O(N__20008),
            .I(N__20004));
    CascadeMux I__3071 (
            .O(N__20007),
            .I(N__20001));
    Span4Mux_v I__3070 (
            .O(N__20004),
            .I(N__19996));
    InMux I__3069 (
            .O(N__20001),
            .I(N__19991));
    InMux I__3068 (
            .O(N__20000),
            .I(N__19991));
    InMux I__3067 (
            .O(N__19999),
            .I(N__19988));
    Odrv4 I__3066 (
            .O(N__19996),
            .I(\b2v_inst11.mult1_un96_sum_s_8 ));
    LocalMux I__3065 (
            .O(N__19991),
            .I(\b2v_inst11.mult1_un96_sum_s_8 ));
    LocalMux I__3064 (
            .O(N__19988),
            .I(\b2v_inst11.mult1_un96_sum_s_8 ));
    InMux I__3063 (
            .O(N__19981),
            .I(\b2v_inst11.mult1_un131_sum_cry_3 ));
    CascadeMux I__3062 (
            .O(N__19978),
            .I(N__19975));
    InMux I__3061 (
            .O(N__19975),
            .I(N__19972));
    LocalMux I__3060 (
            .O(N__19972),
            .I(N__19969));
    Odrv4 I__3059 (
            .O(N__19969),
            .I(\b2v_inst11.mult1_un124_sum_cry_4_s ));
    InMux I__3058 (
            .O(N__19966),
            .I(\b2v_inst11.mult1_un131_sum_cry_4 ));
    InMux I__3057 (
            .O(N__19963),
            .I(N__19960));
    LocalMux I__3056 (
            .O(N__19960),
            .I(\b2v_inst11.mult1_un124_sum_cry_5_s ));
    InMux I__3055 (
            .O(N__19957),
            .I(\b2v_inst11.mult1_un131_sum_cry_5 ));
    InMux I__3054 (
            .O(N__19954),
            .I(N__19951));
    LocalMux I__3053 (
            .O(N__19951),
            .I(\b2v_inst11.mult1_un131_sum_axb_7_l_fx ));
    CascadeMux I__3052 (
            .O(N__19948),
            .I(N__19945));
    InMux I__3051 (
            .O(N__19945),
            .I(N__19941));
    InMux I__3050 (
            .O(N__19944),
            .I(N__19938));
    LocalMux I__3049 (
            .O(N__19941),
            .I(N__19935));
    LocalMux I__3048 (
            .O(N__19938),
            .I(\b2v_inst11.mult1_un124_sum_cry_6_s ));
    Odrv4 I__3047 (
            .O(N__19935),
            .I(\b2v_inst11.mult1_un124_sum_cry_6_s ));
    InMux I__3046 (
            .O(N__19930),
            .I(\b2v_inst11.mult1_un131_sum_cry_6 ));
    InMux I__3045 (
            .O(N__19927),
            .I(N__19924));
    LocalMux I__3044 (
            .O(N__19924),
            .I(\b2v_inst11.mult1_un131_sum_axb_8 ));
    InMux I__3043 (
            .O(N__19921),
            .I(\b2v_inst11.mult1_un131_sum_cry_7 ));
    CascadeMux I__3042 (
            .O(N__19918),
            .I(\b2v_inst11.mult1_un131_sum_s_8_cascade_ ));
    InMux I__3041 (
            .O(N__19915),
            .I(N__19911));
    InMux I__3040 (
            .O(N__19914),
            .I(N__19908));
    LocalMux I__3039 (
            .O(N__19911),
            .I(N__19903));
    LocalMux I__3038 (
            .O(N__19908),
            .I(N__19903));
    Span4Mux_v I__3037 (
            .O(N__19903),
            .I(N__19900));
    Odrv4 I__3036 (
            .O(N__19900),
            .I(\b2v_inst11.mult1_un68_sum ));
    CascadeMux I__3035 (
            .O(N__19897),
            .I(N__19894));
    InMux I__3034 (
            .O(N__19894),
            .I(N__19891));
    LocalMux I__3033 (
            .O(N__19891),
            .I(N__19888));
    Odrv4 I__3032 (
            .O(N__19888),
            .I(\b2v_inst11.mult1_un68_sum_i ));
    InMux I__3031 (
            .O(N__19885),
            .I(N__19881));
    CascadeMux I__3030 (
            .O(N__19884),
            .I(N__19878));
    LocalMux I__3029 (
            .O(N__19881),
            .I(N__19873));
    InMux I__3028 (
            .O(N__19878),
            .I(N__19868));
    InMux I__3027 (
            .O(N__19877),
            .I(N__19868));
    InMux I__3026 (
            .O(N__19876),
            .I(N__19865));
    Odrv12 I__3025 (
            .O(N__19873),
            .I(\b2v_inst11.mult1_un117_sum_s_8 ));
    LocalMux I__3024 (
            .O(N__19868),
            .I(\b2v_inst11.mult1_un117_sum_s_8 ));
    LocalMux I__3023 (
            .O(N__19865),
            .I(\b2v_inst11.mult1_un117_sum_s_8 ));
    InMux I__3022 (
            .O(N__19858),
            .I(N__19855));
    LocalMux I__3021 (
            .O(N__19855),
            .I(N__19851));
    InMux I__3020 (
            .O(N__19854),
            .I(N__19848));
    Span4Mux_s2_v I__3019 (
            .O(N__19851),
            .I(N__19843));
    LocalMux I__3018 (
            .O(N__19848),
            .I(N__19843));
    Odrv4 I__3017 (
            .O(N__19843),
            .I(\b2v_inst11.mult1_un117_sum ));
    CascadeMux I__3016 (
            .O(N__19840),
            .I(N__19837));
    InMux I__3015 (
            .O(N__19837),
            .I(N__19834));
    LocalMux I__3014 (
            .O(N__19834),
            .I(N__19831));
    Odrv4 I__3013 (
            .O(N__19831),
            .I(\b2v_inst11.mult1_un117_sum_i ));
    InMux I__3012 (
            .O(N__19828),
            .I(N__19825));
    LocalMux I__3011 (
            .O(N__19825),
            .I(\b2v_inst11.mult1_un117_sum_cry_3_s ));
    InMux I__3010 (
            .O(N__19822),
            .I(\b2v_inst11.mult1_un124_sum_cry_3 ));
    CascadeMux I__3009 (
            .O(N__19819),
            .I(N__19816));
    InMux I__3008 (
            .O(N__19816),
            .I(N__19813));
    LocalMux I__3007 (
            .O(N__19813),
            .I(\b2v_inst11.mult1_un117_sum_cry_4_s ));
    InMux I__3006 (
            .O(N__19810),
            .I(\b2v_inst11.mult1_un124_sum_cry_4 ));
    InMux I__3005 (
            .O(N__19807),
            .I(N__19804));
    LocalMux I__3004 (
            .O(N__19804),
            .I(\b2v_inst11.mult1_un117_sum_cry_5_s ));
    InMux I__3003 (
            .O(N__19801),
            .I(\b2v_inst11.mult1_un124_sum_cry_5 ));
    CascadeMux I__3002 (
            .O(N__19798),
            .I(N__19794));
    InMux I__3001 (
            .O(N__19797),
            .I(N__19786));
    InMux I__3000 (
            .O(N__19794),
            .I(N__19786));
    InMux I__2999 (
            .O(N__19793),
            .I(N__19786));
    LocalMux I__2998 (
            .O(N__19786),
            .I(\b2v_inst11.mult1_un117_sum_i_0_8 ));
    CascadeMux I__2997 (
            .O(N__19783),
            .I(N__19780));
    InMux I__2996 (
            .O(N__19780),
            .I(N__19777));
    LocalMux I__2995 (
            .O(N__19777),
            .I(\b2v_inst11.mult1_un117_sum_cry_6_s ));
    InMux I__2994 (
            .O(N__19774),
            .I(\b2v_inst11.mult1_un124_sum_cry_6 ));
    InMux I__2993 (
            .O(N__19771),
            .I(N__19768));
    LocalMux I__2992 (
            .O(N__19768),
            .I(\b2v_inst11.mult1_un124_sum_axb_8 ));
    InMux I__2991 (
            .O(N__19765),
            .I(\b2v_inst11.mult1_un124_sum_cry_7 ));
    CascadeMux I__2990 (
            .O(N__19762),
            .I(N__19758));
    InMux I__2989 (
            .O(N__19761),
            .I(N__19750));
    InMux I__2988 (
            .O(N__19758),
            .I(N__19750));
    InMux I__2987 (
            .O(N__19757),
            .I(N__19750));
    LocalMux I__2986 (
            .O(N__19750),
            .I(\b2v_inst11.mult1_un110_sum_i_0_8 ));
    CascadeMux I__2985 (
            .O(N__19747),
            .I(N__19744));
    InMux I__2984 (
            .O(N__19744),
            .I(N__19741));
    LocalMux I__2983 (
            .O(N__19741),
            .I(\b2v_inst11.mult1_un124_sum_i_0_8 ));
    InMux I__2982 (
            .O(N__19738),
            .I(\b2v_inst11.mult1_un131_sum_cry_2 ));
    InMux I__2981 (
            .O(N__19735),
            .I(N__19732));
    LocalMux I__2980 (
            .O(N__19732),
            .I(\b2v_inst11.mult1_un131_sum_axb_4_l_fx ));
    CascadeMux I__2979 (
            .O(N__19729),
            .I(N__19725));
    InMux I__2978 (
            .O(N__19728),
            .I(N__19722));
    InMux I__2977 (
            .O(N__19725),
            .I(N__19719));
    LocalMux I__2976 (
            .O(N__19722),
            .I(\b2v_inst11.mult1_un124_sum_cry_3_s ));
    LocalMux I__2975 (
            .O(N__19719),
            .I(\b2v_inst11.mult1_un124_sum_cry_3_s ));
    CascadeMux I__2974 (
            .O(N__19714),
            .I(N__19711));
    InMux I__2973 (
            .O(N__19711),
            .I(N__19708));
    LocalMux I__2972 (
            .O(N__19708),
            .I(N__19705));
    Odrv4 I__2971 (
            .O(N__19705),
            .I(\b2v_inst11.mult1_un110_sum_i ));
    InMux I__2970 (
            .O(N__19702),
            .I(\b2v_inst11.mult1_un117_sum_cry_2 ));
    InMux I__2969 (
            .O(N__19699),
            .I(N__19696));
    LocalMux I__2968 (
            .O(N__19696),
            .I(\b2v_inst11.mult1_un110_sum_cry_3_s ));
    InMux I__2967 (
            .O(N__19693),
            .I(\b2v_inst11.mult1_un117_sum_cry_3 ));
    CascadeMux I__2966 (
            .O(N__19690),
            .I(N__19687));
    InMux I__2965 (
            .O(N__19687),
            .I(N__19684));
    LocalMux I__2964 (
            .O(N__19684),
            .I(\b2v_inst11.mult1_un110_sum_cry_4_s ));
    InMux I__2963 (
            .O(N__19681),
            .I(\b2v_inst11.mult1_un117_sum_cry_4 ));
    InMux I__2962 (
            .O(N__19678),
            .I(N__19675));
    LocalMux I__2961 (
            .O(N__19675),
            .I(\b2v_inst11.mult1_un110_sum_cry_5_s ));
    InMux I__2960 (
            .O(N__19672),
            .I(\b2v_inst11.mult1_un117_sum_cry_5 ));
    CascadeMux I__2959 (
            .O(N__19669),
            .I(N__19666));
    InMux I__2958 (
            .O(N__19666),
            .I(N__19663));
    LocalMux I__2957 (
            .O(N__19663),
            .I(\b2v_inst11.mult1_un110_sum_cry_6_s ));
    InMux I__2956 (
            .O(N__19660),
            .I(\b2v_inst11.mult1_un117_sum_cry_6 ));
    InMux I__2955 (
            .O(N__19657),
            .I(N__19654));
    LocalMux I__2954 (
            .O(N__19654),
            .I(\b2v_inst11.mult1_un117_sum_axb_8 ));
    InMux I__2953 (
            .O(N__19651),
            .I(\b2v_inst11.mult1_un117_sum_cry_7 ));
    CascadeMux I__2952 (
            .O(N__19648),
            .I(\b2v_inst11.mult1_un117_sum_s_8_cascade_ ));
    InMux I__2951 (
            .O(N__19645),
            .I(\b2v_inst11.mult1_un124_sum_cry_2 ));
    InMux I__2950 (
            .O(N__19642),
            .I(N__19638));
    InMux I__2949 (
            .O(N__19641),
            .I(N__19634));
    LocalMux I__2948 (
            .O(N__19638),
            .I(N__19631));
    CascadeMux I__2947 (
            .O(N__19637),
            .I(N__19628));
    LocalMux I__2946 (
            .O(N__19634),
            .I(N__19625));
    Span4Mux_h I__2945 (
            .O(N__19631),
            .I(N__19622));
    InMux I__2944 (
            .O(N__19628),
            .I(N__19619));
    Span4Mux_h I__2943 (
            .O(N__19625),
            .I(N__19616));
    Odrv4 I__2942 (
            .O(N__19622),
            .I(\b2v_inst11.count_clk_RNI_0Z0Z_1 ));
    LocalMux I__2941 (
            .O(N__19619),
            .I(\b2v_inst11.count_clk_RNI_0Z0Z_1 ));
    Odrv4 I__2940 (
            .O(N__19616),
            .I(\b2v_inst11.count_clk_RNI_0Z0Z_1 ));
    CascadeMux I__2939 (
            .O(N__19609),
            .I(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_1_cascade_ ));
    InMux I__2938 (
            .O(N__19606),
            .I(N__19602));
    InMux I__2937 (
            .O(N__19605),
            .I(N__19599));
    LocalMux I__2936 (
            .O(N__19602),
            .I(N__19596));
    LocalMux I__2935 (
            .O(N__19599),
            .I(N__19593));
    Span4Mux_s2_v I__2934 (
            .O(N__19596),
            .I(N__19590));
    Span4Mux_h I__2933 (
            .O(N__19593),
            .I(N__19585));
    Span4Mux_h I__2932 (
            .O(N__19590),
            .I(N__19585));
    Odrv4 I__2931 (
            .O(N__19585),
            .I(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_0_0 ));
    CascadeMux I__2930 (
            .O(N__19582),
            .I(N__19576));
    CascadeMux I__2929 (
            .O(N__19581),
            .I(N__19558));
    InMux I__2928 (
            .O(N__19580),
            .I(N__19555));
    InMux I__2927 (
            .O(N__19579),
            .I(N__19542));
    InMux I__2926 (
            .O(N__19576),
            .I(N__19542));
    InMux I__2925 (
            .O(N__19575),
            .I(N__19542));
    InMux I__2924 (
            .O(N__19574),
            .I(N__19542));
    InMux I__2923 (
            .O(N__19573),
            .I(N__19542));
    InMux I__2922 (
            .O(N__19572),
            .I(N__19542));
    InMux I__2921 (
            .O(N__19571),
            .I(N__19532));
    InMux I__2920 (
            .O(N__19570),
            .I(N__19532));
    InMux I__2919 (
            .O(N__19569),
            .I(N__19532));
    InMux I__2918 (
            .O(N__19568),
            .I(N__19532));
    InMux I__2917 (
            .O(N__19567),
            .I(N__19523));
    InMux I__2916 (
            .O(N__19566),
            .I(N__19523));
    InMux I__2915 (
            .O(N__19565),
            .I(N__19523));
    InMux I__2914 (
            .O(N__19564),
            .I(N__19523));
    CascadeMux I__2913 (
            .O(N__19563),
            .I(N__19520));
    InMux I__2912 (
            .O(N__19562),
            .I(N__19508));
    InMux I__2911 (
            .O(N__19561),
            .I(N__19508));
    InMux I__2910 (
            .O(N__19558),
            .I(N__19508));
    LocalMux I__2909 (
            .O(N__19555),
            .I(N__19503));
    LocalMux I__2908 (
            .O(N__19542),
            .I(N__19503));
    InMux I__2907 (
            .O(N__19541),
            .I(N__19500));
    LocalMux I__2906 (
            .O(N__19532),
            .I(N__19497));
    LocalMux I__2905 (
            .O(N__19523),
            .I(N__19494));
    InMux I__2904 (
            .O(N__19520),
            .I(N__19481));
    InMux I__2903 (
            .O(N__19519),
            .I(N__19481));
    InMux I__2902 (
            .O(N__19518),
            .I(N__19481));
    InMux I__2901 (
            .O(N__19517),
            .I(N__19481));
    InMux I__2900 (
            .O(N__19516),
            .I(N__19481));
    InMux I__2899 (
            .O(N__19515),
            .I(N__19481));
    LocalMux I__2898 (
            .O(N__19508),
            .I(N__19478));
    Span4Mux_s3_v I__2897 (
            .O(N__19503),
            .I(N__19473));
    LocalMux I__2896 (
            .O(N__19500),
            .I(N__19473));
    Span4Mux_v I__2895 (
            .O(N__19497),
            .I(N__19459));
    Span4Mux_s1_v I__2894 (
            .O(N__19494),
            .I(N__19459));
    LocalMux I__2893 (
            .O(N__19481),
            .I(N__19459));
    Span4Mux_h I__2892 (
            .O(N__19478),
            .I(N__19454));
    Span4Mux_h I__2891 (
            .O(N__19473),
            .I(N__19454));
    InMux I__2890 (
            .O(N__19472),
            .I(N__19439));
    InMux I__2889 (
            .O(N__19471),
            .I(N__19439));
    InMux I__2888 (
            .O(N__19470),
            .I(N__19439));
    InMux I__2887 (
            .O(N__19469),
            .I(N__19439));
    InMux I__2886 (
            .O(N__19468),
            .I(N__19439));
    InMux I__2885 (
            .O(N__19467),
            .I(N__19439));
    InMux I__2884 (
            .O(N__19466),
            .I(N__19439));
    Odrv4 I__2883 (
            .O(N__19459),
            .I(\b2v_inst11.N_122 ));
    Odrv4 I__2882 (
            .O(N__19454),
            .I(\b2v_inst11.N_122 ));
    LocalMux I__2881 (
            .O(N__19439),
            .I(\b2v_inst11.N_122 ));
    InMux I__2880 (
            .O(N__19432),
            .I(N__19423));
    InMux I__2879 (
            .O(N__19431),
            .I(N__19423));
    InMux I__2878 (
            .O(N__19430),
            .I(N__19418));
    InMux I__2877 (
            .O(N__19429),
            .I(N__19418));
    InMux I__2876 (
            .O(N__19428),
            .I(N__19415));
    LocalMux I__2875 (
            .O(N__19423),
            .I(N__19412));
    LocalMux I__2874 (
            .O(N__19418),
            .I(N__19407));
    LocalMux I__2873 (
            .O(N__19415),
            .I(N__19407));
    Odrv4 I__2872 (
            .O(N__19412),
            .I(\b2v_inst11.N_357 ));
    Odrv12 I__2871 (
            .O(N__19407),
            .I(\b2v_inst11.N_357 ));
    InMux I__2870 (
            .O(N__19402),
            .I(N__19399));
    LocalMux I__2869 (
            .O(N__19399),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0 ));
    CascadeMux I__2868 (
            .O(N__19396),
            .I(N__19393));
    InMux I__2867 (
            .O(N__19393),
            .I(N__19390));
    LocalMux I__2866 (
            .O(N__19390),
            .I(N__19387));
    Odrv4 I__2865 (
            .O(N__19387),
            .I(\b2v_inst11.un1_func_state25_6_0_a2_0 ));
    InMux I__2864 (
            .O(N__19384),
            .I(N__19381));
    LocalMux I__2863 (
            .O(N__19381),
            .I(N__19378));
    Span4Mux_s3_v I__2862 (
            .O(N__19378),
            .I(N__19375));
    Odrv4 I__2861 (
            .O(N__19375),
            .I(\b2v_inst11.N_327 ));
    InMux I__2860 (
            .O(N__19372),
            .I(N__19369));
    LocalMux I__2859 (
            .O(N__19369),
            .I(N__19366));
    Span4Mux_s3_v I__2858 (
            .O(N__19366),
            .I(N__19363));
    Odrv4 I__2857 (
            .O(N__19363),
            .I(\b2v_inst11.N_328 ));
    CascadeMux I__2856 (
            .O(N__19360),
            .I(\b2v_inst11.func_state_1_m0_0_0_0_cascade_ ));
    InMux I__2855 (
            .O(N__19357),
            .I(N__19354));
    LocalMux I__2854 (
            .O(N__19354),
            .I(N__19351));
    Odrv12 I__2853 (
            .O(N__19351),
            .I(\b2v_inst11.N_354 ));
    CascadeMux I__2852 (
            .O(N__19348),
            .I(\b2v_inst11.N_354_cascade_ ));
    InMux I__2851 (
            .O(N__19345),
            .I(N__19341));
    CascadeMux I__2850 (
            .O(N__19344),
            .I(N__19334));
    LocalMux I__2849 (
            .O(N__19341),
            .I(N__19329));
    InMux I__2848 (
            .O(N__19340),
            .I(N__19323));
    InMux I__2847 (
            .O(N__19339),
            .I(N__19323));
    InMux I__2846 (
            .O(N__19338),
            .I(N__19320));
    InMux I__2845 (
            .O(N__19337),
            .I(N__19313));
    InMux I__2844 (
            .O(N__19334),
            .I(N__19313));
    InMux I__2843 (
            .O(N__19333),
            .I(N__19308));
    InMux I__2842 (
            .O(N__19332),
            .I(N__19308));
    Span4Mux_v I__2841 (
            .O(N__19329),
            .I(N__19305));
    InMux I__2840 (
            .O(N__19328),
            .I(N__19302));
    LocalMux I__2839 (
            .O(N__19323),
            .I(N__19297));
    LocalMux I__2838 (
            .O(N__19320),
            .I(N__19297));
    InMux I__2837 (
            .O(N__19319),
            .I(N__19292));
    InMux I__2836 (
            .O(N__19318),
            .I(N__19292));
    LocalMux I__2835 (
            .O(N__19313),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_11 ));
    LocalMux I__2834 (
            .O(N__19308),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_11 ));
    Odrv4 I__2833 (
            .O(N__19305),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_11 ));
    LocalMux I__2832 (
            .O(N__19302),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_11 ));
    Odrv4 I__2831 (
            .O(N__19297),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_11 ));
    LocalMux I__2830 (
            .O(N__19292),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_11 ));
    InMux I__2829 (
            .O(N__19279),
            .I(N__19276));
    LocalMux I__2828 (
            .O(N__19276),
            .I(\b2v_inst11.g2_1_1 ));
    CascadeMux I__2827 (
            .O(N__19273),
            .I(\b2v_inst11.g3_0_1_cascade_ ));
    InMux I__2826 (
            .O(N__19270),
            .I(N__19267));
    LocalMux I__2825 (
            .O(N__19267),
            .I(\b2v_inst11.N_14_0 ));
    InMux I__2824 (
            .O(N__19264),
            .I(N__19261));
    LocalMux I__2823 (
            .O(N__19261),
            .I(\b2v_inst11.dutycycle_RNI_6Z0Z_5 ));
    CascadeMux I__2822 (
            .O(N__19258),
            .I(\b2v_inst11.dutycycle_RNI_6Z0Z_5_cascade_ ));
    CascadeMux I__2821 (
            .O(N__19255),
            .I(\b2v_inst11.G_6_i_0_cascade_ ));
    InMux I__2820 (
            .O(N__19252),
            .I(N__19249));
    LocalMux I__2819 (
            .O(N__19249),
            .I(\b2v_inst11.G_6_i_a4_1_1 ));
    InMux I__2818 (
            .O(N__19246),
            .I(N__19243));
    LocalMux I__2817 (
            .O(N__19243),
            .I(\b2v_inst11.un1_dutycycle_53_7_1 ));
    CascadeMux I__2816 (
            .O(N__19240),
            .I(N__19236));
    InMux I__2815 (
            .O(N__19239),
            .I(N__19231));
    InMux I__2814 (
            .O(N__19236),
            .I(N__19231));
    LocalMux I__2813 (
            .O(N__19231),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    InMux I__2812 (
            .O(N__19228),
            .I(N__19222));
    InMux I__2811 (
            .O(N__19227),
            .I(N__19222));
    LocalMux I__2810 (
            .O(N__19222),
            .I(\b2v_inst11.dutycycle_RNIGKEF3Z0Z_11 ));
    CascadeMux I__2809 (
            .O(N__19219),
            .I(\b2v_inst11.dutycycleZ0Z_7_cascade_ ));
    CascadeMux I__2808 (
            .O(N__19216),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_ ));
    CascadeMux I__2807 (
            .O(N__19213),
            .I(N__19210));
    InMux I__2806 (
            .O(N__19210),
            .I(N__19207));
    LocalMux I__2805 (
            .O(N__19207),
            .I(N__19204));
    Odrv12 I__2804 (
            .O(N__19204),
            .I(\b2v_inst11.un1_dutycycle_53_8_0 ));
    InMux I__2803 (
            .O(N__19201),
            .I(N__19198));
    LocalMux I__2802 (
            .O(N__19198),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_11 ));
    CascadeMux I__2801 (
            .O(N__19195),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_7_cascade_ ));
    CascadeMux I__2800 (
            .O(N__19192),
            .I(N__19189));
    InMux I__2799 (
            .O(N__19189),
            .I(N__19186));
    LocalMux I__2798 (
            .O(N__19186),
            .I(N__19183));
    Odrv12 I__2797 (
            .O(N__19183),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_12 ));
    CascadeMux I__2796 (
            .O(N__19180),
            .I(\b2v_inst11.m18_i_1_0_cascade_ ));
    InMux I__2795 (
            .O(N__19177),
            .I(N__19174));
    LocalMux I__2794 (
            .O(N__19174),
            .I(N__19171));
    Odrv4 I__2793 (
            .O(N__19171),
            .I(\b2v_inst11.dutycycle_RNI_11Z0Z_9 ));
    InMux I__2792 (
            .O(N__19168),
            .I(N__19165));
    LocalMux I__2791 (
            .O(N__19165),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_7 ));
    InMux I__2790 (
            .O(N__19162),
            .I(N__19159));
    LocalMux I__2789 (
            .O(N__19159),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_7 ));
    CascadeMux I__2788 (
            .O(N__19156),
            .I(N__19151));
    CascadeMux I__2787 (
            .O(N__19155),
            .I(N__19147));
    CascadeMux I__2786 (
            .O(N__19154),
            .I(N__19144));
    InMux I__2785 (
            .O(N__19151),
            .I(N__19134));
    InMux I__2784 (
            .O(N__19150),
            .I(N__19134));
    InMux I__2783 (
            .O(N__19147),
            .I(N__19125));
    InMux I__2782 (
            .O(N__19144),
            .I(N__19125));
    InMux I__2781 (
            .O(N__19143),
            .I(N__19125));
    InMux I__2780 (
            .O(N__19142),
            .I(N__19125));
    InMux I__2779 (
            .O(N__19141),
            .I(N__19118));
    InMux I__2778 (
            .O(N__19140),
            .I(N__19118));
    InMux I__2777 (
            .O(N__19139),
            .I(N__19118));
    LocalMux I__2776 (
            .O(N__19134),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_9 ));
    LocalMux I__2775 (
            .O(N__19125),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_9 ));
    LocalMux I__2774 (
            .O(N__19118),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_9 ));
    InMux I__2773 (
            .O(N__19111),
            .I(N__19108));
    LocalMux I__2772 (
            .O(N__19108),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_7 ));
    InMux I__2771 (
            .O(N__19105),
            .I(N__19102));
    LocalMux I__2770 (
            .O(N__19102),
            .I(\b2v_inst11.dutycycle_RNI_8Z0Z_9 ));
    CascadeMux I__2769 (
            .O(N__19099),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_7_cascade_ ));
    CascadeMux I__2768 (
            .O(N__19096),
            .I(N__19093));
    InMux I__2767 (
            .O(N__19093),
            .I(N__19090));
    LocalMux I__2766 (
            .O(N__19090),
            .I(N__19087));
    Odrv12 I__2765 (
            .O(N__19087),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_11 ));
    InMux I__2764 (
            .O(N__19084),
            .I(N__19081));
    LocalMux I__2763 (
            .O(N__19081),
            .I(\b2v_inst11.un1_dutycycle_53_13_1 ));
    CascadeMux I__2762 (
            .O(N__19078),
            .I(\b2v_inst11.un1_dutycycle_53_39_0_0_1_cascade_ ));
    InMux I__2761 (
            .O(N__19075),
            .I(N__19072));
    LocalMux I__2760 (
            .O(N__19072),
            .I(\b2v_inst11.un1_dutycycle_53_39_0_0 ));
    CascadeMux I__2759 (
            .O(N__19069),
            .I(\b2v_inst11.un1_dutycycle_53_39_1_cascade_ ));
    InMux I__2758 (
            .O(N__19066),
            .I(N__19063));
    LocalMux I__2757 (
            .O(N__19063),
            .I(\b2v_inst11.un1_dutycycle_53_41_0 ));
    CascadeMux I__2756 (
            .O(N__19060),
            .I(N__19057));
    InMux I__2755 (
            .O(N__19057),
            .I(N__19054));
    LocalMux I__2754 (
            .O(N__19054),
            .I(N__19051));
    Odrv4 I__2753 (
            .O(N__19051),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_13 ));
    CascadeMux I__2752 (
            .O(N__19048),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_9_cascade_ ));
    CascadeMux I__2751 (
            .O(N__19045),
            .I(\b2v_inst11.un1_dutycycle_53_10_1_0_cascade_ ));
    CascadeMux I__2750 (
            .O(N__19042),
            .I(\b2v_inst11.un1_dutycycle_53_44_0_1_cascade_ ));
    CascadeMux I__2749 (
            .O(N__19039),
            .I(\b2v_inst11.dutycycle_RNI_6Z0Z_9_cascade_ ));
    CascadeMux I__2748 (
            .O(N__19036),
            .I(N__19033));
    InMux I__2747 (
            .O(N__19033),
            .I(N__19030));
    LocalMux I__2746 (
            .O(N__19030),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_11 ));
    CascadeMux I__2745 (
            .O(N__19027),
            .I(N__19024));
    InMux I__2744 (
            .O(N__19024),
            .I(N__19021));
    LocalMux I__2743 (
            .O(N__19021),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_15 ));
    CascadeMux I__2742 (
            .O(N__19018),
            .I(\b2v_inst11.un1_m7_1_0_cascade_ ));
    InMux I__2741 (
            .O(N__19015),
            .I(N__19012));
    LocalMux I__2740 (
            .O(N__19012),
            .I(N__19008));
    InMux I__2739 (
            .O(N__19011),
            .I(N__19005));
    Span4Mux_v I__2738 (
            .O(N__19008),
            .I(N__19002));
    LocalMux I__2737 (
            .O(N__19005),
            .I(\b2v_inst11.un1_i3_mux ));
    Odrv4 I__2736 (
            .O(N__19002),
            .I(\b2v_inst11.un1_i3_mux ));
    InMux I__2735 (
            .O(N__18997),
            .I(N__18994));
    LocalMux I__2734 (
            .O(N__18994),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_11 ));
    InMux I__2733 (
            .O(N__18991),
            .I(N__18988));
    LocalMux I__2732 (
            .O(N__18988),
            .I(\b2v_inst11.un1_dutycycle_53_44_0_2_tz ));
    InMux I__2731 (
            .O(N__18985),
            .I(\b2v_inst11.un1_dutycycle_53_cry_11 ));
    CascadeMux I__2730 (
            .O(N__18982),
            .I(N__18979));
    InMux I__2729 (
            .O(N__18979),
            .I(N__18976));
    LocalMux I__2728 (
            .O(N__18976),
            .I(N__18973));
    Span4Mux_v I__2727 (
            .O(N__18973),
            .I(N__18970));
    Odrv4 I__2726 (
            .O(N__18970),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_13 ));
    InMux I__2725 (
            .O(N__18967),
            .I(\b2v_inst11.un1_dutycycle_53_cry_12 ));
    InMux I__2724 (
            .O(N__18964),
            .I(N__18961));
    LocalMux I__2723 (
            .O(N__18961),
            .I(N__18958));
    Odrv4 I__2722 (
            .O(N__18958),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_13 ));
    CascadeMux I__2721 (
            .O(N__18955),
            .I(N__18952));
    InMux I__2720 (
            .O(N__18952),
            .I(N__18948));
    InMux I__2719 (
            .O(N__18951),
            .I(N__18945));
    LocalMux I__2718 (
            .O(N__18948),
            .I(N__18942));
    LocalMux I__2717 (
            .O(N__18945),
            .I(\b2v_inst11.mult1_un47_sum ));
    Odrv4 I__2716 (
            .O(N__18942),
            .I(\b2v_inst11.mult1_un47_sum ));
    InMux I__2715 (
            .O(N__18937),
            .I(\b2v_inst11.un1_dutycycle_53_cry_13 ));
    InMux I__2714 (
            .O(N__18934),
            .I(N__18931));
    LocalMux I__2713 (
            .O(N__18931),
            .I(N__18928));
    Span4Mux_h I__2712 (
            .O(N__18928),
            .I(N__18922));
    InMux I__2711 (
            .O(N__18927),
            .I(N__18915));
    InMux I__2710 (
            .O(N__18926),
            .I(N__18915));
    InMux I__2709 (
            .O(N__18925),
            .I(N__18915));
    Odrv4 I__2708 (
            .O(N__18922),
            .I(\b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0 ));
    LocalMux I__2707 (
            .O(N__18915),
            .I(\b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0 ));
    InMux I__2706 (
            .O(N__18910),
            .I(\b2v_inst11.un1_dutycycle_53_cry_14 ));
    CascadeMux I__2705 (
            .O(N__18907),
            .I(N__18904));
    InMux I__2704 (
            .O(N__18904),
            .I(N__18901));
    LocalMux I__2703 (
            .O(N__18901),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_14 ));
    InMux I__2702 (
            .O(N__18898),
            .I(N__18893));
    CascadeMux I__2701 (
            .O(N__18897),
            .I(N__18890));
    CascadeMux I__2700 (
            .O(N__18896),
            .I(N__18887));
    LocalMux I__2699 (
            .O(N__18893),
            .I(N__18884));
    InMux I__2698 (
            .O(N__18890),
            .I(N__18879));
    InMux I__2697 (
            .O(N__18887),
            .I(N__18879));
    Span4Mux_h I__2696 (
            .O(N__18884),
            .I(N__18874));
    LocalMux I__2695 (
            .O(N__18879),
            .I(N__18874));
    Odrv4 I__2694 (
            .O(N__18874),
            .I(\b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ));
    InMux I__2693 (
            .O(N__18871),
            .I(bfn_5_9_0_));
    InMux I__2692 (
            .O(N__18868),
            .I(\b2v_inst11.CO2 ));
    CascadeMux I__2691 (
            .O(N__18865),
            .I(N__18862));
    InMux I__2690 (
            .O(N__18862),
            .I(N__18859));
    LocalMux I__2689 (
            .O(N__18859),
            .I(N__18855));
    InMux I__2688 (
            .O(N__18858),
            .I(N__18852));
    Span4Mux_h I__2687 (
            .O(N__18855),
            .I(N__18847));
    LocalMux I__2686 (
            .O(N__18852),
            .I(N__18847));
    Odrv4 I__2685 (
            .O(N__18847),
            .I(\b2v_inst11.CO2_THRU_CO ));
    InMux I__2684 (
            .O(N__18844),
            .I(N__18841));
    LocalMux I__2683 (
            .O(N__18841),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_10 ));
    InMux I__2682 (
            .O(N__18838),
            .I(N__18835));
    LocalMux I__2681 (
            .O(N__18835),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_15 ));
    InMux I__2680 (
            .O(N__18832),
            .I(\b2v_inst11.un1_dutycycle_53_cry_2_cZ0 ));
    InMux I__2679 (
            .O(N__18829),
            .I(\b2v_inst11.un1_dutycycle_53_cry_3_cZ0 ));
    InMux I__2678 (
            .O(N__18826),
            .I(N__18822));
    InMux I__2677 (
            .O(N__18825),
            .I(N__18819));
    LocalMux I__2676 (
            .O(N__18822),
            .I(N__18814));
    LocalMux I__2675 (
            .O(N__18819),
            .I(N__18814));
    Odrv12 I__2674 (
            .O(N__18814),
            .I(\b2v_inst11.mult1_un110_sum ));
    InMux I__2673 (
            .O(N__18811),
            .I(\b2v_inst11.un1_dutycycle_53_cry_4_cZ0 ));
    InMux I__2672 (
            .O(N__18808),
            .I(N__18804));
    InMux I__2671 (
            .O(N__18807),
            .I(N__18801));
    LocalMux I__2670 (
            .O(N__18804),
            .I(N__18796));
    LocalMux I__2669 (
            .O(N__18801),
            .I(N__18796));
    Odrv12 I__2668 (
            .O(N__18796),
            .I(\b2v_inst11.mult1_un103_sum ));
    InMux I__2667 (
            .O(N__18793),
            .I(\b2v_inst11.un1_dutycycle_53_cry_5_cZ0 ));
    InMux I__2666 (
            .O(N__18790),
            .I(N__18787));
    LocalMux I__2665 (
            .O(N__18787),
            .I(N__18784));
    Span4Mux_s3_v I__2664 (
            .O(N__18784),
            .I(N__18780));
    InMux I__2663 (
            .O(N__18783),
            .I(N__18777));
    Odrv4 I__2662 (
            .O(N__18780),
            .I(\b2v_inst11.mult1_un96_sum ));
    LocalMux I__2661 (
            .O(N__18777),
            .I(\b2v_inst11.mult1_un96_sum ));
    InMux I__2660 (
            .O(N__18772),
            .I(\b2v_inst11.un1_dutycycle_53_cry_6_cZ0 ));
    InMux I__2659 (
            .O(N__18769),
            .I(bfn_5_8_0_));
    InMux I__2658 (
            .O(N__18766),
            .I(N__18763));
    LocalMux I__2657 (
            .O(N__18763),
            .I(N__18759));
    InMux I__2656 (
            .O(N__18762),
            .I(N__18756));
    Sp12to4 I__2655 (
            .O(N__18759),
            .I(N__18751));
    LocalMux I__2654 (
            .O(N__18756),
            .I(N__18751));
    Odrv12 I__2653 (
            .O(N__18751),
            .I(\b2v_inst11.mult1_un82_sum ));
    InMux I__2652 (
            .O(N__18748),
            .I(\b2v_inst11.un1_dutycycle_53_cry_8_cZ0 ));
    InMux I__2651 (
            .O(N__18745),
            .I(N__18742));
    LocalMux I__2650 (
            .O(N__18742),
            .I(N__18738));
    InMux I__2649 (
            .O(N__18741),
            .I(N__18735));
    Sp12to4 I__2648 (
            .O(N__18738),
            .I(N__18730));
    LocalMux I__2647 (
            .O(N__18735),
            .I(N__18730));
    Odrv12 I__2646 (
            .O(N__18730),
            .I(\b2v_inst11.mult1_un75_sum ));
    InMux I__2645 (
            .O(N__18727),
            .I(\b2v_inst11.un1_dutycycle_53_cry_9_cZ0 ));
    InMux I__2644 (
            .O(N__18724),
            .I(\b2v_inst11.un1_dutycycle_53_cry_10 ));
    CascadeMux I__2643 (
            .O(N__18721),
            .I(N__18718));
    InMux I__2642 (
            .O(N__18718),
            .I(N__18715));
    LocalMux I__2641 (
            .O(N__18715),
            .I(\b2v_inst11.mult1_un47_sum_cry_4_s ));
    CascadeMux I__2640 (
            .O(N__18712),
            .I(N__18709));
    InMux I__2639 (
            .O(N__18709),
            .I(N__18706));
    LocalMux I__2638 (
            .O(N__18706),
            .I(\b2v_inst11.mult1_un54_sum_cry_5_s ));
    InMux I__2637 (
            .O(N__18703),
            .I(\b2v_inst11.mult1_un54_sum_cry_4 ));
    CascadeMux I__2636 (
            .O(N__18700),
            .I(N__18697));
    InMux I__2635 (
            .O(N__18697),
            .I(N__18694));
    LocalMux I__2634 (
            .O(N__18694),
            .I(\b2v_inst11.mult1_un47_sum_cry_5_s ));
    InMux I__2633 (
            .O(N__18691),
            .I(N__18688));
    LocalMux I__2632 (
            .O(N__18688),
            .I(\b2v_inst11.mult1_un54_sum_cry_6_s ));
    InMux I__2631 (
            .O(N__18685),
            .I(\b2v_inst11.mult1_un54_sum_cry_5 ));
    InMux I__2630 (
            .O(N__18682),
            .I(N__18679));
    LocalMux I__2629 (
            .O(N__18679),
            .I(\b2v_inst11.mult1_un47_sum_l_fx_6 ));
    CascadeMux I__2628 (
            .O(N__18676),
            .I(N__18673));
    InMux I__2627 (
            .O(N__18673),
            .I(N__18668));
    InMux I__2626 (
            .O(N__18672),
            .I(N__18665));
    InMux I__2625 (
            .O(N__18671),
            .I(N__18662));
    LocalMux I__2624 (
            .O(N__18668),
            .I(\b2v_inst11.mult1_un47_sum_s_6 ));
    LocalMux I__2623 (
            .O(N__18665),
            .I(\b2v_inst11.mult1_un47_sum_s_6 ));
    LocalMux I__2622 (
            .O(N__18662),
            .I(\b2v_inst11.mult1_un47_sum_s_6 ));
    CascadeMux I__2621 (
            .O(N__18655),
            .I(N__18652));
    InMux I__2620 (
            .O(N__18652),
            .I(N__18649));
    LocalMux I__2619 (
            .O(N__18649),
            .I(\b2v_inst11.mult1_un61_sum_axb_8 ));
    InMux I__2618 (
            .O(N__18646),
            .I(\b2v_inst11.mult1_un54_sum_cry_6 ));
    InMux I__2617 (
            .O(N__18643),
            .I(N__18640));
    LocalMux I__2616 (
            .O(N__18640),
            .I(\b2v_inst11.mult1_un40_sum_i_5 ));
    CascadeMux I__2615 (
            .O(N__18637),
            .I(N__18634));
    InMux I__2614 (
            .O(N__18634),
            .I(N__18630));
    InMux I__2613 (
            .O(N__18633),
            .I(N__18627));
    LocalMux I__2612 (
            .O(N__18630),
            .I(\b2v_inst11.mult1_un47_sum_cry_5_THRU_CO ));
    LocalMux I__2611 (
            .O(N__18627),
            .I(\b2v_inst11.mult1_un47_sum_cry_5_THRU_CO ));
    InMux I__2610 (
            .O(N__18622),
            .I(\b2v_inst11.mult1_un54_sum_cry_7 ));
    CascadeMux I__2609 (
            .O(N__18619),
            .I(N__18615));
    InMux I__2608 (
            .O(N__18618),
            .I(N__18609));
    InMux I__2607 (
            .O(N__18615),
            .I(N__18609));
    InMux I__2606 (
            .O(N__18614),
            .I(N__18606));
    LocalMux I__2605 (
            .O(N__18609),
            .I(\b2v_inst11.mult1_un54_sum_s_8 ));
    LocalMux I__2604 (
            .O(N__18606),
            .I(\b2v_inst11.mult1_un54_sum_s_8 ));
    CascadeMux I__2603 (
            .O(N__18601),
            .I(\b2v_inst11.mult1_un54_sum_s_8_cascade_ ));
    CascadeMux I__2602 (
            .O(N__18598),
            .I(N__18594));
    CascadeMux I__2601 (
            .O(N__18597),
            .I(N__18590));
    InMux I__2600 (
            .O(N__18594),
            .I(N__18583));
    InMux I__2599 (
            .O(N__18593),
            .I(N__18583));
    InMux I__2598 (
            .O(N__18590),
            .I(N__18583));
    LocalMux I__2597 (
            .O(N__18583),
            .I(\b2v_inst11.mult1_un54_sum_i_8 ));
    InMux I__2596 (
            .O(N__18580),
            .I(N__18577));
    LocalMux I__2595 (
            .O(N__18577),
            .I(N__18574));
    Span4Mux_v I__2594 (
            .O(N__18574),
            .I(N__18571));
    Odrv4 I__2593 (
            .O(N__18571),
            .I(\b2v_inst11.m15_e_2 ));
    InMux I__2592 (
            .O(N__18568),
            .I(\b2v_inst11.un1_dutycycle_53_cry_0_cZ0 ));
    InMux I__2591 (
            .O(N__18565),
            .I(\b2v_inst11.un1_dutycycle_53_cry_1_cZ0 ));
    InMux I__2590 (
            .O(N__18562),
            .I(N__18559));
    LocalMux I__2589 (
            .O(N__18559),
            .I(\b2v_inst11.mult1_un61_sum_cry_4_s ));
    InMux I__2588 (
            .O(N__18556),
            .I(\b2v_inst11.mult1_un61_sum_cry_3 ));
    InMux I__2587 (
            .O(N__18553),
            .I(N__18550));
    LocalMux I__2586 (
            .O(N__18550),
            .I(\b2v_inst11.mult1_un61_sum_cry_5_s ));
    InMux I__2585 (
            .O(N__18547),
            .I(\b2v_inst11.mult1_un61_sum_cry_4 ));
    CascadeMux I__2584 (
            .O(N__18544),
            .I(N__18541));
    InMux I__2583 (
            .O(N__18541),
            .I(N__18538));
    LocalMux I__2582 (
            .O(N__18538),
            .I(\b2v_inst11.mult1_un61_sum_cry_6_s ));
    InMux I__2581 (
            .O(N__18535),
            .I(\b2v_inst11.mult1_un61_sum_cry_5 ));
    InMux I__2580 (
            .O(N__18532),
            .I(N__18529));
    LocalMux I__2579 (
            .O(N__18529),
            .I(\b2v_inst11.mult1_un68_sum_axb_8 ));
    InMux I__2578 (
            .O(N__18526),
            .I(\b2v_inst11.mult1_un61_sum_cry_6 ));
    InMux I__2577 (
            .O(N__18523),
            .I(\b2v_inst11.mult1_un61_sum_cry_7 ));
    InMux I__2576 (
            .O(N__18520),
            .I(N__18517));
    LocalMux I__2575 (
            .O(N__18517),
            .I(\b2v_inst11.mult1_un47_sum_i ));
    CascadeMux I__2574 (
            .O(N__18514),
            .I(N__18511));
    InMux I__2573 (
            .O(N__18511),
            .I(N__18508));
    LocalMux I__2572 (
            .O(N__18508),
            .I(\b2v_inst11.mult1_un54_sum_cry_3_s ));
    InMux I__2571 (
            .O(N__18505),
            .I(\b2v_inst11.mult1_un54_sum_cry_2 ));
    InMux I__2570 (
            .O(N__18502),
            .I(N__18497));
    InMux I__2569 (
            .O(N__18501),
            .I(N__18494));
    InMux I__2568 (
            .O(N__18500),
            .I(N__18491));
    LocalMux I__2567 (
            .O(N__18497),
            .I(\b2v_inst11.mult1_un47_sum_cry_3_s ));
    LocalMux I__2566 (
            .O(N__18494),
            .I(\b2v_inst11.mult1_un47_sum_cry_3_s ));
    LocalMux I__2565 (
            .O(N__18491),
            .I(\b2v_inst11.mult1_un47_sum_cry_3_s ));
    CascadeMux I__2564 (
            .O(N__18484),
            .I(N__18481));
    InMux I__2563 (
            .O(N__18481),
            .I(N__18478));
    LocalMux I__2562 (
            .O(N__18478),
            .I(\b2v_inst11.mult1_un47_sum_l_fx_3 ));
    InMux I__2561 (
            .O(N__18475),
            .I(N__18472));
    LocalMux I__2560 (
            .O(N__18472),
            .I(\b2v_inst11.mult1_un54_sum_cry_4_s ));
    InMux I__2559 (
            .O(N__18469),
            .I(\b2v_inst11.mult1_un54_sum_cry_3 ));
    InMux I__2558 (
            .O(N__18466),
            .I(N__18463));
    LocalMux I__2557 (
            .O(N__18463),
            .I(\b2v_inst11.mult1_un68_sum_cry_3_s ));
    InMux I__2556 (
            .O(N__18460),
            .I(\b2v_inst11.mult1_un68_sum_cry_2_c ));
    CascadeMux I__2555 (
            .O(N__18457),
            .I(N__18454));
    InMux I__2554 (
            .O(N__18454),
            .I(N__18451));
    LocalMux I__2553 (
            .O(N__18451),
            .I(\b2v_inst11.mult1_un68_sum_cry_4_s ));
    InMux I__2552 (
            .O(N__18448),
            .I(\b2v_inst11.mult1_un68_sum_cry_3_c ));
    InMux I__2551 (
            .O(N__18445),
            .I(N__18442));
    LocalMux I__2550 (
            .O(N__18442),
            .I(\b2v_inst11.mult1_un68_sum_cry_5_s ));
    InMux I__2549 (
            .O(N__18439),
            .I(\b2v_inst11.mult1_un68_sum_cry_4_c ));
    CascadeMux I__2548 (
            .O(N__18436),
            .I(N__18433));
    InMux I__2547 (
            .O(N__18433),
            .I(N__18430));
    LocalMux I__2546 (
            .O(N__18430),
            .I(\b2v_inst11.mult1_un68_sum_cry_6_s ));
    InMux I__2545 (
            .O(N__18427),
            .I(\b2v_inst11.mult1_un68_sum_cry_5_c ));
    InMux I__2544 (
            .O(N__18424),
            .I(N__18421));
    LocalMux I__2543 (
            .O(N__18421),
            .I(\b2v_inst11.mult1_un75_sum_axb_8 ));
    InMux I__2542 (
            .O(N__18418),
            .I(\b2v_inst11.mult1_un68_sum_cry_6_c ));
    InMux I__2541 (
            .O(N__18415),
            .I(\b2v_inst11.mult1_un68_sum_cry_7 ));
    CascadeMux I__2540 (
            .O(N__18412),
            .I(\b2v_inst11.mult1_un68_sum_s_8_cascade_ ));
    CascadeMux I__2539 (
            .O(N__18409),
            .I(N__18405));
    InMux I__2538 (
            .O(N__18408),
            .I(N__18397));
    InMux I__2537 (
            .O(N__18405),
            .I(N__18397));
    InMux I__2536 (
            .O(N__18404),
            .I(N__18397));
    LocalMux I__2535 (
            .O(N__18397),
            .I(\b2v_inst11.mult1_un68_sum_i_0_8 ));
    InMux I__2534 (
            .O(N__18394),
            .I(N__18391));
    LocalMux I__2533 (
            .O(N__18391),
            .I(\b2v_inst11.mult1_un61_sum_cry_3_s ));
    InMux I__2532 (
            .O(N__18388),
            .I(\b2v_inst11.mult1_un61_sum_cry_2 ));
    CascadeMux I__2531 (
            .O(N__18385),
            .I(N__18382));
    InMux I__2530 (
            .O(N__18382),
            .I(N__18379));
    LocalMux I__2529 (
            .O(N__18379),
            .I(\b2v_inst11.mult1_un82_sum_i ));
    CascadeMux I__2528 (
            .O(N__18376),
            .I(N__18373));
    InMux I__2527 (
            .O(N__18373),
            .I(N__18370));
    LocalMux I__2526 (
            .O(N__18370),
            .I(\b2v_inst11.mult1_un75_sum_i ));
    CascadeMux I__2525 (
            .O(N__18367),
            .I(N__18364));
    InMux I__2524 (
            .O(N__18364),
            .I(N__18361));
    LocalMux I__2523 (
            .O(N__18361),
            .I(N__18358));
    Odrv12 I__2522 (
            .O(N__18358),
            .I(\b2v_inst11.mult1_un103_sum_i ));
    CascadeMux I__2521 (
            .O(N__18355),
            .I(N__18352));
    InMux I__2520 (
            .O(N__18352),
            .I(N__18344));
    InMux I__2519 (
            .O(N__18351),
            .I(N__18344));
    InMux I__2518 (
            .O(N__18350),
            .I(N__18341));
    InMux I__2517 (
            .O(N__18349),
            .I(N__18338));
    LocalMux I__2516 (
            .O(N__18344),
            .I(\b2v_inst11.mult1_un103_sum_s_8 ));
    LocalMux I__2515 (
            .O(N__18341),
            .I(\b2v_inst11.mult1_un103_sum_s_8 ));
    LocalMux I__2514 (
            .O(N__18338),
            .I(\b2v_inst11.mult1_un103_sum_s_8 ));
    CascadeMux I__2513 (
            .O(N__18331),
            .I(N__18328));
    InMux I__2512 (
            .O(N__18328),
            .I(N__18319));
    InMux I__2511 (
            .O(N__18327),
            .I(N__18319));
    InMux I__2510 (
            .O(N__18326),
            .I(N__18319));
    LocalMux I__2509 (
            .O(N__18319),
            .I(\b2v_inst11.mult1_un89_sum_i_0_8 ));
    CascadeMux I__2508 (
            .O(N__18316),
            .I(N__18313));
    InMux I__2507 (
            .O(N__18313),
            .I(N__18310));
    LocalMux I__2506 (
            .O(N__18310),
            .I(N__18307));
    Span4Mux_s3_v I__2505 (
            .O(N__18307),
            .I(N__18304));
    Span4Mux_v I__2504 (
            .O(N__18304),
            .I(N__18301));
    Odrv4 I__2503 (
            .O(N__18301),
            .I(\b2v_inst11.mult1_un96_sum_i ));
    InMux I__2502 (
            .O(N__18298),
            .I(N__18295));
    LocalMux I__2501 (
            .O(N__18295),
            .I(\b2v_inst11.mult1_un103_sum_cry_3_s ));
    InMux I__2500 (
            .O(N__18292),
            .I(\b2v_inst11.mult1_un103_sum_cry_2 ));
    InMux I__2499 (
            .O(N__18289),
            .I(N__18286));
    LocalMux I__2498 (
            .O(N__18286),
            .I(\b2v_inst11.mult1_un96_sum_cry_3_s ));
    CascadeMux I__2497 (
            .O(N__18283),
            .I(N__18280));
    InMux I__2496 (
            .O(N__18280),
            .I(N__18277));
    LocalMux I__2495 (
            .O(N__18277),
            .I(\b2v_inst11.mult1_un103_sum_cry_4_s ));
    InMux I__2494 (
            .O(N__18274),
            .I(\b2v_inst11.mult1_un103_sum_cry_3 ));
    CascadeMux I__2493 (
            .O(N__18271),
            .I(N__18268));
    InMux I__2492 (
            .O(N__18268),
            .I(N__18265));
    LocalMux I__2491 (
            .O(N__18265),
            .I(\b2v_inst11.mult1_un96_sum_cry_4_s ));
    InMux I__2490 (
            .O(N__18262),
            .I(N__18259));
    LocalMux I__2489 (
            .O(N__18259),
            .I(\b2v_inst11.mult1_un103_sum_cry_5_s ));
    InMux I__2488 (
            .O(N__18256),
            .I(\b2v_inst11.mult1_un103_sum_cry_4 ));
    InMux I__2487 (
            .O(N__18253),
            .I(N__18250));
    LocalMux I__2486 (
            .O(N__18250),
            .I(\b2v_inst11.mult1_un96_sum_cry_5_s ));
    CascadeMux I__2485 (
            .O(N__18247),
            .I(N__18244));
    InMux I__2484 (
            .O(N__18244),
            .I(N__18241));
    LocalMux I__2483 (
            .O(N__18241),
            .I(\b2v_inst11.mult1_un103_sum_cry_6_s ));
    InMux I__2482 (
            .O(N__18238),
            .I(\b2v_inst11.mult1_un103_sum_cry_5 ));
    CascadeMux I__2481 (
            .O(N__18235),
            .I(N__18231));
    InMux I__2480 (
            .O(N__18234),
            .I(N__18223));
    InMux I__2479 (
            .O(N__18231),
            .I(N__18223));
    InMux I__2478 (
            .O(N__18230),
            .I(N__18223));
    LocalMux I__2477 (
            .O(N__18223),
            .I(\b2v_inst11.mult1_un96_sum_i_0_8 ));
    CascadeMux I__2476 (
            .O(N__18220),
            .I(N__18217));
    InMux I__2475 (
            .O(N__18217),
            .I(N__18214));
    LocalMux I__2474 (
            .O(N__18214),
            .I(\b2v_inst11.mult1_un96_sum_cry_6_s ));
    InMux I__2473 (
            .O(N__18211),
            .I(N__18208));
    LocalMux I__2472 (
            .O(N__18208),
            .I(\b2v_inst11.mult1_un110_sum_axb_8 ));
    InMux I__2471 (
            .O(N__18205),
            .I(\b2v_inst11.mult1_un103_sum_cry_6 ));
    InMux I__2470 (
            .O(N__18202),
            .I(N__18199));
    LocalMux I__2469 (
            .O(N__18199),
            .I(\b2v_inst11.mult1_un103_sum_axb_8 ));
    InMux I__2468 (
            .O(N__18196),
            .I(\b2v_inst11.mult1_un103_sum_cry_7 ));
    CascadeMux I__2467 (
            .O(N__18193),
            .I(\b2v_inst11.mult1_un103_sum_s_8_cascade_ ));
    CascadeMux I__2466 (
            .O(N__18190),
            .I(N__18186));
    InMux I__2465 (
            .O(N__18189),
            .I(N__18178));
    InMux I__2464 (
            .O(N__18186),
            .I(N__18178));
    InMux I__2463 (
            .O(N__18185),
            .I(N__18178));
    LocalMux I__2462 (
            .O(N__18178),
            .I(\b2v_inst11.mult1_un103_sum_i_0_8 ));
    CascadeMux I__2461 (
            .O(N__18175),
            .I(N__18172));
    InMux I__2460 (
            .O(N__18172),
            .I(N__18169));
    LocalMux I__2459 (
            .O(N__18169),
            .I(N__18166));
    Odrv4 I__2458 (
            .O(N__18166),
            .I(\b2v_inst11.count_off_0_13 ));
    CascadeMux I__2457 (
            .O(N__18163),
            .I(N__18159));
    InMux I__2456 (
            .O(N__18162),
            .I(N__18144));
    InMux I__2455 (
            .O(N__18159),
            .I(N__18144));
    CEMux I__2454 (
            .O(N__18158),
            .I(N__18144));
    CascadeMux I__2453 (
            .O(N__18157),
            .I(N__18140));
    CEMux I__2452 (
            .O(N__18156),
            .I(N__18127));
    InMux I__2451 (
            .O(N__18155),
            .I(N__18120));
    InMux I__2450 (
            .O(N__18154),
            .I(N__18120));
    CEMux I__2449 (
            .O(N__18153),
            .I(N__18120));
    InMux I__2448 (
            .O(N__18152),
            .I(N__18115));
    CEMux I__2447 (
            .O(N__18151),
            .I(N__18115));
    LocalMux I__2446 (
            .O(N__18144),
            .I(N__18112));
    InMux I__2445 (
            .O(N__18143),
            .I(N__18109));
    InMux I__2444 (
            .O(N__18140),
            .I(N__18106));
    InMux I__2443 (
            .O(N__18139),
            .I(N__18103));
    InMux I__2442 (
            .O(N__18138),
            .I(N__18097));
    InMux I__2441 (
            .O(N__18137),
            .I(N__18094));
    InMux I__2440 (
            .O(N__18136),
            .I(N__18083));
    CEMux I__2439 (
            .O(N__18135),
            .I(N__18083));
    InMux I__2438 (
            .O(N__18134),
            .I(N__18083));
    InMux I__2437 (
            .O(N__18133),
            .I(N__18083));
    InMux I__2436 (
            .O(N__18132),
            .I(N__18083));
    InMux I__2435 (
            .O(N__18131),
            .I(N__18078));
    InMux I__2434 (
            .O(N__18130),
            .I(N__18078));
    LocalMux I__2433 (
            .O(N__18127),
            .I(N__18074));
    LocalMux I__2432 (
            .O(N__18120),
            .I(N__18071));
    LocalMux I__2431 (
            .O(N__18115),
            .I(N__18068));
    Span4Mux_s2_v I__2430 (
            .O(N__18112),
            .I(N__18065));
    LocalMux I__2429 (
            .O(N__18109),
            .I(N__18062));
    LocalMux I__2428 (
            .O(N__18106),
            .I(N__18057));
    LocalMux I__2427 (
            .O(N__18103),
            .I(N__18057));
    InMux I__2426 (
            .O(N__18102),
            .I(N__18050));
    InMux I__2425 (
            .O(N__18101),
            .I(N__18050));
    InMux I__2424 (
            .O(N__18100),
            .I(N__18050));
    LocalMux I__2423 (
            .O(N__18097),
            .I(N__18047));
    LocalMux I__2422 (
            .O(N__18094),
            .I(N__18042));
    LocalMux I__2421 (
            .O(N__18083),
            .I(N__18042));
    LocalMux I__2420 (
            .O(N__18078),
            .I(N__18039));
    CascadeMux I__2419 (
            .O(N__18077),
            .I(N__18034));
    Span4Mux_s3_h I__2418 (
            .O(N__18074),
            .I(N__18030));
    Span4Mux_h I__2417 (
            .O(N__18071),
            .I(N__18027));
    Span4Mux_s2_h I__2416 (
            .O(N__18068),
            .I(N__18018));
    Span4Mux_s2_h I__2415 (
            .O(N__18065),
            .I(N__18018));
    Span4Mux_s2_v I__2414 (
            .O(N__18062),
            .I(N__18018));
    Span4Mux_s2_v I__2413 (
            .O(N__18057),
            .I(N__18018));
    LocalMux I__2412 (
            .O(N__18050),
            .I(N__18011));
    Span4Mux_v I__2411 (
            .O(N__18047),
            .I(N__18011));
    Span4Mux_s2_v I__2410 (
            .O(N__18042),
            .I(N__18011));
    Span4Mux_s3_h I__2409 (
            .O(N__18039),
            .I(N__18008));
    InMux I__2408 (
            .O(N__18038),
            .I(N__17999));
    CEMux I__2407 (
            .O(N__18037),
            .I(N__17999));
    InMux I__2406 (
            .O(N__18034),
            .I(N__17999));
    InMux I__2405 (
            .O(N__18033),
            .I(N__17999));
    Odrv4 I__2404 (
            .O(N__18030),
            .I(\b2v_inst11.count_off_enZ0 ));
    Odrv4 I__2403 (
            .O(N__18027),
            .I(\b2v_inst11.count_off_enZ0 ));
    Odrv4 I__2402 (
            .O(N__18018),
            .I(\b2v_inst11.count_off_enZ0 ));
    Odrv4 I__2401 (
            .O(N__18011),
            .I(\b2v_inst11.count_off_enZ0 ));
    Odrv4 I__2400 (
            .O(N__18008),
            .I(\b2v_inst11.count_off_enZ0 ));
    LocalMux I__2399 (
            .O(N__17999),
            .I(\b2v_inst11.count_off_enZ0 ));
    InMux I__2398 (
            .O(N__17986),
            .I(N__17983));
    LocalMux I__2397 (
            .O(N__17983),
            .I(N__17980));
    Odrv12 I__2396 (
            .O(N__17980),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2 ));
    InMux I__2395 (
            .O(N__17977),
            .I(\b2v_inst11.mult1_un110_sum_cry_2 ));
    InMux I__2394 (
            .O(N__17974),
            .I(\b2v_inst11.mult1_un110_sum_cry_3 ));
    InMux I__2393 (
            .O(N__17971),
            .I(\b2v_inst11.mult1_un110_sum_cry_4 ));
    InMux I__2392 (
            .O(N__17968),
            .I(\b2v_inst11.mult1_un110_sum_cry_5 ));
    InMux I__2391 (
            .O(N__17965),
            .I(\b2v_inst11.mult1_un110_sum_cry_6 ));
    InMux I__2390 (
            .O(N__17962),
            .I(\b2v_inst11.mult1_un110_sum_cry_7 ));
    CascadeMux I__2389 (
            .O(N__17959),
            .I(N__17955));
    InMux I__2388 (
            .O(N__17958),
            .I(N__17949));
    InMux I__2387 (
            .O(N__17955),
            .I(N__17944));
    InMux I__2386 (
            .O(N__17954),
            .I(N__17944));
    InMux I__2385 (
            .O(N__17953),
            .I(N__17941));
    InMux I__2384 (
            .O(N__17952),
            .I(N__17938));
    LocalMux I__2383 (
            .O(N__17949),
            .I(\b2v_inst11.mult1_un89_sum_s_8 ));
    LocalMux I__2382 (
            .O(N__17944),
            .I(\b2v_inst11.mult1_un89_sum_s_8 ));
    LocalMux I__2381 (
            .O(N__17941),
            .I(\b2v_inst11.mult1_un89_sum_s_8 ));
    LocalMux I__2380 (
            .O(N__17938),
            .I(\b2v_inst11.mult1_un89_sum_s_8 ));
    InMux I__2379 (
            .O(N__17929),
            .I(N__17926));
    LocalMux I__2378 (
            .O(N__17926),
            .I(N__17923));
    Span4Mux_s2_h I__2377 (
            .O(N__17923),
            .I(N__17920));
    Span4Mux_v I__2376 (
            .O(N__17920),
            .I(N__17917));
    Odrv4 I__2375 (
            .O(N__17917),
            .I(\b2v_inst11.N_322 ));
    CascadeMux I__2374 (
            .O(N__17914),
            .I(\b2v_inst11.count_offZ0Z_0_cascade_ ));
    InMux I__2373 (
            .O(N__17911),
            .I(N__17907));
    CascadeMux I__2372 (
            .O(N__17910),
            .I(N__17904));
    LocalMux I__2371 (
            .O(N__17907),
            .I(N__17901));
    InMux I__2370 (
            .O(N__17904),
            .I(N__17898));
    Span4Mux_v I__2369 (
            .O(N__17901),
            .I(N__17894));
    LocalMux I__2368 (
            .O(N__17898),
            .I(N__17891));
    InMux I__2367 (
            .O(N__17897),
            .I(N__17888));
    Span4Mux_s1_v I__2366 (
            .O(N__17894),
            .I(N__17883));
    Span4Mux_v I__2365 (
            .O(N__17891),
            .I(N__17883));
    LocalMux I__2364 (
            .O(N__17888),
            .I(\b2v_inst11.count_offZ0Z_1 ));
    Odrv4 I__2363 (
            .O(N__17883),
            .I(\b2v_inst11.count_offZ0Z_1 ));
    InMux I__2362 (
            .O(N__17878),
            .I(N__17875));
    LocalMux I__2361 (
            .O(N__17875),
            .I(\b2v_inst11.count_off_RNIZ0Z_1 ));
    CascadeMux I__2360 (
            .O(N__17872),
            .I(\b2v_inst11.count_off_RNIZ0Z_1_cascade_ ));
    InMux I__2359 (
            .O(N__17869),
            .I(N__17866));
    LocalMux I__2358 (
            .O(N__17866),
            .I(\b2v_inst11.count_off_0_1 ));
    InMux I__2357 (
            .O(N__17863),
            .I(N__17859));
    InMux I__2356 (
            .O(N__17862),
            .I(N__17856));
    LocalMux I__2355 (
            .O(N__17859),
            .I(N__17853));
    LocalMux I__2354 (
            .O(N__17856),
            .I(N__17849));
    Span4Mux_v I__2353 (
            .O(N__17853),
            .I(N__17846));
    CascadeMux I__2352 (
            .O(N__17852),
            .I(N__17842));
    Span4Mux_s1_v I__2351 (
            .O(N__17849),
            .I(N__17837));
    Span4Mux_s1_h I__2350 (
            .O(N__17846),
            .I(N__17837));
    InMux I__2349 (
            .O(N__17845),
            .I(N__17832));
    InMux I__2348 (
            .O(N__17842),
            .I(N__17832));
    Odrv4 I__2347 (
            .O(N__17837),
            .I(\b2v_inst11.count_offZ0Z_0 ));
    LocalMux I__2346 (
            .O(N__17832),
            .I(\b2v_inst11.count_offZ0Z_0 ));
    InMux I__2345 (
            .O(N__17827),
            .I(N__17824));
    LocalMux I__2344 (
            .O(N__17824),
            .I(\b2v_inst11.count_off_0_0 ));
    InMux I__2343 (
            .O(N__17821),
            .I(N__17818));
    LocalMux I__2342 (
            .O(N__17818),
            .I(\b2v_inst11.count_off_0_10 ));
    CascadeMux I__2341 (
            .O(N__17815),
            .I(N__17812));
    InMux I__2340 (
            .O(N__17812),
            .I(N__17806));
    InMux I__2339 (
            .O(N__17811),
            .I(N__17806));
    LocalMux I__2338 (
            .O(N__17806),
            .I(N__17803));
    Odrv4 I__2337 (
            .O(N__17803),
            .I(\b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2 ));
    CascadeMux I__2336 (
            .O(N__17800),
            .I(N__17796));
    InMux I__2335 (
            .O(N__17799),
            .I(N__17793));
    InMux I__2334 (
            .O(N__17796),
            .I(N__17790));
    LocalMux I__2333 (
            .O(N__17793),
            .I(N__17787));
    LocalMux I__2332 (
            .O(N__17790),
            .I(N__17784));
    Span4Mux_s3_h I__2331 (
            .O(N__17787),
            .I(N__17781));
    Odrv4 I__2330 (
            .O(N__17784),
            .I(\b2v_inst11.count_offZ0Z_10 ));
    Odrv4 I__2329 (
            .O(N__17781),
            .I(\b2v_inst11.count_offZ0Z_10 ));
    InMux I__2328 (
            .O(N__17776),
            .I(N__17773));
    LocalMux I__2327 (
            .O(N__17773),
            .I(N__17769));
    InMux I__2326 (
            .O(N__17772),
            .I(N__17766));
    Odrv4 I__2325 (
            .O(N__17769),
            .I(\b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5 ));
    LocalMux I__2324 (
            .O(N__17766),
            .I(\b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5 ));
    InMux I__2323 (
            .O(N__17761),
            .I(N__17758));
    LocalMux I__2322 (
            .O(N__17758),
            .I(\b2v_inst11.dutycycle_RNIGKEF3Z0Z_12 ));
    CascadeMux I__2321 (
            .O(N__17755),
            .I(N__17752));
    InMux I__2320 (
            .O(N__17752),
            .I(N__17746));
    InMux I__2319 (
            .O(N__17751),
            .I(N__17746));
    LocalMux I__2318 (
            .O(N__17746),
            .I(\b2v_inst11.dutycycleZ1Z_12 ));
    CascadeMux I__2317 (
            .O(N__17743),
            .I(\b2v_inst11.dutycycle_RNIGKEF3Z0Z_12_cascade_ ));
    CascadeMux I__2316 (
            .O(N__17740),
            .I(\b2v_inst11.dutycycleZ0Z_10_cascade_ ));
    CascadeMux I__2315 (
            .O(N__17737),
            .I(\b2v_inst11.un1_dutycycle_53_56_a0_3_0_cascade_ ));
    InMux I__2314 (
            .O(N__17734),
            .I(N__17728));
    InMux I__2313 (
            .O(N__17733),
            .I(N__17728));
    LocalMux I__2312 (
            .O(N__17728),
            .I(\b2v_inst11.N_232_N ));
    CascadeMux I__2311 (
            .O(N__17725),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_325_N_cascade_ ));
    CascadeMux I__2310 (
            .O(N__17722),
            .I(\b2v_inst11.un1_func_state25_6_0_1_cascade_ ));
    InMux I__2309 (
            .O(N__17719),
            .I(N__17716));
    LocalMux I__2308 (
            .O(N__17716),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_323_N ));
    InMux I__2307 (
            .O(N__17713),
            .I(N__17710));
    LocalMux I__2306 (
            .O(N__17710),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_324_N ));
    CascadeMux I__2305 (
            .O(N__17707),
            .I(\b2v_inst11.N_289_cascade_ ));
    CascadeMux I__2304 (
            .O(N__17704),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_0_2_cascade_ ));
    CascadeMux I__2303 (
            .O(N__17701),
            .I(\b2v_inst11.N_302_cascade_ ));
    CascadeMux I__2302 (
            .O(N__17698),
            .I(\b2v_inst11.N_301_cascade_ ));
    CascadeMux I__2301 (
            .O(N__17695),
            .I(\b2v_inst11.dutycycle_RNIJU083Z0Z_8_cascade_ ));
    CascadeMux I__2300 (
            .O(N__17692),
            .I(\b2v_inst11.N_108_f0_cascade_ ));
    InMux I__2299 (
            .O(N__17689),
            .I(N__17686));
    LocalMux I__2298 (
            .O(N__17686),
            .I(\b2v_inst11.dutycycle_RNIHTFQZ0Z_8 ));
    CascadeMux I__2297 (
            .O(N__17683),
            .I(\b2v_inst11.dutycycle_RNI2NK31Z0Z_8_cascade_ ));
    InMux I__2296 (
            .O(N__17680),
            .I(N__17677));
    LocalMux I__2295 (
            .O(N__17677),
            .I(\b2v_inst11.dutycycle_e_1_8 ));
    InMux I__2294 (
            .O(N__17674),
            .I(N__17662));
    InMux I__2293 (
            .O(N__17673),
            .I(N__17662));
    InMux I__2292 (
            .O(N__17672),
            .I(N__17662));
    InMux I__2291 (
            .O(N__17671),
            .I(N__17662));
    LocalMux I__2290 (
            .O(N__17662),
            .I(\b2v_inst11.dutycycleZ1Z_8 ));
    InMux I__2289 (
            .O(N__17659),
            .I(N__17656));
    LocalMux I__2288 (
            .O(N__17656),
            .I(\b2v_inst11.N_108_f0 ));
    CascadeMux I__2287 (
            .O(N__17653),
            .I(\b2v_inst11.dutycycle_e_1_8_cascade_ ));
    CascadeMux I__2286 (
            .O(N__17650),
            .I(\b2v_inst11.dutycycleZ0Z_1_cascade_ ));
    InMux I__2285 (
            .O(N__17647),
            .I(N__17644));
    LocalMux I__2284 (
            .O(N__17644),
            .I(\b2v_inst11.dutycycle_RNIJU083_0Z0Z_8 ));
    IoInMux I__2283 (
            .O(N__17641),
            .I(N__17637));
    IoInMux I__2282 (
            .O(N__17640),
            .I(N__17634));
    LocalMux I__2281 (
            .O(N__17637),
            .I(N__17629));
    LocalMux I__2280 (
            .O(N__17634),
            .I(N__17629));
    IoSpan4Mux I__2279 (
            .O(N__17629),
            .I(N__17626));
    Span4Mux_s0_h I__2278 (
            .O(N__17626),
            .I(N__17622));
    IoInMux I__2277 (
            .O(N__17625),
            .I(N__17619));
    Sp12to4 I__2276 (
            .O(N__17622),
            .I(N__17614));
    LocalMux I__2275 (
            .O(N__17619),
            .I(N__17614));
    Odrv12 I__2274 (
            .O(N__17614),
            .I(delayed_vccin_vccinaux_ok_RNIM6F44_0));
    CascadeMux I__2273 (
            .O(N__17611),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_12_cascade_ ));
    CascadeMux I__2272 (
            .O(N__17608),
            .I(\b2v_inst11.dutycycle_RNI_10Z0Z_9_cascade_ ));
    InMux I__2271 (
            .O(N__17605),
            .I(N__17599));
    InMux I__2270 (
            .O(N__17604),
            .I(N__17599));
    LocalMux I__2269 (
            .O(N__17599),
            .I(\b2v_inst11.dutycycle_en_10 ));
    CascadeMux I__2268 (
            .O(N__17596),
            .I(N__17592));
    CascadeMux I__2267 (
            .O(N__17595),
            .I(N__17589));
    InMux I__2266 (
            .O(N__17592),
            .I(N__17584));
    InMux I__2265 (
            .O(N__17589),
            .I(N__17584));
    LocalMux I__2264 (
            .O(N__17584),
            .I(\b2v_inst11.dutycycleZ1Z_13 ));
    CascadeMux I__2263 (
            .O(N__17581),
            .I(\b2v_inst11.dutycycleZ0Z_9_cascade_ ));
    CascadeMux I__2262 (
            .O(N__17578),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_13_cascade_ ));
    CascadeMux I__2261 (
            .O(N__17575),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_10_cascade_ ));
    InMux I__2260 (
            .O(N__17572),
            .I(N__17569));
    LocalMux I__2259 (
            .O(N__17569),
            .I(N__17566));
    Span4Mux_v I__2258 (
            .O(N__17566),
            .I(N__17562));
    InMux I__2257 (
            .O(N__17565),
            .I(N__17559));
    Odrv4 I__2256 (
            .O(N__17562),
            .I(\b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5 ));
    LocalMux I__2255 (
            .O(N__17559),
            .I(\b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5 ));
    InMux I__2254 (
            .O(N__17554),
            .I(N__17551));
    LocalMux I__2253 (
            .O(N__17551),
            .I(N__17548));
    Span4Mux_s3_h I__2252 (
            .O(N__17548),
            .I(N__17545));
    Odrv4 I__2251 (
            .O(N__17545),
            .I(\b2v_inst11.count_clk_0_3 ));
    CEMux I__2250 (
            .O(N__17542),
            .I(N__17539));
    LocalMux I__2249 (
            .O(N__17539),
            .I(N__17534));
    CEMux I__2248 (
            .O(N__17538),
            .I(N__17531));
    CEMux I__2247 (
            .O(N__17537),
            .I(N__17528));
    Span4Mux_s2_h I__2246 (
            .O(N__17534),
            .I(N__17520));
    LocalMux I__2245 (
            .O(N__17531),
            .I(N__17515));
    LocalMux I__2244 (
            .O(N__17528),
            .I(N__17515));
    CEMux I__2243 (
            .O(N__17527),
            .I(N__17512));
    CEMux I__2242 (
            .O(N__17526),
            .I(N__17508));
    InMux I__2241 (
            .O(N__17525),
            .I(N__17501));
    InMux I__2240 (
            .O(N__17524),
            .I(N__17501));
    InMux I__2239 (
            .O(N__17523),
            .I(N__17501));
    Span4Mux_v I__2238 (
            .O(N__17520),
            .I(N__17496));
    Span4Mux_v I__2237 (
            .O(N__17515),
            .I(N__17489));
    LocalMux I__2236 (
            .O(N__17512),
            .I(N__17489));
    CEMux I__2235 (
            .O(N__17511),
            .I(N__17486));
    LocalMux I__2234 (
            .O(N__17508),
            .I(N__17477));
    LocalMux I__2233 (
            .O(N__17501),
            .I(N__17474));
    CascadeMux I__2232 (
            .O(N__17500),
            .I(N__17471));
    CascadeMux I__2231 (
            .O(N__17499),
            .I(N__17468));
    IoSpan4Mux I__2230 (
            .O(N__17496),
            .I(N__17463));
    InMux I__2229 (
            .O(N__17495),
            .I(N__17458));
    InMux I__2228 (
            .O(N__17494),
            .I(N__17458));
    Span4Mux_h I__2227 (
            .O(N__17489),
            .I(N__17455));
    LocalMux I__2226 (
            .O(N__17486),
            .I(N__17452));
    InMux I__2225 (
            .O(N__17485),
            .I(N__17447));
    InMux I__2224 (
            .O(N__17484),
            .I(N__17447));
    InMux I__2223 (
            .O(N__17483),
            .I(N__17438));
    InMux I__2222 (
            .O(N__17482),
            .I(N__17438));
    InMux I__2221 (
            .O(N__17481),
            .I(N__17438));
    InMux I__2220 (
            .O(N__17480),
            .I(N__17438));
    Span4Mux_h I__2219 (
            .O(N__17477),
            .I(N__17433));
    Span4Mux_s2_h I__2218 (
            .O(N__17474),
            .I(N__17433));
    InMux I__2217 (
            .O(N__17471),
            .I(N__17430));
    InMux I__2216 (
            .O(N__17468),
            .I(N__17423));
    InMux I__2215 (
            .O(N__17467),
            .I(N__17423));
    InMux I__2214 (
            .O(N__17466),
            .I(N__17423));
    Span4Mux_s3_v I__2213 (
            .O(N__17463),
            .I(N__17418));
    LocalMux I__2212 (
            .O(N__17458),
            .I(N__17418));
    Odrv4 I__2211 (
            .O(N__17455),
            .I(\b2v_inst11.count_clk_en ));
    Odrv12 I__2210 (
            .O(N__17452),
            .I(\b2v_inst11.count_clk_en ));
    LocalMux I__2209 (
            .O(N__17447),
            .I(\b2v_inst11.count_clk_en ));
    LocalMux I__2208 (
            .O(N__17438),
            .I(\b2v_inst11.count_clk_en ));
    Odrv4 I__2207 (
            .O(N__17433),
            .I(\b2v_inst11.count_clk_en ));
    LocalMux I__2206 (
            .O(N__17430),
            .I(\b2v_inst11.count_clk_en ));
    LocalMux I__2205 (
            .O(N__17423),
            .I(\b2v_inst11.count_clk_en ));
    Odrv4 I__2204 (
            .O(N__17418),
            .I(\b2v_inst11.count_clk_en ));
    CascadeMux I__2203 (
            .O(N__17401),
            .I(N__17398));
    InMux I__2202 (
            .O(N__17398),
            .I(N__17395));
    LocalMux I__2201 (
            .O(N__17395),
            .I(\b2v_inst11.N_150_N ));
    CascadeMux I__2200 (
            .O(N__17392),
            .I(\b2v_inst11.N_152_N_cascade_ ));
    CascadeMux I__2199 (
            .O(N__17389),
            .I(\b2v_inst11.dutycycleZ0Z_12_cascade_ ));
    CascadeMux I__2198 (
            .O(N__17386),
            .I(\b2v_inst11.N_155_N_cascade_ ));
    InMux I__2197 (
            .O(N__17383),
            .I(N__17380));
    LocalMux I__2196 (
            .O(N__17380),
            .I(\b2v_inst11.dutycycle_en_12 ));
    CascadeMux I__2195 (
            .O(N__17377),
            .I(\b2v_inst11.dutycycle_en_12_cascade_ ));
    InMux I__2194 (
            .O(N__17374),
            .I(N__17370));
    InMux I__2193 (
            .O(N__17373),
            .I(N__17367));
    LocalMux I__2192 (
            .O(N__17370),
            .I(\b2v_inst11.dutycycleZ0Z_15 ));
    LocalMux I__2191 (
            .O(N__17367),
            .I(\b2v_inst11.dutycycleZ0Z_15 ));
    IoInMux I__2190 (
            .O(N__17362),
            .I(N__17359));
    LocalMux I__2189 (
            .O(N__17359),
            .I(N__17356));
    Span4Mux_s3_h I__2188 (
            .O(N__17356),
            .I(N__17353));
    Odrv4 I__2187 (
            .O(N__17353),
            .I(\b2v_inst200.count_enZ0 ));
    CascadeMux I__2186 (
            .O(N__17350),
            .I(N__17347));
    InMux I__2185 (
            .O(N__17347),
            .I(N__17344));
    LocalMux I__2184 (
            .O(N__17344),
            .I(\b2v_inst11.un1_dutycycle_53_i_29 ));
    CascadeMux I__2183 (
            .O(N__17341),
            .I(N__17338));
    InMux I__2182 (
            .O(N__17338),
            .I(N__17335));
    LocalMux I__2181 (
            .O(N__17335),
            .I(\b2v_inst11.mult1_un40_sum_i_l_ofx_4 ));
    CascadeMux I__2180 (
            .O(N__17332),
            .I(N__17329));
    InMux I__2179 (
            .O(N__17329),
            .I(N__17326));
    LocalMux I__2178 (
            .O(N__17326),
            .I(\b2v_inst11.mult1_un47_sum_s_4_sf ));
    CascadeMux I__2177 (
            .O(N__17323),
            .I(\b2v_inst11.mult1_un40_sum_i_5_cascade_ ));
    InMux I__2176 (
            .O(N__17320),
            .I(N__17316));
    InMux I__2175 (
            .O(N__17319),
            .I(N__17313));
    LocalMux I__2174 (
            .O(N__17316),
            .I(N__17310));
    LocalMux I__2173 (
            .O(N__17313),
            .I(N__17307));
    Span4Mux_s3_h I__2172 (
            .O(N__17310),
            .I(N__17304));
    Span4Mux_s3_h I__2171 (
            .O(N__17307),
            .I(N__17301));
    Odrv4 I__2170 (
            .O(N__17304),
            .I(\b2v_inst16.countZ0Z_10 ));
    Odrv4 I__2169 (
            .O(N__17301),
            .I(\b2v_inst16.countZ0Z_10 ));
    InMux I__2168 (
            .O(N__17296),
            .I(N__17290));
    InMux I__2167 (
            .O(N__17295),
            .I(N__17290));
    LocalMux I__2166 (
            .O(N__17290),
            .I(N__17287));
    Span4Mux_h I__2165 (
            .O(N__17287),
            .I(N__17284));
    Odrv4 I__2164 (
            .O(N__17284),
            .I(\b2v_inst16.count_rst ));
    InMux I__2163 (
            .O(N__17281),
            .I(N__17278));
    LocalMux I__2162 (
            .O(N__17278),
            .I(\b2v_inst16.count_4_10 ));
    InMux I__2161 (
            .O(N__17275),
            .I(\b2v_inst11.mult1_un47_sum_cry_2 ));
    InMux I__2160 (
            .O(N__17272),
            .I(\b2v_inst11.mult1_un47_sum_cry_3 ));
    InMux I__2159 (
            .O(N__17269),
            .I(\b2v_inst11.mult1_un47_sum_cry_4 ));
    InMux I__2158 (
            .O(N__17266),
            .I(\b2v_inst11.mult1_un47_sum_cry_5 ));
    InMux I__2157 (
            .O(N__17263),
            .I(N__17260));
    LocalMux I__2156 (
            .O(N__17260),
            .I(\b2v_inst11.mult1_un75_sum_cry_3_s ));
    InMux I__2155 (
            .O(N__17257),
            .I(\b2v_inst11.mult1_un75_sum_cry_2 ));
    CascadeMux I__2154 (
            .O(N__17254),
            .I(N__17251));
    InMux I__2153 (
            .O(N__17251),
            .I(N__17248));
    LocalMux I__2152 (
            .O(N__17248),
            .I(\b2v_inst11.mult1_un75_sum_cry_4_s ));
    InMux I__2151 (
            .O(N__17245),
            .I(\b2v_inst11.mult1_un75_sum_cry_3 ));
    InMux I__2150 (
            .O(N__17242),
            .I(N__17239));
    LocalMux I__2149 (
            .O(N__17239),
            .I(\b2v_inst11.mult1_un75_sum_cry_5_s ));
    InMux I__2148 (
            .O(N__17236),
            .I(\b2v_inst11.mult1_un75_sum_cry_4 ));
    CascadeMux I__2147 (
            .O(N__17233),
            .I(N__17230));
    InMux I__2146 (
            .O(N__17230),
            .I(N__17227));
    LocalMux I__2145 (
            .O(N__17227),
            .I(\b2v_inst11.mult1_un75_sum_cry_6_s ));
    InMux I__2144 (
            .O(N__17224),
            .I(\b2v_inst11.mult1_un75_sum_cry_5 ));
    InMux I__2143 (
            .O(N__17221),
            .I(N__17218));
    LocalMux I__2142 (
            .O(N__17218),
            .I(\b2v_inst11.mult1_un82_sum_axb_8 ));
    InMux I__2141 (
            .O(N__17215),
            .I(\b2v_inst11.mult1_un75_sum_cry_6 ));
    InMux I__2140 (
            .O(N__17212),
            .I(\b2v_inst11.mult1_un75_sum_cry_7 ));
    CascadeMux I__2139 (
            .O(N__17209),
            .I(\b2v_inst11.mult1_un75_sum_s_8_cascade_ ));
    CascadeMux I__2138 (
            .O(N__17206),
            .I(N__17202));
    InMux I__2137 (
            .O(N__17205),
            .I(N__17194));
    InMux I__2136 (
            .O(N__17202),
            .I(N__17194));
    InMux I__2135 (
            .O(N__17201),
            .I(N__17194));
    LocalMux I__2134 (
            .O(N__17194),
            .I(\b2v_inst11.mult1_un75_sum_i_0_8 ));
    InMux I__2133 (
            .O(N__17191),
            .I(\b2v_inst11.mult1_un89_sum_cry_7 ));
    CascadeMux I__2132 (
            .O(N__17188),
            .I(N__17184));
    InMux I__2131 (
            .O(N__17187),
            .I(N__17176));
    InMux I__2130 (
            .O(N__17184),
            .I(N__17176));
    InMux I__2129 (
            .O(N__17183),
            .I(N__17176));
    LocalMux I__2128 (
            .O(N__17176),
            .I(\b2v_inst11.mult1_un82_sum_i_0_8 ));
    InMux I__2127 (
            .O(N__17173),
            .I(N__17170));
    LocalMux I__2126 (
            .O(N__17170),
            .I(\b2v_inst11.mult1_un82_sum_cry_3_s ));
    InMux I__2125 (
            .O(N__17167),
            .I(\b2v_inst11.mult1_un82_sum_cry_2 ));
    CascadeMux I__2124 (
            .O(N__17164),
            .I(N__17161));
    InMux I__2123 (
            .O(N__17161),
            .I(N__17158));
    LocalMux I__2122 (
            .O(N__17158),
            .I(\b2v_inst11.mult1_un82_sum_cry_4_s ));
    InMux I__2121 (
            .O(N__17155),
            .I(\b2v_inst11.mult1_un82_sum_cry_3 ));
    InMux I__2120 (
            .O(N__17152),
            .I(N__17149));
    LocalMux I__2119 (
            .O(N__17149),
            .I(\b2v_inst11.mult1_un82_sum_cry_5_s ));
    InMux I__2118 (
            .O(N__17146),
            .I(\b2v_inst11.mult1_un82_sum_cry_4 ));
    CascadeMux I__2117 (
            .O(N__17143),
            .I(N__17140));
    InMux I__2116 (
            .O(N__17140),
            .I(N__17137));
    LocalMux I__2115 (
            .O(N__17137),
            .I(\b2v_inst11.mult1_un82_sum_cry_6_s ));
    InMux I__2114 (
            .O(N__17134),
            .I(\b2v_inst11.mult1_un82_sum_cry_5 ));
    InMux I__2113 (
            .O(N__17131),
            .I(N__17128));
    LocalMux I__2112 (
            .O(N__17128),
            .I(\b2v_inst11.mult1_un89_sum_axb_8 ));
    InMux I__2111 (
            .O(N__17125),
            .I(\b2v_inst11.mult1_un82_sum_cry_6 ));
    InMux I__2110 (
            .O(N__17122),
            .I(\b2v_inst11.mult1_un82_sum_cry_7 ));
    InMux I__2109 (
            .O(N__17119),
            .I(\b2v_inst11.mult1_un96_sum_cry_6 ));
    InMux I__2108 (
            .O(N__17116),
            .I(\b2v_inst11.mult1_un96_sum_cry_7 ));
    CascadeMux I__2107 (
            .O(N__17113),
            .I(\b2v_inst11.mult1_un96_sum_s_8_cascade_ ));
    InMux I__2106 (
            .O(N__17110),
            .I(N__17107));
    LocalMux I__2105 (
            .O(N__17107),
            .I(\b2v_inst11.mult1_un89_sum_cry_3_s ));
    InMux I__2104 (
            .O(N__17104),
            .I(\b2v_inst11.mult1_un89_sum_cry_2 ));
    CascadeMux I__2103 (
            .O(N__17101),
            .I(N__17098));
    InMux I__2102 (
            .O(N__17098),
            .I(N__17095));
    LocalMux I__2101 (
            .O(N__17095),
            .I(\b2v_inst11.mult1_un89_sum_cry_4_s ));
    InMux I__2100 (
            .O(N__17092),
            .I(\b2v_inst11.mult1_un89_sum_cry_3 ));
    InMux I__2099 (
            .O(N__17089),
            .I(N__17086));
    LocalMux I__2098 (
            .O(N__17086),
            .I(\b2v_inst11.mult1_un89_sum_cry_5_s ));
    InMux I__2097 (
            .O(N__17083),
            .I(\b2v_inst11.mult1_un89_sum_cry_4 ));
    CascadeMux I__2096 (
            .O(N__17080),
            .I(N__17077));
    InMux I__2095 (
            .O(N__17077),
            .I(N__17074));
    LocalMux I__2094 (
            .O(N__17074),
            .I(\b2v_inst11.mult1_un89_sum_cry_6_s ));
    InMux I__2093 (
            .O(N__17071),
            .I(\b2v_inst11.mult1_un89_sum_cry_5 ));
    InMux I__2092 (
            .O(N__17068),
            .I(N__17065));
    LocalMux I__2091 (
            .O(N__17065),
            .I(\b2v_inst11.mult1_un96_sum_axb_8 ));
    InMux I__2090 (
            .O(N__17062),
            .I(\b2v_inst11.mult1_un89_sum_cry_6 ));
    InMux I__2089 (
            .O(N__17059),
            .I(N__17056));
    LocalMux I__2088 (
            .O(N__17056),
            .I(\b2v_inst11.count_off_0_8 ));
    CascadeMux I__2087 (
            .O(N__17053),
            .I(N__17050));
    InMux I__2086 (
            .O(N__17050),
            .I(N__17044));
    InMux I__2085 (
            .O(N__17049),
            .I(N__17044));
    LocalMux I__2084 (
            .O(N__17044),
            .I(N__17041));
    Odrv4 I__2083 (
            .O(N__17041),
            .I(\b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2 ));
    CascadeMux I__2082 (
            .O(N__17038),
            .I(N__17035));
    InMux I__2081 (
            .O(N__17035),
            .I(N__17032));
    LocalMux I__2080 (
            .O(N__17032),
            .I(N__17029));
    Odrv4 I__2079 (
            .O(N__17029),
            .I(\b2v_inst11.count_offZ0Z_8 ));
    CascadeMux I__2078 (
            .O(N__17026),
            .I(\b2v_inst11.count_offZ0Z_8_cascade_ ));
    InMux I__2077 (
            .O(N__17023),
            .I(N__17020));
    LocalMux I__2076 (
            .O(N__17020),
            .I(N__17017));
    Span4Mux_v I__2075 (
            .O(N__17017),
            .I(N__17014));
    Odrv4 I__2074 (
            .O(N__17014),
            .I(\b2v_inst11.un34_clk_100khz_3 ));
    InMux I__2073 (
            .O(N__17011),
            .I(N__17005));
    InMux I__2072 (
            .O(N__17010),
            .I(N__17005));
    LocalMux I__2071 (
            .O(N__17005),
            .I(\b2v_inst11.count_offZ0Z_7 ));
    InMux I__2070 (
            .O(N__17002),
            .I(N__16998));
    InMux I__2069 (
            .O(N__17001),
            .I(N__16995));
    LocalMux I__2068 (
            .O(N__16998),
            .I(\b2v_inst11.count_off_1_7 ));
    LocalMux I__2067 (
            .O(N__16995),
            .I(\b2v_inst11.count_off_1_7 ));
    CascadeMux I__2066 (
            .O(N__16990),
            .I(N__16987));
    InMux I__2065 (
            .O(N__16987),
            .I(N__16984));
    LocalMux I__2064 (
            .O(N__16984),
            .I(N__16981));
    Odrv4 I__2063 (
            .O(N__16981),
            .I(\b2v_inst11.un3_count_off_1_axb_7 ));
    InMux I__2062 (
            .O(N__16978),
            .I(\b2v_inst11.mult1_un96_sum_cry_2 ));
    InMux I__2061 (
            .O(N__16975),
            .I(\b2v_inst11.mult1_un96_sum_cry_3 ));
    InMux I__2060 (
            .O(N__16972),
            .I(\b2v_inst11.mult1_un96_sum_cry_4 ));
    InMux I__2059 (
            .O(N__16969),
            .I(\b2v_inst11.mult1_un96_sum_cry_5 ));
    CascadeMux I__2058 (
            .O(N__16966),
            .I(\b2v_inst11.count_off_1_9_cascade_ ));
    CascadeMux I__2057 (
            .O(N__16963),
            .I(N__16959));
    InMux I__2056 (
            .O(N__16962),
            .I(N__16956));
    InMux I__2055 (
            .O(N__16959),
            .I(N__16953));
    LocalMux I__2054 (
            .O(N__16956),
            .I(\b2v_inst11.count_offZ0Z_9 ));
    LocalMux I__2053 (
            .O(N__16953),
            .I(\b2v_inst11.count_offZ0Z_9 ));
    CascadeMux I__2052 (
            .O(N__16948),
            .I(N__16945));
    InMux I__2051 (
            .O(N__16945),
            .I(N__16942));
    LocalMux I__2050 (
            .O(N__16942),
            .I(\b2v_inst11.un3_count_off_1_axb_9 ));
    InMux I__2049 (
            .O(N__16939),
            .I(N__16933));
    InMux I__2048 (
            .O(N__16938),
            .I(N__16933));
    LocalMux I__2047 (
            .O(N__16933),
            .I(\b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92 ));
    CascadeMux I__2046 (
            .O(N__16930),
            .I(N__16927));
    InMux I__2045 (
            .O(N__16927),
            .I(N__16924));
    LocalMux I__2044 (
            .O(N__16924),
            .I(N__16920));
    InMux I__2043 (
            .O(N__16923),
            .I(N__16917));
    Span4Mux_s1_h I__2042 (
            .O(N__16920),
            .I(N__16914));
    LocalMux I__2041 (
            .O(N__16917),
            .I(N__16911));
    Odrv4 I__2040 (
            .O(N__16914),
            .I(\b2v_inst11.count_off_1_6 ));
    Odrv4 I__2039 (
            .O(N__16911),
            .I(\b2v_inst11.count_off_1_6 ));
    InMux I__2038 (
            .O(N__16906),
            .I(N__16902));
    InMux I__2037 (
            .O(N__16905),
            .I(N__16899));
    LocalMux I__2036 (
            .O(N__16902),
            .I(\b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2 ));
    LocalMux I__2035 (
            .O(N__16899),
            .I(\b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2 ));
    InMux I__2034 (
            .O(N__16894),
            .I(N__16891));
    LocalMux I__2033 (
            .O(N__16891),
            .I(\b2v_inst11.count_off_0_15 ));
    InMux I__2032 (
            .O(N__16888),
            .I(N__16884));
    InMux I__2031 (
            .O(N__16887),
            .I(N__16881));
    LocalMux I__2030 (
            .O(N__16884),
            .I(\b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5 ));
    LocalMux I__2029 (
            .O(N__16881),
            .I(\b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5 ));
    InMux I__2028 (
            .O(N__16876),
            .I(N__16873));
    LocalMux I__2027 (
            .O(N__16873),
            .I(\b2v_inst11.count_offZ0Z_15 ));
    CascadeMux I__2026 (
            .O(N__16870),
            .I(N__16866));
    InMux I__2025 (
            .O(N__16869),
            .I(N__16863));
    InMux I__2024 (
            .O(N__16866),
            .I(N__16860));
    LocalMux I__2023 (
            .O(N__16863),
            .I(\b2v_inst11.count_offZ0Z_13 ));
    LocalMux I__2022 (
            .O(N__16860),
            .I(\b2v_inst11.count_offZ0Z_13 ));
    InMux I__2021 (
            .O(N__16855),
            .I(N__16851));
    CascadeMux I__2020 (
            .O(N__16854),
            .I(N__16848));
    LocalMux I__2019 (
            .O(N__16851),
            .I(N__16845));
    InMux I__2018 (
            .O(N__16848),
            .I(N__16842));
    Odrv4 I__2017 (
            .O(N__16845),
            .I(\b2v_inst11.count_offZ0Z_14 ));
    LocalMux I__2016 (
            .O(N__16842),
            .I(\b2v_inst11.count_offZ0Z_14 ));
    CascadeMux I__2015 (
            .O(N__16837),
            .I(\b2v_inst11.count_offZ0Z_15_cascade_ ));
    InMux I__2014 (
            .O(N__16834),
            .I(N__16831));
    LocalMux I__2013 (
            .O(N__16831),
            .I(N__16828));
    Odrv4 I__2012 (
            .O(N__16828),
            .I(\b2v_inst11.un34_clk_100khz_11 ));
    InMux I__2011 (
            .O(N__16825),
            .I(N__16819));
    InMux I__2010 (
            .O(N__16824),
            .I(N__16819));
    LocalMux I__2009 (
            .O(N__16819),
            .I(\b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5 ));
    InMux I__2008 (
            .O(N__16816),
            .I(N__16813));
    LocalMux I__2007 (
            .O(N__16813),
            .I(\b2v_inst11.un34_clk_100khz_12 ));
    CascadeMux I__2006 (
            .O(N__16810),
            .I(\b2v_inst11.un34_clk_100khz_4_cascade_ ));
    CascadeMux I__2005 (
            .O(N__16807),
            .I(N__16804));
    InMux I__2004 (
            .O(N__16804),
            .I(N__16801));
    LocalMux I__2003 (
            .O(N__16801),
            .I(\b2v_inst11.count_off_0_12 ));
    CascadeMux I__2002 (
            .O(N__16798),
            .I(N__16795));
    InMux I__2001 (
            .O(N__16795),
            .I(N__16789));
    InMux I__2000 (
            .O(N__16794),
            .I(N__16789));
    LocalMux I__1999 (
            .O(N__16789),
            .I(\b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5 ));
    CascadeMux I__1998 (
            .O(N__16786),
            .I(N__16783));
    InMux I__1997 (
            .O(N__16783),
            .I(N__16780));
    LocalMux I__1996 (
            .O(N__16780),
            .I(\b2v_inst11.count_offZ0Z_12 ));
    InMux I__1995 (
            .O(N__16777),
            .I(N__16774));
    LocalMux I__1994 (
            .O(N__16774),
            .I(\b2v_inst11.count_off_1_11 ));
    InMux I__1993 (
            .O(N__16771),
            .I(N__16765));
    InMux I__1992 (
            .O(N__16770),
            .I(N__16765));
    LocalMux I__1991 (
            .O(N__16765),
            .I(\b2v_inst11.count_offZ0Z_11 ));
    CascadeMux I__1990 (
            .O(N__16762),
            .I(\b2v_inst11.count_offZ0Z_12_cascade_ ));
    InMux I__1989 (
            .O(N__16759),
            .I(N__16756));
    LocalMux I__1988 (
            .O(N__16756),
            .I(\b2v_inst11.un34_clk_100khz_5 ));
    InMux I__1987 (
            .O(N__16753),
            .I(N__16749));
    InMux I__1986 (
            .O(N__16752),
            .I(N__16746));
    LocalMux I__1985 (
            .O(N__16749),
            .I(N__16743));
    LocalMux I__1984 (
            .O(N__16746),
            .I(N__16740));
    Odrv4 I__1983 (
            .O(N__16743),
            .I(\b2v_inst11.count_offZ0Z_6 ));
    Odrv4 I__1982 (
            .O(N__16740),
            .I(\b2v_inst11.count_offZ0Z_6 ));
    CascadeMux I__1981 (
            .O(N__16735),
            .I(N__16732));
    InMux I__1980 (
            .O(N__16732),
            .I(N__16726));
    InMux I__1979 (
            .O(N__16731),
            .I(N__16726));
    LocalMux I__1978 (
            .O(N__16726),
            .I(\b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2 ));
    InMux I__1977 (
            .O(N__16723),
            .I(N__16720));
    LocalMux I__1976 (
            .O(N__16720),
            .I(\b2v_inst11.count_off_1_9 ));
    CascadeMux I__1975 (
            .O(N__16717),
            .I(N__16714));
    InMux I__1974 (
            .O(N__16714),
            .I(N__16709));
    InMux I__1973 (
            .O(N__16713),
            .I(N__16704));
    InMux I__1972 (
            .O(N__16712),
            .I(N__16704));
    LocalMux I__1971 (
            .O(N__16709),
            .I(N__16701));
    LocalMux I__1970 (
            .O(N__16704),
            .I(\b2v_inst11.count_clkZ0Z_9 ));
    Odrv4 I__1969 (
            .O(N__16701),
            .I(\b2v_inst11.count_clkZ0Z_9 ));
    CascadeMux I__1968 (
            .O(N__16696),
            .I(N__16693));
    InMux I__1967 (
            .O(N__16693),
            .I(N__16687));
    InMux I__1966 (
            .O(N__16692),
            .I(N__16680));
    InMux I__1965 (
            .O(N__16691),
            .I(N__16680));
    InMux I__1964 (
            .O(N__16690),
            .I(N__16680));
    LocalMux I__1963 (
            .O(N__16687),
            .I(N__16677));
    LocalMux I__1962 (
            .O(N__16680),
            .I(\b2v_inst11.count_clkZ0Z_1 ));
    Odrv4 I__1961 (
            .O(N__16677),
            .I(\b2v_inst11.count_clkZ0Z_1 ));
    CascadeMux I__1960 (
            .O(N__16672),
            .I(N__16669));
    InMux I__1959 (
            .O(N__16669),
            .I(N__16666));
    LocalMux I__1958 (
            .O(N__16666),
            .I(\b2v_inst11.count_clk_RNIZ0Z_5 ));
    InMux I__1957 (
            .O(N__16663),
            .I(N__16657));
    InMux I__1956 (
            .O(N__16662),
            .I(N__16657));
    LocalMux I__1955 (
            .O(N__16657),
            .I(N__16654));
    Odrv4 I__1954 (
            .O(N__16654),
            .I(\b2v_inst11.N_172 ));
    CascadeMux I__1953 (
            .O(N__16651),
            .I(N__16648));
    InMux I__1952 (
            .O(N__16648),
            .I(N__16645));
    LocalMux I__1951 (
            .O(N__16645),
            .I(N__16642));
    Span4Mux_v I__1950 (
            .O(N__16642),
            .I(N__16638));
    InMux I__1949 (
            .O(N__16641),
            .I(N__16635));
    Odrv4 I__1948 (
            .O(N__16638),
            .I(\b2v_inst11.N_421 ));
    LocalMux I__1947 (
            .O(N__16635),
            .I(\b2v_inst11.N_421 ));
    CascadeMux I__1946 (
            .O(N__16630),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ));
    InMux I__1945 (
            .O(N__16627),
            .I(N__16624));
    LocalMux I__1944 (
            .O(N__16624),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_i_1 ));
    CascadeMux I__1943 (
            .O(N__16621),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_0_cascade_ ));
    InMux I__1942 (
            .O(N__16618),
            .I(N__16614));
    CascadeMux I__1941 (
            .O(N__16617),
            .I(N__16607));
    LocalMux I__1940 (
            .O(N__16614),
            .I(N__16596));
    InMux I__1939 (
            .O(N__16613),
            .I(N__16582));
    InMux I__1938 (
            .O(N__16612),
            .I(N__16582));
    InMux I__1937 (
            .O(N__16611),
            .I(N__16582));
    InMux I__1936 (
            .O(N__16610),
            .I(N__16582));
    InMux I__1935 (
            .O(N__16607),
            .I(N__16582));
    InMux I__1934 (
            .O(N__16606),
            .I(N__16573));
    InMux I__1933 (
            .O(N__16605),
            .I(N__16573));
    InMux I__1932 (
            .O(N__16604),
            .I(N__16573));
    InMux I__1931 (
            .O(N__16603),
            .I(N__16573));
    InMux I__1930 (
            .O(N__16602),
            .I(N__16566));
    InMux I__1929 (
            .O(N__16601),
            .I(N__16566));
    InMux I__1928 (
            .O(N__16600),
            .I(N__16566));
    CascadeMux I__1927 (
            .O(N__16599),
            .I(N__16561));
    Span4Mux_v I__1926 (
            .O(N__16596),
            .I(N__16558));
    InMux I__1925 (
            .O(N__16595),
            .I(N__16551));
    InMux I__1924 (
            .O(N__16594),
            .I(N__16551));
    InMux I__1923 (
            .O(N__16593),
            .I(N__16551));
    LocalMux I__1922 (
            .O(N__16582),
            .I(N__16544));
    LocalMux I__1921 (
            .O(N__16573),
            .I(N__16544));
    LocalMux I__1920 (
            .O(N__16566),
            .I(N__16544));
    InMux I__1919 (
            .O(N__16565),
            .I(N__16535));
    InMux I__1918 (
            .O(N__16564),
            .I(N__16535));
    InMux I__1917 (
            .O(N__16561),
            .I(N__16535));
    Span4Mux_s1_h I__1916 (
            .O(N__16558),
            .I(N__16530));
    LocalMux I__1915 (
            .O(N__16551),
            .I(N__16530));
    Span4Mux_s2_h I__1914 (
            .O(N__16544),
            .I(N__16527));
    InMux I__1913 (
            .O(N__16543),
            .I(N__16522));
    InMux I__1912 (
            .O(N__16542),
            .I(N__16522));
    LocalMux I__1911 (
            .O(N__16535),
            .I(\b2v_inst11.func_state_RNICC5V2_0_1 ));
    Odrv4 I__1910 (
            .O(N__16530),
            .I(\b2v_inst11.func_state_RNICC5V2_0_1 ));
    Odrv4 I__1909 (
            .O(N__16527),
            .I(\b2v_inst11.func_state_RNICC5V2_0_1 ));
    LocalMux I__1908 (
            .O(N__16522),
            .I(\b2v_inst11.func_state_RNICC5V2_0_1 ));
    CascadeMux I__1907 (
            .O(N__16513),
            .I(\b2v_inst11.count_off_1_11_cascade_ ));
    CascadeMux I__1906 (
            .O(N__16510),
            .I(N__16507));
    InMux I__1905 (
            .O(N__16507),
            .I(N__16504));
    LocalMux I__1904 (
            .O(N__16504),
            .I(\b2v_inst11.un3_count_off_1_axb_11 ));
    CascadeMux I__1903 (
            .O(N__16501),
            .I(\b2v_inst11.count_clk_RNIZ0Z_3_cascade_ ));
    CascadeMux I__1902 (
            .O(N__16498),
            .I(N__16495));
    InMux I__1901 (
            .O(N__16495),
            .I(N__16492));
    LocalMux I__1900 (
            .O(N__16492),
            .I(\b2v_inst11.count_clk_en_0 ));
    CascadeMux I__1899 (
            .O(N__16489),
            .I(N__16485));
    InMux I__1898 (
            .O(N__16488),
            .I(N__16482));
    InMux I__1897 (
            .O(N__16485),
            .I(N__16479));
    LocalMux I__1896 (
            .O(N__16482),
            .I(N__16474));
    LocalMux I__1895 (
            .O(N__16479),
            .I(N__16474));
    Odrv4 I__1894 (
            .O(N__16474),
            .I(\b2v_inst11.count_clkZ0Z_12 ));
    CascadeMux I__1893 (
            .O(N__16471),
            .I(N__16468));
    InMux I__1892 (
            .O(N__16468),
            .I(N__16462));
    InMux I__1891 (
            .O(N__16467),
            .I(N__16462));
    LocalMux I__1890 (
            .O(N__16462),
            .I(N__16459));
    Odrv4 I__1889 (
            .O(N__16459),
            .I(\b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BAZ0 ));
    InMux I__1888 (
            .O(N__16456),
            .I(N__16453));
    LocalMux I__1887 (
            .O(N__16453),
            .I(\b2v_inst11.count_clk_0_12 ));
    InMux I__1886 (
            .O(N__16450),
            .I(N__16447));
    LocalMux I__1885 (
            .O(N__16447),
            .I(N__16444));
    Odrv4 I__1884 (
            .O(N__16444),
            .I(\b2v_inst11.count_clk_RNI_0Z0Z_0 ));
    InMux I__1883 (
            .O(N__16441),
            .I(N__16432));
    InMux I__1882 (
            .O(N__16440),
            .I(N__16432));
    InMux I__1881 (
            .O(N__16439),
            .I(N__16432));
    LocalMux I__1880 (
            .O(N__16432),
            .I(N__16427));
    InMux I__1879 (
            .O(N__16431),
            .I(N__16424));
    InMux I__1878 (
            .O(N__16430),
            .I(N__16421));
    Odrv12 I__1877 (
            .O(N__16427),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    LocalMux I__1876 (
            .O(N__16424),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    LocalMux I__1875 (
            .O(N__16421),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    InMux I__1874 (
            .O(N__16414),
            .I(N__16411));
    LocalMux I__1873 (
            .O(N__16411),
            .I(\b2v_inst11.count_clk_0_1 ));
    CascadeMux I__1872 (
            .O(N__16408),
            .I(\b2v_inst11.count_clk_RNIZ0Z_0_cascade_ ));
    CascadeMux I__1871 (
            .O(N__16405),
            .I(\b2v_inst11.count_clkZ0Z_1_cascade_ ));
    CascadeMux I__1870 (
            .O(N__16402),
            .I(N__16399));
    InMux I__1869 (
            .O(N__16399),
            .I(N__16394));
    InMux I__1868 (
            .O(N__16398),
            .I(N__16391));
    InMux I__1867 (
            .O(N__16397),
            .I(N__16388));
    LocalMux I__1866 (
            .O(N__16394),
            .I(N__16385));
    LocalMux I__1865 (
            .O(N__16391),
            .I(\b2v_inst11.count_clkZ0Z_5 ));
    LocalMux I__1864 (
            .O(N__16388),
            .I(\b2v_inst11.count_clkZ0Z_5 ));
    Odrv4 I__1863 (
            .O(N__16385),
            .I(\b2v_inst11.count_clkZ0Z_5 ));
    InMux I__1862 (
            .O(N__16378),
            .I(N__16372));
    InMux I__1861 (
            .O(N__16377),
            .I(N__16372));
    LocalMux I__1860 (
            .O(N__16372),
            .I(\b2v_inst11.N_187 ));
    CascadeMux I__1859 (
            .O(N__16369),
            .I(\b2v_inst11.count_clk_en_cascade_ ));
    InMux I__1858 (
            .O(N__16366),
            .I(N__16360));
    InMux I__1857 (
            .O(N__16365),
            .I(N__16360));
    LocalMux I__1856 (
            .O(N__16360),
            .I(\b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5 ));
    InMux I__1855 (
            .O(N__16357),
            .I(N__16354));
    LocalMux I__1854 (
            .O(N__16354),
            .I(\b2v_inst11.count_clk_0_2 ));
    CascadeMux I__1853 (
            .O(N__16351),
            .I(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_ ));
    InMux I__1852 (
            .O(N__16348),
            .I(N__16345));
    LocalMux I__1851 (
            .O(N__16345),
            .I(\b2v_inst11.N_373 ));
    CascadeMux I__1850 (
            .O(N__16342),
            .I(\b2v_inst11.N_373_cascade_ ));
    CascadeMux I__1849 (
            .O(N__16339),
            .I(N__16336));
    InMux I__1848 (
            .O(N__16336),
            .I(N__16331));
    InMux I__1847 (
            .O(N__16335),
            .I(N__16326));
    InMux I__1846 (
            .O(N__16334),
            .I(N__16326));
    LocalMux I__1845 (
            .O(N__16331),
            .I(N__16323));
    LocalMux I__1844 (
            .O(N__16326),
            .I(\b2v_inst11.count_clkZ0Z_8 ));
    Odrv4 I__1843 (
            .O(N__16323),
            .I(\b2v_inst11.count_clkZ0Z_8 ));
    CascadeMux I__1842 (
            .O(N__16318),
            .I(N__16315));
    InMux I__1841 (
            .O(N__16315),
            .I(N__16310));
    InMux I__1840 (
            .O(N__16314),
            .I(N__16305));
    InMux I__1839 (
            .O(N__16313),
            .I(N__16305));
    LocalMux I__1838 (
            .O(N__16310),
            .I(N__16302));
    LocalMux I__1837 (
            .O(N__16305),
            .I(\b2v_inst11.count_clkZ0Z_6 ));
    Odrv4 I__1836 (
            .O(N__16302),
            .I(\b2v_inst11.count_clkZ0Z_6 ));
    CascadeMux I__1835 (
            .O(N__16297),
            .I(N__16293));
    CascadeMux I__1834 (
            .O(N__16296),
            .I(N__16290));
    InMux I__1833 (
            .O(N__16293),
            .I(N__16286));
    InMux I__1832 (
            .O(N__16290),
            .I(N__16283));
    InMux I__1831 (
            .O(N__16289),
            .I(N__16280));
    LocalMux I__1830 (
            .O(N__16286),
            .I(N__16277));
    LocalMux I__1829 (
            .O(N__16283),
            .I(\b2v_inst11.count_clkZ0Z_4 ));
    LocalMux I__1828 (
            .O(N__16280),
            .I(\b2v_inst11.count_clkZ0Z_4 ));
    Odrv4 I__1827 (
            .O(N__16277),
            .I(\b2v_inst11.count_clkZ0Z_4 ));
    InMux I__1826 (
            .O(N__16270),
            .I(N__16265));
    InMux I__1825 (
            .O(N__16269),
            .I(N__16260));
    InMux I__1824 (
            .O(N__16268),
            .I(N__16260));
    LocalMux I__1823 (
            .O(N__16265),
            .I(\b2v_inst11.count_clkZ0Z_2 ));
    LocalMux I__1822 (
            .O(N__16260),
            .I(\b2v_inst11.count_clkZ0Z_2 ));
    InMux I__1821 (
            .O(N__16255),
            .I(N__16248));
    InMux I__1820 (
            .O(N__16254),
            .I(N__16248));
    InMux I__1819 (
            .O(N__16253),
            .I(N__16245));
    LocalMux I__1818 (
            .O(N__16248),
            .I(\b2v_inst11.count_clkZ0Z_3 ));
    LocalMux I__1817 (
            .O(N__16245),
            .I(\b2v_inst11.count_clkZ0Z_3 ));
    CascadeMux I__1816 (
            .O(N__16240),
            .I(\b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_ ));
    CascadeMux I__1815 (
            .O(N__16237),
            .I(N__16234));
    InMux I__1814 (
            .O(N__16234),
            .I(N__16228));
    InMux I__1813 (
            .O(N__16233),
            .I(N__16221));
    InMux I__1812 (
            .O(N__16232),
            .I(N__16221));
    InMux I__1811 (
            .O(N__16231),
            .I(N__16221));
    LocalMux I__1810 (
            .O(N__16228),
            .I(N__16218));
    LocalMux I__1809 (
            .O(N__16221),
            .I(\b2v_inst11.count_clkZ0Z_7 ));
    Odrv4 I__1808 (
            .O(N__16218),
            .I(\b2v_inst11.count_clkZ0Z_7 ));
    InMux I__1807 (
            .O(N__16213),
            .I(N__16210));
    LocalMux I__1806 (
            .O(N__16210),
            .I(\b2v_inst11.count_clk_0_0 ));
    InMux I__1805 (
            .O(N__16207),
            .I(N__16204));
    LocalMux I__1804 (
            .O(N__16204),
            .I(\b2v_inst11.count_clk_0_10 ));
    InMux I__1803 (
            .O(N__16201),
            .I(N__16195));
    InMux I__1802 (
            .O(N__16200),
            .I(N__16195));
    LocalMux I__1801 (
            .O(N__16195),
            .I(\b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5 ));
    CascadeMux I__1800 (
            .O(N__16192),
            .I(N__16189));
    InMux I__1799 (
            .O(N__16189),
            .I(N__16186));
    LocalMux I__1798 (
            .O(N__16186),
            .I(\b2v_inst11.count_clkZ0Z_10 ));
    CascadeMux I__1797 (
            .O(N__16183),
            .I(N__16179));
    InMux I__1796 (
            .O(N__16182),
            .I(N__16176));
    InMux I__1795 (
            .O(N__16179),
            .I(N__16173));
    LocalMux I__1794 (
            .O(N__16176),
            .I(\b2v_inst11.count_clkZ0Z_11 ));
    LocalMux I__1793 (
            .O(N__16173),
            .I(\b2v_inst11.count_clkZ0Z_11 ));
    CascadeMux I__1792 (
            .O(N__16168),
            .I(\b2v_inst11.count_clkZ0Z_10_cascade_ ));
    InMux I__1791 (
            .O(N__16165),
            .I(N__16161));
    InMux I__1790 (
            .O(N__16164),
            .I(N__16158));
    LocalMux I__1789 (
            .O(N__16161),
            .I(N__16155));
    LocalMux I__1788 (
            .O(N__16158),
            .I(\b2v_inst11.count_clkZ0Z_15 ));
    Odrv4 I__1787 (
            .O(N__16155),
            .I(\b2v_inst11.count_clkZ0Z_15 ));
    CascadeMux I__1786 (
            .O(N__16150),
            .I(\b2v_inst11.un2_count_clk_17_0_o2_1_4_cascade_ ));
    CascadeMux I__1785 (
            .O(N__16147),
            .I(N__16143));
    InMux I__1784 (
            .O(N__16146),
            .I(N__16140));
    InMux I__1783 (
            .O(N__16143),
            .I(N__16137));
    LocalMux I__1782 (
            .O(N__16140),
            .I(\b2v_inst11.count_clkZ0Z_14 ));
    LocalMux I__1781 (
            .O(N__16137),
            .I(\b2v_inst11.count_clkZ0Z_14 ));
    InMux I__1780 (
            .O(N__16132),
            .I(N__16129));
    LocalMux I__1779 (
            .O(N__16129),
            .I(\b2v_inst11.count_clk_0_13 ));
    InMux I__1778 (
            .O(N__16126),
            .I(N__16120));
    InMux I__1777 (
            .O(N__16125),
            .I(N__16120));
    LocalMux I__1776 (
            .O(N__16120),
            .I(\b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CAZ0 ));
    CascadeMux I__1775 (
            .O(N__16117),
            .I(N__16113));
    InMux I__1774 (
            .O(N__16116),
            .I(N__16110));
    InMux I__1773 (
            .O(N__16113),
            .I(N__16107));
    LocalMux I__1772 (
            .O(N__16110),
            .I(\b2v_inst11.count_clkZ0Z_13 ));
    LocalMux I__1771 (
            .O(N__16107),
            .I(\b2v_inst11.count_clkZ0Z_13 ));
    InMux I__1770 (
            .O(N__16102),
            .I(N__16096));
    InMux I__1769 (
            .O(N__16101),
            .I(N__16096));
    LocalMux I__1768 (
            .O(N__16096),
            .I(\b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DAZ0 ));
    InMux I__1767 (
            .O(N__16093),
            .I(N__16090));
    LocalMux I__1766 (
            .O(N__16090),
            .I(\b2v_inst11.count_clk_0_14 ));
    InMux I__1765 (
            .O(N__16087),
            .I(N__16083));
    InMux I__1764 (
            .O(N__16086),
            .I(N__16080));
    LocalMux I__1763 (
            .O(N__16083),
            .I(\b2v_inst200.countZ0Z_14 ));
    LocalMux I__1762 (
            .O(N__16080),
            .I(\b2v_inst200.countZ0Z_14 ));
    InMux I__1761 (
            .O(N__16075),
            .I(N__16069));
    InMux I__1760 (
            .O(N__16074),
            .I(N__16069));
    LocalMux I__1759 (
            .O(N__16069),
            .I(\b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59 ));
    InMux I__1758 (
            .O(N__16066),
            .I(\b2v_inst200.un2_count_1_cry_13 ));
    InMux I__1757 (
            .O(N__16063),
            .I(N__16059));
    InMux I__1756 (
            .O(N__16062),
            .I(N__16056));
    LocalMux I__1755 (
            .O(N__16059),
            .I(\b2v_inst200.countZ0Z_15 ));
    LocalMux I__1754 (
            .O(N__16056),
            .I(\b2v_inst200.countZ0Z_15 ));
    InMux I__1753 (
            .O(N__16051),
            .I(N__16048));
    LocalMux I__1752 (
            .O(N__16048),
            .I(N__16044));
    InMux I__1751 (
            .O(N__16047),
            .I(N__16041));
    Odrv12 I__1750 (
            .O(N__16044),
            .I(\b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69 ));
    LocalMux I__1749 (
            .O(N__16041),
            .I(\b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69 ));
    InMux I__1748 (
            .O(N__16036),
            .I(\b2v_inst200.un2_count_1_cry_14 ));
    InMux I__1747 (
            .O(N__16033),
            .I(N__16030));
    LocalMux I__1746 (
            .O(N__16030),
            .I(N__16027));
    Span4Mux_v I__1745 (
            .O(N__16027),
            .I(N__16023));
    InMux I__1744 (
            .O(N__16026),
            .I(N__16020));
    Odrv4 I__1743 (
            .O(N__16023),
            .I(\b2v_inst200.countZ0Z_16 ));
    LocalMux I__1742 (
            .O(N__16020),
            .I(\b2v_inst200.countZ0Z_16 ));
    InMux I__1741 (
            .O(N__16015),
            .I(N__16009));
    InMux I__1740 (
            .O(N__16014),
            .I(N__16009));
    LocalMux I__1739 (
            .O(N__16009),
            .I(N__16006));
    Odrv4 I__1738 (
            .O(N__16006),
            .I(\b2v_inst200.count_1_16 ));
    InMux I__1737 (
            .O(N__16003),
            .I(bfn_2_8_0_));
    InMux I__1736 (
            .O(N__16000),
            .I(N__15997));
    LocalMux I__1735 (
            .O(N__15997),
            .I(N__15993));
    InMux I__1734 (
            .O(N__15996),
            .I(N__15990));
    Odrv12 I__1733 (
            .O(N__15993),
            .I(\b2v_inst200.countZ0Z_17 ));
    LocalMux I__1732 (
            .O(N__15990),
            .I(\b2v_inst200.countZ0Z_17 ));
    InMux I__1731 (
            .O(N__15985),
            .I(\b2v_inst200.un2_count_1_cry_16 ));
    InMux I__1730 (
            .O(N__15982),
            .I(N__15976));
    InMux I__1729 (
            .O(N__15981),
            .I(N__15976));
    LocalMux I__1728 (
            .O(N__15976),
            .I(N__15973));
    Odrv4 I__1727 (
            .O(N__15973),
            .I(\b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ));
    InMux I__1726 (
            .O(N__15970),
            .I(N__15964));
    InMux I__1725 (
            .O(N__15969),
            .I(N__15964));
    LocalMux I__1724 (
            .O(N__15964),
            .I(\b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AAZ0 ));
    InMux I__1723 (
            .O(N__15961),
            .I(N__15958));
    LocalMux I__1722 (
            .O(N__15958),
            .I(\b2v_inst11.count_clk_0_11 ));
    CascadeMux I__1721 (
            .O(N__15955),
            .I(\b2v_inst11.count_clkZ0Z_0_cascade_ ));
    CascadeMux I__1720 (
            .O(N__15952),
            .I(N__15949));
    InMux I__1719 (
            .O(N__15949),
            .I(N__15945));
    InMux I__1718 (
            .O(N__15948),
            .I(N__15942));
    LocalMux I__1717 (
            .O(N__15945),
            .I(\b2v_inst200.countZ0Z_6 ));
    LocalMux I__1716 (
            .O(N__15942),
            .I(\b2v_inst200.countZ0Z_6 ));
    InMux I__1715 (
            .O(N__15937),
            .I(N__15933));
    InMux I__1714 (
            .O(N__15936),
            .I(N__15930));
    LocalMux I__1713 (
            .O(N__15933),
            .I(\b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0 ));
    LocalMux I__1712 (
            .O(N__15930),
            .I(\b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0 ));
    InMux I__1711 (
            .O(N__15925),
            .I(\b2v_inst200.un2_count_1_cry_5 ));
    InMux I__1710 (
            .O(N__15922),
            .I(N__15918));
    InMux I__1709 (
            .O(N__15921),
            .I(N__15915));
    LocalMux I__1708 (
            .O(N__15918),
            .I(\b2v_inst200.countZ0Z_7 ));
    LocalMux I__1707 (
            .O(N__15915),
            .I(\b2v_inst200.countZ0Z_7 ));
    InMux I__1706 (
            .O(N__15910),
            .I(N__15907));
    LocalMux I__1705 (
            .O(N__15907),
            .I(N__15903));
    InMux I__1704 (
            .O(N__15906),
            .I(N__15900));
    Odrv4 I__1703 (
            .O(N__15903),
            .I(\b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ));
    LocalMux I__1702 (
            .O(N__15900),
            .I(\b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ));
    InMux I__1701 (
            .O(N__15895),
            .I(\b2v_inst200.un2_count_1_cry_6 ));
    InMux I__1700 (
            .O(N__15892),
            .I(N__15888));
    InMux I__1699 (
            .O(N__15891),
            .I(N__15885));
    LocalMux I__1698 (
            .O(N__15888),
            .I(\b2v_inst200.countZ0Z_8 ));
    LocalMux I__1697 (
            .O(N__15885),
            .I(\b2v_inst200.countZ0Z_8 ));
    CascadeMux I__1696 (
            .O(N__15880),
            .I(N__15877));
    InMux I__1695 (
            .O(N__15877),
            .I(N__15871));
    InMux I__1694 (
            .O(N__15876),
            .I(N__15871));
    LocalMux I__1693 (
            .O(N__15871),
            .I(\b2v_inst200.un2_count_1_cry_7_c_RNIP33EZ0 ));
    InMux I__1692 (
            .O(N__15868),
            .I(bfn_2_7_0_));
    InMux I__1691 (
            .O(N__15865),
            .I(N__15862));
    LocalMux I__1690 (
            .O(N__15862),
            .I(\b2v_inst200.countZ0Z_9 ));
    InMux I__1689 (
            .O(N__15859),
            .I(N__15853));
    InMux I__1688 (
            .O(N__15858),
            .I(N__15853));
    LocalMux I__1687 (
            .O(N__15853),
            .I(\b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0 ));
    InMux I__1686 (
            .O(N__15850),
            .I(\b2v_inst200.un2_count_1_cry_8 ));
    InMux I__1685 (
            .O(N__15847),
            .I(N__15844));
    LocalMux I__1684 (
            .O(N__15844),
            .I(N__15840));
    InMux I__1683 (
            .O(N__15843),
            .I(N__15837));
    Odrv4 I__1682 (
            .O(N__15840),
            .I(\b2v_inst200.countZ0Z_10 ));
    LocalMux I__1681 (
            .O(N__15837),
            .I(\b2v_inst200.countZ0Z_10 ));
    CascadeMux I__1680 (
            .O(N__15832),
            .I(N__15829));
    InMux I__1679 (
            .O(N__15829),
            .I(N__15823));
    InMux I__1678 (
            .O(N__15828),
            .I(N__15823));
    LocalMux I__1677 (
            .O(N__15823),
            .I(N__15820));
    Odrv4 I__1676 (
            .O(N__15820),
            .I(\b2v_inst200.un2_count_1_cry_9_c_RNIR75EZ0 ));
    InMux I__1675 (
            .O(N__15817),
            .I(\b2v_inst200.un2_count_1_cry_9 ));
    InMux I__1674 (
            .O(N__15814),
            .I(N__15810));
    CascadeMux I__1673 (
            .O(N__15813),
            .I(N__15807));
    LocalMux I__1672 (
            .O(N__15810),
            .I(N__15804));
    InMux I__1671 (
            .O(N__15807),
            .I(N__15801));
    Odrv4 I__1670 (
            .O(N__15804),
            .I(\b2v_inst200.countZ0Z_11 ));
    LocalMux I__1669 (
            .O(N__15801),
            .I(\b2v_inst200.countZ0Z_11 ));
    InMux I__1668 (
            .O(N__15796),
            .I(N__15790));
    InMux I__1667 (
            .O(N__15795),
            .I(N__15790));
    LocalMux I__1666 (
            .O(N__15790),
            .I(N__15787));
    Odrv4 I__1665 (
            .O(N__15787),
            .I(\b2v_inst200.un2_count_1_cry_10_c_RNI3AZ0Z29 ));
    InMux I__1664 (
            .O(N__15784),
            .I(\b2v_inst200.un2_count_1_cry_10 ));
    InMux I__1663 (
            .O(N__15781),
            .I(N__15777));
    InMux I__1662 (
            .O(N__15780),
            .I(N__15774));
    LocalMux I__1661 (
            .O(N__15777),
            .I(\b2v_inst200.countZ0Z_12 ));
    LocalMux I__1660 (
            .O(N__15774),
            .I(\b2v_inst200.countZ0Z_12 ));
    InMux I__1659 (
            .O(N__15769),
            .I(N__15763));
    InMux I__1658 (
            .O(N__15768),
            .I(N__15763));
    LocalMux I__1657 (
            .O(N__15763),
            .I(\b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39 ));
    InMux I__1656 (
            .O(N__15760),
            .I(\b2v_inst200.un2_count_1_cry_11 ));
    InMux I__1655 (
            .O(N__15757),
            .I(N__15753));
    InMux I__1654 (
            .O(N__15756),
            .I(N__15750));
    LocalMux I__1653 (
            .O(N__15753),
            .I(\b2v_inst200.countZ0Z_13 ));
    LocalMux I__1652 (
            .O(N__15750),
            .I(\b2v_inst200.countZ0Z_13 ));
    InMux I__1651 (
            .O(N__15745),
            .I(N__15739));
    InMux I__1650 (
            .O(N__15744),
            .I(N__15739));
    LocalMux I__1649 (
            .O(N__15739),
            .I(\b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49 ));
    InMux I__1648 (
            .O(N__15736),
            .I(\b2v_inst200.un2_count_1_cry_12 ));
    InMux I__1647 (
            .O(N__15733),
            .I(N__15730));
    LocalMux I__1646 (
            .O(N__15730),
            .I(\b2v_inst200.count_2_1 ));
    InMux I__1645 (
            .O(N__15727),
            .I(N__15724));
    LocalMux I__1644 (
            .O(N__15724),
            .I(\b2v_inst200.count_2_2 ));
    InMux I__1643 (
            .O(N__15721),
            .I(N__15701));
    InMux I__1642 (
            .O(N__15720),
            .I(N__15696));
    InMux I__1641 (
            .O(N__15719),
            .I(N__15696));
    InMux I__1640 (
            .O(N__15718),
            .I(N__15689));
    InMux I__1639 (
            .O(N__15717),
            .I(N__15689));
    InMux I__1638 (
            .O(N__15716),
            .I(N__15689));
    InMux I__1637 (
            .O(N__15715),
            .I(N__15680));
    InMux I__1636 (
            .O(N__15714),
            .I(N__15680));
    InMux I__1635 (
            .O(N__15713),
            .I(N__15680));
    InMux I__1634 (
            .O(N__15712),
            .I(N__15680));
    InMux I__1633 (
            .O(N__15711),
            .I(N__15671));
    InMux I__1632 (
            .O(N__15710),
            .I(N__15671));
    InMux I__1631 (
            .O(N__15709),
            .I(N__15671));
    InMux I__1630 (
            .O(N__15708),
            .I(N__15671));
    InMux I__1629 (
            .O(N__15707),
            .I(N__15662));
    InMux I__1628 (
            .O(N__15706),
            .I(N__15662));
    InMux I__1627 (
            .O(N__15705),
            .I(N__15662));
    InMux I__1626 (
            .O(N__15704),
            .I(N__15662));
    LocalMux I__1625 (
            .O(N__15701),
            .I(N__15653));
    LocalMux I__1624 (
            .O(N__15696),
            .I(N__15650));
    LocalMux I__1623 (
            .O(N__15689),
            .I(N__15647));
    LocalMux I__1622 (
            .O(N__15680),
            .I(N__15644));
    LocalMux I__1621 (
            .O(N__15671),
            .I(N__15641));
    LocalMux I__1620 (
            .O(N__15662),
            .I(N__15638));
    CEMux I__1619 (
            .O(N__15661),
            .I(N__15613));
    CEMux I__1618 (
            .O(N__15660),
            .I(N__15613));
    CEMux I__1617 (
            .O(N__15659),
            .I(N__15613));
    CEMux I__1616 (
            .O(N__15658),
            .I(N__15613));
    CEMux I__1615 (
            .O(N__15657),
            .I(N__15613));
    CEMux I__1614 (
            .O(N__15656),
            .I(N__15613));
    Glb2LocalMux I__1613 (
            .O(N__15653),
            .I(N__15613));
    Glb2LocalMux I__1612 (
            .O(N__15650),
            .I(N__15613));
    Glb2LocalMux I__1611 (
            .O(N__15647),
            .I(N__15613));
    Glb2LocalMux I__1610 (
            .O(N__15644),
            .I(N__15613));
    Glb2LocalMux I__1609 (
            .O(N__15641),
            .I(N__15613));
    Glb2LocalMux I__1608 (
            .O(N__15638),
            .I(N__15613));
    GlobalMux I__1607 (
            .O(N__15613),
            .I(N__15610));
    gio2CtrlBuf I__1606 (
            .O(N__15610),
            .I(\b2v_inst200.count_en_g ));
    InMux I__1605 (
            .O(N__15607),
            .I(N__15603));
    InMux I__1604 (
            .O(N__15606),
            .I(N__15600));
    LocalMux I__1603 (
            .O(N__15603),
            .I(\b2v_inst200.countZ0Z_0 ));
    LocalMux I__1602 (
            .O(N__15600),
            .I(\b2v_inst200.countZ0Z_0 ));
    InMux I__1601 (
            .O(N__15595),
            .I(N__15592));
    LocalMux I__1600 (
            .O(N__15592),
            .I(\b2v_inst200.count_1_0 ));
    CascadeMux I__1599 (
            .O(N__15589),
            .I(N__15586));
    InMux I__1598 (
            .O(N__15586),
            .I(N__15582));
    InMux I__1597 (
            .O(N__15585),
            .I(N__15579));
    LocalMux I__1596 (
            .O(N__15582),
            .I(\b2v_inst200.countZ0Z_1 ));
    LocalMux I__1595 (
            .O(N__15579),
            .I(\b2v_inst200.countZ0Z_1 ));
    InMux I__1594 (
            .O(N__15574),
            .I(N__15568));
    InMux I__1593 (
            .O(N__15573),
            .I(N__15568));
    LocalMux I__1592 (
            .O(N__15568),
            .I(\b2v_inst200.count_RNIC03N_5Z0Z_0 ));
    InMux I__1591 (
            .O(N__15565),
            .I(\b2v_inst200.un2_count_1_cry_1_cy ));
    InMux I__1590 (
            .O(N__15562),
            .I(N__15558));
    InMux I__1589 (
            .O(N__15561),
            .I(N__15555));
    LocalMux I__1588 (
            .O(N__15558),
            .I(\b2v_inst200.countZ0Z_2 ));
    LocalMux I__1587 (
            .O(N__15555),
            .I(\b2v_inst200.countZ0Z_2 ));
    InMux I__1586 (
            .O(N__15550),
            .I(N__15546));
    InMux I__1585 (
            .O(N__15549),
            .I(N__15543));
    LocalMux I__1584 (
            .O(N__15546),
            .I(N__15540));
    LocalMux I__1583 (
            .O(N__15543),
            .I(\b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ));
    Odrv4 I__1582 (
            .O(N__15540),
            .I(\b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ));
    InMux I__1581 (
            .O(N__15535),
            .I(\b2v_inst200.un2_count_1_cry_1 ));
    InMux I__1580 (
            .O(N__15532),
            .I(N__15528));
    InMux I__1579 (
            .O(N__15531),
            .I(N__15525));
    LocalMux I__1578 (
            .O(N__15528),
            .I(\b2v_inst200.countZ0Z_3 ));
    LocalMux I__1577 (
            .O(N__15525),
            .I(\b2v_inst200.countZ0Z_3 ));
    InMux I__1576 (
            .O(N__15520),
            .I(N__15514));
    InMux I__1575 (
            .O(N__15519),
            .I(N__15514));
    LocalMux I__1574 (
            .O(N__15514),
            .I(\b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0 ));
    InMux I__1573 (
            .O(N__15511),
            .I(\b2v_inst200.un2_count_1_cry_2 ));
    CascadeMux I__1572 (
            .O(N__15508),
            .I(N__15505));
    InMux I__1571 (
            .O(N__15505),
            .I(N__15501));
    InMux I__1570 (
            .O(N__15504),
            .I(N__15498));
    LocalMux I__1569 (
            .O(N__15501),
            .I(\b2v_inst200.countZ0Z_4 ));
    LocalMux I__1568 (
            .O(N__15498),
            .I(\b2v_inst200.countZ0Z_4 ));
    InMux I__1567 (
            .O(N__15493),
            .I(N__15487));
    InMux I__1566 (
            .O(N__15492),
            .I(N__15487));
    LocalMux I__1565 (
            .O(N__15487),
            .I(\b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ));
    InMux I__1564 (
            .O(N__15484),
            .I(\b2v_inst200.un2_count_1_cry_3 ));
    InMux I__1563 (
            .O(N__15481),
            .I(N__15477));
    InMux I__1562 (
            .O(N__15480),
            .I(N__15474));
    LocalMux I__1561 (
            .O(N__15477),
            .I(\b2v_inst200.countZ0Z_5 ));
    LocalMux I__1560 (
            .O(N__15474),
            .I(\b2v_inst200.countZ0Z_5 ));
    InMux I__1559 (
            .O(N__15469),
            .I(N__15463));
    InMux I__1558 (
            .O(N__15468),
            .I(N__15463));
    LocalMux I__1557 (
            .O(N__15463),
            .I(\b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ));
    InMux I__1556 (
            .O(N__15460),
            .I(\b2v_inst200.un2_count_1_cry_4 ));
    InMux I__1555 (
            .O(N__15457),
            .I(N__15454));
    LocalMux I__1554 (
            .O(N__15454),
            .I(N__15451));
    Span4Mux_v I__1553 (
            .O(N__15451),
            .I(N__15448));
    Odrv4 I__1552 (
            .O(N__15448),
            .I(\b2v_inst200.count_2_15 ));
    InMux I__1551 (
            .O(N__15445),
            .I(N__15442));
    LocalMux I__1550 (
            .O(N__15442),
            .I(N__15439));
    Span4Mux_s1_h I__1549 (
            .O(N__15439),
            .I(N__15436));
    Odrv4 I__1548 (
            .O(N__15436),
            .I(\b2v_inst200.count_2_7 ));
    InMux I__1547 (
            .O(N__15433),
            .I(N__15430));
    LocalMux I__1546 (
            .O(N__15430),
            .I(\b2v_inst200.un25_clk_100khz_11 ));
    InMux I__1545 (
            .O(N__15427),
            .I(N__15424));
    LocalMux I__1544 (
            .O(N__15424),
            .I(\b2v_inst200.count_0_16 ));
    InMux I__1543 (
            .O(N__15421),
            .I(N__15418));
    LocalMux I__1542 (
            .O(N__15418),
            .I(\b2v_inst200.count_0_17 ));
    CascadeMux I__1541 (
            .O(N__15415),
            .I(\b2v_inst16.un13_clk_100khz_i_cascade_ ));
    InMux I__1540 (
            .O(N__15412),
            .I(N__15409));
    LocalMux I__1539 (
            .O(N__15409),
            .I(\b2v_inst16.count_4_0 ));
    CascadeMux I__1538 (
            .O(N__15406),
            .I(\b2v_inst16.count_rst_5_cascade_ ));
    InMux I__1537 (
            .O(N__15403),
            .I(N__15400));
    LocalMux I__1536 (
            .O(N__15400),
            .I(\b2v_inst16.count_4_13 ));
    InMux I__1535 (
            .O(N__15397),
            .I(N__15391));
    InMux I__1534 (
            .O(N__15396),
            .I(N__15391));
    LocalMux I__1533 (
            .O(N__15391),
            .I(\b2v_inst16.count_rst_2 ));
    InMux I__1532 (
            .O(N__15388),
            .I(N__15385));
    LocalMux I__1531 (
            .O(N__15385),
            .I(\b2v_inst16.countZ0Z_13 ));
    InMux I__1530 (
            .O(N__15382),
            .I(N__15372));
    InMux I__1529 (
            .O(N__15381),
            .I(N__15372));
    InMux I__1528 (
            .O(N__15380),
            .I(N__15369));
    InMux I__1527 (
            .O(N__15379),
            .I(N__15362));
    InMux I__1526 (
            .O(N__15378),
            .I(N__15362));
    InMux I__1525 (
            .O(N__15377),
            .I(N__15362));
    LocalMux I__1524 (
            .O(N__15372),
            .I(\b2v_inst16.countZ0Z_0 ));
    LocalMux I__1523 (
            .O(N__15369),
            .I(\b2v_inst16.countZ0Z_0 ));
    LocalMux I__1522 (
            .O(N__15362),
            .I(\b2v_inst16.countZ0Z_0 ));
    CascadeMux I__1521 (
            .O(N__15355),
            .I(\b2v_inst16.countZ0Z_13_cascade_ ));
    InMux I__1520 (
            .O(N__15352),
            .I(N__15349));
    LocalMux I__1519 (
            .O(N__15349),
            .I(\b2v_inst16.un13_clk_100khz_11 ));
    InMux I__1518 (
            .O(N__15346),
            .I(N__15342));
    InMux I__1517 (
            .O(N__15345),
            .I(N__15339));
    LocalMux I__1516 (
            .O(N__15342),
            .I(\b2v_inst16.countZ0Z_15 ));
    LocalMux I__1515 (
            .O(N__15339),
            .I(\b2v_inst16.countZ0Z_15 ));
    InMux I__1514 (
            .O(N__15334),
            .I(N__15328));
    InMux I__1513 (
            .O(N__15333),
            .I(N__15328));
    LocalMux I__1512 (
            .O(N__15328),
            .I(\b2v_inst16.count_rst_4 ));
    InMux I__1511 (
            .O(N__15325),
            .I(N__15322));
    LocalMux I__1510 (
            .O(N__15322),
            .I(\b2v_inst16.count_4_15 ));
    InMux I__1509 (
            .O(N__15319),
            .I(N__15316));
    LocalMux I__1508 (
            .O(N__15316),
            .I(\b2v_inst16.count_4_14 ));
    InMux I__1507 (
            .O(N__15313),
            .I(N__15309));
    InMux I__1506 (
            .O(N__15312),
            .I(N__15306));
    LocalMux I__1505 (
            .O(N__15309),
            .I(\b2v_inst16.count_rst_3 ));
    LocalMux I__1504 (
            .O(N__15306),
            .I(\b2v_inst16.count_rst_3 ));
    InMux I__1503 (
            .O(N__15301),
            .I(N__15297));
    InMux I__1502 (
            .O(N__15300),
            .I(N__15294));
    LocalMux I__1501 (
            .O(N__15297),
            .I(\b2v_inst16.countZ0Z_14 ));
    LocalMux I__1500 (
            .O(N__15294),
            .I(\b2v_inst16.countZ0Z_14 ));
    InMux I__1499 (
            .O(N__15289),
            .I(N__15285));
    InMux I__1498 (
            .O(N__15288),
            .I(N__15282));
    LocalMux I__1497 (
            .O(N__15285),
            .I(\b2v_inst16.count_rst_12 ));
    LocalMux I__1496 (
            .O(N__15282),
            .I(\b2v_inst16.count_rst_12 ));
    InMux I__1495 (
            .O(N__15277),
            .I(N__15274));
    LocalMux I__1494 (
            .O(N__15274),
            .I(\b2v_inst16.count_4_7 ));
    InMux I__1493 (
            .O(N__15271),
            .I(N__15267));
    InMux I__1492 (
            .O(N__15270),
            .I(N__15264));
    LocalMux I__1491 (
            .O(N__15267),
            .I(\b2v_inst16.count_rst_9 ));
    LocalMux I__1490 (
            .O(N__15264),
            .I(\b2v_inst16.count_rst_9 ));
    InMux I__1489 (
            .O(N__15259),
            .I(N__15256));
    LocalMux I__1488 (
            .O(N__15256),
            .I(\b2v_inst16.count_4_4 ));
    CascadeMux I__1487 (
            .O(N__15253),
            .I(\b2v_inst16.count_rst_6_cascade_ ));
    InMux I__1486 (
            .O(N__15250),
            .I(N__15247));
    LocalMux I__1485 (
            .O(N__15247),
            .I(\b2v_inst16.count_rst_6 ));
    InMux I__1484 (
            .O(N__15244),
            .I(N__15241));
    LocalMux I__1483 (
            .O(N__15241),
            .I(N__15237));
    InMux I__1482 (
            .O(N__15240),
            .I(N__15234));
    Odrv4 I__1481 (
            .O(N__15237),
            .I(\b2v_inst16.countZ0Z_11 ));
    LocalMux I__1480 (
            .O(N__15234),
            .I(\b2v_inst16.countZ0Z_11 ));
    CascadeMux I__1479 (
            .O(N__15229),
            .I(\b2v_inst16.countZ0Z_1_cascade_ ));
    CascadeMux I__1478 (
            .O(N__15226),
            .I(N__15223));
    InMux I__1477 (
            .O(N__15223),
            .I(N__15218));
    InMux I__1476 (
            .O(N__15222),
            .I(N__15213));
    InMux I__1475 (
            .O(N__15221),
            .I(N__15213));
    LocalMux I__1474 (
            .O(N__15218),
            .I(N__15210));
    LocalMux I__1473 (
            .O(N__15213),
            .I(\b2v_inst16.un4_count_1_axb_1 ));
    Odrv4 I__1472 (
            .O(N__15210),
            .I(\b2v_inst16.un4_count_1_axb_1 ));
    InMux I__1471 (
            .O(N__15205),
            .I(N__15199));
    InMux I__1470 (
            .O(N__15204),
            .I(N__15199));
    LocalMux I__1469 (
            .O(N__15199),
            .I(\b2v_inst16.count_4_1 ));
    InMux I__1468 (
            .O(N__15196),
            .I(N__15193));
    LocalMux I__1467 (
            .O(N__15193),
            .I(N__15189));
    InMux I__1466 (
            .O(N__15192),
            .I(N__15186));
    Span4Mux_s1_v I__1465 (
            .O(N__15189),
            .I(N__15183));
    LocalMux I__1464 (
            .O(N__15186),
            .I(N__15180));
    Odrv4 I__1463 (
            .O(N__15183),
            .I(\b2v_inst16.countZ0Z_2 ));
    Odrv4 I__1462 (
            .O(N__15180),
            .I(\b2v_inst16.countZ0Z_2 ));
    CascadeMux I__1461 (
            .O(N__15175),
            .I(N__15172));
    InMux I__1460 (
            .O(N__15172),
            .I(N__15168));
    InMux I__1459 (
            .O(N__15171),
            .I(N__15165));
    LocalMux I__1458 (
            .O(N__15168),
            .I(N__15162));
    LocalMux I__1457 (
            .O(N__15165),
            .I(N__15159));
    Odrv4 I__1456 (
            .O(N__15162),
            .I(\b2v_inst16.countZ0Z_6 ));
    Odrv4 I__1455 (
            .O(N__15159),
            .I(\b2v_inst16.countZ0Z_6 ));
    InMux I__1454 (
            .O(N__15154),
            .I(N__15151));
    LocalMux I__1453 (
            .O(N__15151),
            .I(N__15147));
    InMux I__1452 (
            .O(N__15150),
            .I(N__15144));
    Odrv4 I__1451 (
            .O(N__15147),
            .I(\b2v_inst16.countZ0Z_12 ));
    LocalMux I__1450 (
            .O(N__15144),
            .I(\b2v_inst16.countZ0Z_12 ));
    InMux I__1449 (
            .O(N__15139),
            .I(N__15136));
    LocalMux I__1448 (
            .O(N__15136),
            .I(\b2v_inst16.un13_clk_100khz_9 ));
    InMux I__1447 (
            .O(N__15133),
            .I(N__15130));
    LocalMux I__1446 (
            .O(N__15130),
            .I(\b2v_inst16.un13_clk_100khz_8 ));
    CascadeMux I__1445 (
            .O(N__15127),
            .I(\b2v_inst16.un13_clk_100khz_10_cascade_ ));
    CascadeMux I__1444 (
            .O(N__15124),
            .I(\b2v_inst11.count_off_1_3_cascade_ ));
    CascadeMux I__1443 (
            .O(N__15121),
            .I(N__15118));
    InMux I__1442 (
            .O(N__15118),
            .I(N__15115));
    LocalMux I__1441 (
            .O(N__15115),
            .I(N__15112));
    Odrv4 I__1440 (
            .O(N__15112),
            .I(\b2v_inst11.un3_count_off_1_axb_3 ));
    CascadeMux I__1439 (
            .O(N__15109),
            .I(N__15106));
    InMux I__1438 (
            .O(N__15106),
            .I(N__15103));
    LocalMux I__1437 (
            .O(N__15103),
            .I(N__15100));
    Odrv4 I__1436 (
            .O(N__15100),
            .I(\b2v_inst11.count_offZ0Z_4 ));
    InMux I__1435 (
            .O(N__15097),
            .I(N__15094));
    LocalMux I__1434 (
            .O(N__15094),
            .I(\b2v_inst11.count_off_1_3 ));
    CascadeMux I__1433 (
            .O(N__15091),
            .I(\b2v_inst11.count_offZ0Z_4_cascade_ ));
    InMux I__1432 (
            .O(N__15088),
            .I(N__15085));
    LocalMux I__1431 (
            .O(N__15085),
            .I(N__15082));
    Odrv4 I__1430 (
            .O(N__15082),
            .I(\b2v_inst11.un34_clk_100khz_2 ));
    InMux I__1429 (
            .O(N__15079),
            .I(N__15073));
    InMux I__1428 (
            .O(N__15078),
            .I(N__15073));
    LocalMux I__1427 (
            .O(N__15073),
            .I(N__15070));
    Odrv4 I__1426 (
            .O(N__15070),
            .I(\b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362 ));
    InMux I__1425 (
            .O(N__15067),
            .I(N__15061));
    InMux I__1424 (
            .O(N__15066),
            .I(N__15061));
    LocalMux I__1423 (
            .O(N__15061),
            .I(\b2v_inst11.count_offZ0Z_3 ));
    InMux I__1422 (
            .O(N__15058),
            .I(N__15052));
    InMux I__1421 (
            .O(N__15057),
            .I(N__15052));
    LocalMux I__1420 (
            .O(N__15052),
            .I(N__15049));
    Odrv4 I__1419 (
            .O(N__15049),
            .I(\b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672 ));
    CascadeMux I__1418 (
            .O(N__15046),
            .I(N__15043));
    InMux I__1417 (
            .O(N__15043),
            .I(N__15040));
    LocalMux I__1416 (
            .O(N__15040),
            .I(\b2v_inst11.count_off_0_4 ));
    CascadeMux I__1415 (
            .O(N__15037),
            .I(N__15034));
    InMux I__1414 (
            .O(N__15034),
            .I(N__15031));
    LocalMux I__1413 (
            .O(N__15031),
            .I(\b2v_inst11.count_off_0_14 ));
    CascadeMux I__1412 (
            .O(N__15028),
            .I(N__15025));
    InMux I__1411 (
            .O(N__15025),
            .I(N__15019));
    InMux I__1410 (
            .O(N__15024),
            .I(N__15019));
    LocalMux I__1409 (
            .O(N__15019),
            .I(\b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5 ));
    InMux I__1408 (
            .O(N__15016),
            .I(\b2v_inst11.un3_count_off_1_cry_6 ));
    InMux I__1407 (
            .O(N__15013),
            .I(\b2v_inst11.un3_count_off_1_cry_7 ));
    InMux I__1406 (
            .O(N__15010),
            .I(bfn_1_15_0_));
    InMux I__1405 (
            .O(N__15007),
            .I(\b2v_inst11.un3_count_off_1_cry_9 ));
    InMux I__1404 (
            .O(N__15004),
            .I(\b2v_inst11.un3_count_off_1_cry_10 ));
    InMux I__1403 (
            .O(N__15001),
            .I(\b2v_inst11.un3_count_off_1_cry_11 ));
    InMux I__1402 (
            .O(N__14998),
            .I(\b2v_inst11.un3_count_off_1_cry_12 ));
    InMux I__1401 (
            .O(N__14995),
            .I(\b2v_inst11.un3_count_off_1_cry_13 ));
    InMux I__1400 (
            .O(N__14992),
            .I(\b2v_inst11.un3_count_off_1_cry_14 ));
    CascadeMux I__1399 (
            .O(N__14989),
            .I(\b2v_inst11.un34_clk_100khz_1_cascade_ ));
    InMux I__1398 (
            .O(N__14986),
            .I(N__14983));
    LocalMux I__1397 (
            .O(N__14983),
            .I(\b2v_inst11.un34_clk_100khz_0 ));
    InMux I__1396 (
            .O(N__14980),
            .I(N__14977));
    LocalMux I__1395 (
            .O(N__14977),
            .I(\b2v_inst11.count_off_0_5 ));
    InMux I__1394 (
            .O(N__14974),
            .I(N__14971));
    LocalMux I__1393 (
            .O(N__14971),
            .I(\b2v_inst11.un3_count_off_1_axb_2 ));
    InMux I__1392 (
            .O(N__14968),
            .I(N__14962));
    InMux I__1391 (
            .O(N__14967),
            .I(N__14962));
    LocalMux I__1390 (
            .O(N__14962),
            .I(\b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152 ));
    InMux I__1389 (
            .O(N__14959),
            .I(\b2v_inst11.un3_count_off_1_cry_1 ));
    InMux I__1388 (
            .O(N__14956),
            .I(\b2v_inst11.un3_count_off_1_cry_2_cZ0 ));
    InMux I__1387 (
            .O(N__14953),
            .I(\b2v_inst11.un3_count_off_1_cry_3_cZ0 ));
    CascadeMux I__1386 (
            .O(N__14950),
            .I(N__14946));
    InMux I__1385 (
            .O(N__14949),
            .I(N__14943));
    InMux I__1384 (
            .O(N__14946),
            .I(N__14940));
    LocalMux I__1383 (
            .O(N__14943),
            .I(\b2v_inst11.count_offZ0Z_5 ));
    LocalMux I__1382 (
            .O(N__14940),
            .I(\b2v_inst11.count_offZ0Z_5 ));
    InMux I__1381 (
            .O(N__14935),
            .I(N__14929));
    InMux I__1380 (
            .O(N__14934),
            .I(N__14929));
    LocalMux I__1379 (
            .O(N__14929),
            .I(\b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882 ));
    InMux I__1378 (
            .O(N__14926),
            .I(\b2v_inst11.un3_count_off_1_cry_4_cZ0 ));
    CascadeMux I__1377 (
            .O(N__14923),
            .I(N__14920));
    InMux I__1376 (
            .O(N__14920),
            .I(N__14917));
    LocalMux I__1375 (
            .O(N__14917),
            .I(N__14914));
    Odrv4 I__1374 (
            .O(N__14914),
            .I(\b2v_inst11.un3_count_off_1_axb_6 ));
    InMux I__1373 (
            .O(N__14911),
            .I(\b2v_inst11.un3_count_off_1_cry_5 ));
    InMux I__1372 (
            .O(N__14908),
            .I(N__14902));
    InMux I__1371 (
            .O(N__14907),
            .I(N__14902));
    LocalMux I__1370 (
            .O(N__14902),
            .I(N__14899));
    Odrv4 I__1369 (
            .O(N__14899),
            .I(\b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5 ));
    InMux I__1368 (
            .O(N__14896),
            .I(N__14893));
    LocalMux I__1367 (
            .O(N__14893),
            .I(\b2v_inst11.count_clk_0_4 ));
    InMux I__1366 (
            .O(N__14890),
            .I(N__14887));
    LocalMux I__1365 (
            .O(N__14887),
            .I(\b2v_inst11.count_off_1_2 ));
    InMux I__1364 (
            .O(N__14884),
            .I(N__14878));
    InMux I__1363 (
            .O(N__14883),
            .I(N__14878));
    LocalMux I__1362 (
            .O(N__14878),
            .I(\b2v_inst11.count_offZ0Z_2 ));
    CascadeMux I__1361 (
            .O(N__14875),
            .I(\b2v_inst11.count_off_1_2_cascade_ ));
    InMux I__1360 (
            .O(N__14872),
            .I(N__14869));
    LocalMux I__1359 (
            .O(N__14869),
            .I(N__14865));
    InMux I__1358 (
            .O(N__14868),
            .I(N__14862));
    Odrv4 I__1357 (
            .O(N__14865),
            .I(\b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0 ));
    LocalMux I__1356 (
            .O(N__14862),
            .I(\b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0 ));
    InMux I__1355 (
            .O(N__14857),
            .I(N__14854));
    LocalMux I__1354 (
            .O(N__14854),
            .I(\b2v_inst11.count_clk_0_15 ));
    InMux I__1353 (
            .O(N__14851),
            .I(N__14845));
    InMux I__1352 (
            .O(N__14850),
            .I(N__14845));
    LocalMux I__1351 (
            .O(N__14845),
            .I(N__14842));
    Odrv4 I__1350 (
            .O(N__14842),
            .I(\b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ));
    InMux I__1349 (
            .O(N__14839),
            .I(N__14836));
    LocalMux I__1348 (
            .O(N__14836),
            .I(\b2v_inst11.count_clk_0_6 ));
    CascadeMux I__1347 (
            .O(N__14833),
            .I(N__14829));
    InMux I__1346 (
            .O(N__14832),
            .I(N__14824));
    InMux I__1345 (
            .O(N__14829),
            .I(N__14824));
    LocalMux I__1344 (
            .O(N__14824),
            .I(N__14821));
    Odrv4 I__1343 (
            .O(N__14821),
            .I(\b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5 ));
    InMux I__1342 (
            .O(N__14818),
            .I(N__14815));
    LocalMux I__1341 (
            .O(N__14815),
            .I(\b2v_inst11.count_clk_0_8 ));
    CascadeMux I__1340 (
            .O(N__14812),
            .I(N__14808));
    InMux I__1339 (
            .O(N__14811),
            .I(N__14803));
    InMux I__1338 (
            .O(N__14808),
            .I(N__14803));
    LocalMux I__1337 (
            .O(N__14803),
            .I(N__14800));
    Odrv4 I__1336 (
            .O(N__14800),
            .I(\b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5 ));
    InMux I__1335 (
            .O(N__14797),
            .I(N__14794));
    LocalMux I__1334 (
            .O(N__14794),
            .I(\b2v_inst11.count_clk_0_7 ));
    InMux I__1333 (
            .O(N__14791),
            .I(N__14785));
    InMux I__1332 (
            .O(N__14790),
            .I(N__14785));
    LocalMux I__1331 (
            .O(N__14785),
            .I(N__14782));
    Odrv4 I__1330 (
            .O(N__14782),
            .I(\b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5 ));
    InMux I__1329 (
            .O(N__14779),
            .I(N__14776));
    LocalMux I__1328 (
            .O(N__14776),
            .I(\b2v_inst11.count_clk_0_9 ));
    InMux I__1327 (
            .O(N__14773),
            .I(\b2v_inst11.un1_count_clk_2_cry_9_cZ0 ));
    InMux I__1326 (
            .O(N__14770),
            .I(\b2v_inst11.un1_count_clk_2_cry_10_cZ0 ));
    InMux I__1325 (
            .O(N__14767),
            .I(\b2v_inst11.un1_count_clk_2_cry_11 ));
    InMux I__1324 (
            .O(N__14764),
            .I(\b2v_inst11.un1_count_clk_2_cry_12 ));
    InMux I__1323 (
            .O(N__14761),
            .I(\b2v_inst11.un1_count_clk_2_cry_13 ));
    InMux I__1322 (
            .O(N__14758),
            .I(\b2v_inst11.un1_count_clk_2_cry_14 ));
    InMux I__1321 (
            .O(N__14755),
            .I(N__14749));
    InMux I__1320 (
            .O(N__14754),
            .I(N__14749));
    LocalMux I__1319 (
            .O(N__14749),
            .I(N__14746));
    Odrv4 I__1318 (
            .O(N__14746),
            .I(\b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5 ));
    InMux I__1317 (
            .O(N__14743),
            .I(N__14740));
    LocalMux I__1316 (
            .O(N__14740),
            .I(\b2v_inst11.count_clk_0_5 ));
    InMux I__1315 (
            .O(N__14737),
            .I(\b2v_inst11.un1_count_clk_2_cry_1 ));
    InMux I__1314 (
            .O(N__14734),
            .I(\b2v_inst11.un1_count_clk_2_cry_2 ));
    InMux I__1313 (
            .O(N__14731),
            .I(\b2v_inst11.un1_count_clk_2_cry_3 ));
    InMux I__1312 (
            .O(N__14728),
            .I(\b2v_inst11.un1_count_clk_2_cry_4 ));
    InMux I__1311 (
            .O(N__14725),
            .I(\b2v_inst11.un1_count_clk_2_cry_5 ));
    InMux I__1310 (
            .O(N__14722),
            .I(\b2v_inst11.un1_count_clk_2_cry_6 ));
    InMux I__1309 (
            .O(N__14719),
            .I(\b2v_inst11.un1_count_clk_2_cry_7_cZ0 ));
    InMux I__1308 (
            .O(N__14716),
            .I(bfn_1_10_0_));
    InMux I__1307 (
            .O(N__14713),
            .I(N__14710));
    LocalMux I__1306 (
            .O(N__14710),
            .I(\b2v_inst200.count_2_5 ));
    InMux I__1305 (
            .O(N__14707),
            .I(N__14704));
    LocalMux I__1304 (
            .O(N__14704),
            .I(\b2v_inst200.count_2_9 ));
    CascadeMux I__1303 (
            .O(N__14701),
            .I(\b2v_inst200.countZ0Z_9_cascade_ ));
    InMux I__1302 (
            .O(N__14698),
            .I(N__14695));
    LocalMux I__1301 (
            .O(N__14695),
            .I(N__14692));
    Odrv4 I__1300 (
            .O(N__14692),
            .I(\b2v_inst200.un25_clk_100khz_9 ));
    InMux I__1299 (
            .O(N__14689),
            .I(N__14686));
    LocalMux I__1298 (
            .O(N__14686),
            .I(\b2v_inst200.count_2_12 ));
    InMux I__1297 (
            .O(N__14683),
            .I(N__14680));
    LocalMux I__1296 (
            .O(N__14680),
            .I(\b2v_inst200.count_2_13 ));
    CascadeMux I__1295 (
            .O(N__14677),
            .I(\b2v_inst200.countZ0Z_0_cascade_ ));
    InMux I__1294 (
            .O(N__14674),
            .I(N__14671));
    LocalMux I__1293 (
            .O(N__14671),
            .I(\b2v_inst200.un25_clk_100khz_13 ));
    InMux I__1292 (
            .O(N__14668),
            .I(N__14665));
    LocalMux I__1291 (
            .O(N__14665),
            .I(\b2v_inst200.count_2_6 ));
    InMux I__1290 (
            .O(N__14662),
            .I(N__14659));
    LocalMux I__1289 (
            .O(N__14659),
            .I(\b2v_inst200.count_2_14 ));
    InMux I__1288 (
            .O(N__14656),
            .I(N__14653));
    LocalMux I__1287 (
            .O(N__14653),
            .I(N__14650));
    Odrv4 I__1286 (
            .O(N__14650),
            .I(\b2v_inst200.un25_clk_100khz_10 ));
    InMux I__1285 (
            .O(N__14647),
            .I(N__14644));
    LocalMux I__1284 (
            .O(N__14644),
            .I(\b2v_inst200.count_2_3 ));
    InMux I__1283 (
            .O(N__14641),
            .I(N__14638));
    LocalMux I__1282 (
            .O(N__14638),
            .I(\b2v_inst200.count_2_4 ));
    CascadeMux I__1281 (
            .O(N__14635),
            .I(\b2v_inst200.count_RNI_0_0_cascade_ ));
    InMux I__1280 (
            .O(N__14632),
            .I(N__14629));
    LocalMux I__1279 (
            .O(N__14629),
            .I(\b2v_inst200.count_2_11 ));
    InMux I__1278 (
            .O(N__14626),
            .I(N__14623));
    LocalMux I__1277 (
            .O(N__14623),
            .I(\b2v_inst200.count_2_10 ));
    InMux I__1276 (
            .O(N__14620),
            .I(N__14617));
    LocalMux I__1275 (
            .O(N__14617),
            .I(\b2v_inst200.count_2_8 ));
    InMux I__1274 (
            .O(N__14614),
            .I(N__14611));
    LocalMux I__1273 (
            .O(N__14611),
            .I(\b2v_inst200.count_2_0 ));
    InMux I__1272 (
            .O(N__14608),
            .I(N__14602));
    InMux I__1271 (
            .O(N__14607),
            .I(N__14602));
    LocalMux I__1270 (
            .O(N__14602),
            .I(\b2v_inst16.count_rst_1 ));
    InMux I__1269 (
            .O(N__14599),
            .I(N__14596));
    LocalMux I__1268 (
            .O(N__14596),
            .I(\b2v_inst16.count_4_12 ));
    InMux I__1267 (
            .O(N__14593),
            .I(N__14587));
    InMux I__1266 (
            .O(N__14592),
            .I(N__14587));
    LocalMux I__1265 (
            .O(N__14587),
            .I(\b2v_inst16.count_rst_0 ));
    InMux I__1264 (
            .O(N__14584),
            .I(N__14581));
    LocalMux I__1263 (
            .O(N__14581),
            .I(\b2v_inst16.count_4_11 ));
    InMux I__1262 (
            .O(N__14578),
            .I(N__14572));
    InMux I__1261 (
            .O(N__14577),
            .I(N__14572));
    LocalMux I__1260 (
            .O(N__14572),
            .I(N__14569));
    Odrv4 I__1259 (
            .O(N__14569),
            .I(\b2v_inst16.count_rst_11 ));
    InMux I__1258 (
            .O(N__14566),
            .I(N__14563));
    LocalMux I__1257 (
            .O(N__14563),
            .I(\b2v_inst16.count_4_6 ));
    CascadeMux I__1256 (
            .O(N__14560),
            .I(\b2v_inst200.un25_clk_100khz_12_cascade_ ));
    CascadeMux I__1255 (
            .O(N__14557),
            .I(\b2v_inst200.count_RNIC03N_3Z0Z_0_cascade_ ));
    InMux I__1254 (
            .O(N__14554),
            .I(\b2v_inst16.un4_count_1_cry_9 ));
    InMux I__1253 (
            .O(N__14551),
            .I(\b2v_inst16.un4_count_1_cry_10_cZ0 ));
    InMux I__1252 (
            .O(N__14548),
            .I(\b2v_inst16.un4_count_1_cry_11 ));
    InMux I__1251 (
            .O(N__14545),
            .I(\b2v_inst16.un4_count_1_cry_12 ));
    InMux I__1250 (
            .O(N__14542),
            .I(\b2v_inst16.un4_count_1_cry_13 ));
    InMux I__1249 (
            .O(N__14539),
            .I(\b2v_inst16.un4_count_1_cry_14 ));
    InMux I__1248 (
            .O(N__14536),
            .I(N__14530));
    InMux I__1247 (
            .O(N__14535),
            .I(N__14530));
    LocalMux I__1246 (
            .O(N__14530),
            .I(N__14527));
    Odrv4 I__1245 (
            .O(N__14527),
            .I(\b2v_inst16.count_rst_7 ));
    InMux I__1244 (
            .O(N__14524),
            .I(N__14521));
    LocalMux I__1243 (
            .O(N__14521),
            .I(\b2v_inst16.count_4_2 ));
    InMux I__1242 (
            .O(N__14518),
            .I(\b2v_inst16.un4_count_1_cry_1 ));
    InMux I__1241 (
            .O(N__14515),
            .I(N__14511));
    InMux I__1240 (
            .O(N__14514),
            .I(N__14508));
    LocalMux I__1239 (
            .O(N__14511),
            .I(\b2v_inst16.countZ0Z_3 ));
    LocalMux I__1238 (
            .O(N__14508),
            .I(\b2v_inst16.countZ0Z_3 ));
    InMux I__1237 (
            .O(N__14503),
            .I(N__14497));
    InMux I__1236 (
            .O(N__14502),
            .I(N__14497));
    LocalMux I__1235 (
            .O(N__14497),
            .I(\b2v_inst16.count_rst_8 ));
    InMux I__1234 (
            .O(N__14494),
            .I(\b2v_inst16.un4_count_1_cry_2_cZ0 ));
    InMux I__1233 (
            .O(N__14491),
            .I(N__14487));
    InMux I__1232 (
            .O(N__14490),
            .I(N__14484));
    LocalMux I__1231 (
            .O(N__14487),
            .I(\b2v_inst16.countZ0Z_4 ));
    LocalMux I__1230 (
            .O(N__14484),
            .I(\b2v_inst16.countZ0Z_4 ));
    InMux I__1229 (
            .O(N__14479),
            .I(\b2v_inst16.un4_count_1_cry_3 ));
    CascadeMux I__1228 (
            .O(N__14476),
            .I(N__14473));
    InMux I__1227 (
            .O(N__14473),
            .I(N__14469));
    InMux I__1226 (
            .O(N__14472),
            .I(N__14466));
    LocalMux I__1225 (
            .O(N__14469),
            .I(\b2v_inst16.countZ0Z_5 ));
    LocalMux I__1224 (
            .O(N__14466),
            .I(\b2v_inst16.countZ0Z_5 ));
    InMux I__1223 (
            .O(N__14461),
            .I(N__14455));
    InMux I__1222 (
            .O(N__14460),
            .I(N__14455));
    LocalMux I__1221 (
            .O(N__14455),
            .I(\b2v_inst16.count_rst_10 ));
    InMux I__1220 (
            .O(N__14452),
            .I(\b2v_inst16.un4_count_1_cry_4 ));
    InMux I__1219 (
            .O(N__14449),
            .I(\b2v_inst16.un4_count_1_cry_5 ));
    InMux I__1218 (
            .O(N__14446),
            .I(N__14442));
    InMux I__1217 (
            .O(N__14445),
            .I(N__14439));
    LocalMux I__1216 (
            .O(N__14442),
            .I(\b2v_inst16.countZ0Z_7 ));
    LocalMux I__1215 (
            .O(N__14439),
            .I(\b2v_inst16.countZ0Z_7 ));
    InMux I__1214 (
            .O(N__14434),
            .I(\b2v_inst16.un4_count_1_cry_6 ));
    InMux I__1213 (
            .O(N__14431),
            .I(\b2v_inst16.un4_count_1_cry_7 ));
    InMux I__1212 (
            .O(N__14428),
            .I(bfn_1_3_0_));
    InMux I__1211 (
            .O(N__14425),
            .I(N__14422));
    LocalMux I__1210 (
            .O(N__14422),
            .I(\b2v_inst16.count_4_3 ));
    InMux I__1209 (
            .O(N__14419),
            .I(N__14416));
    LocalMux I__1208 (
            .O(N__14416),
            .I(\b2v_inst16.count_4_5 ));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\b2v_inst6.un2_count_1_cry_8 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(\b2v_inst5.un2_count_1_cry_8 ),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_9_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_1_0_));
    defparam IN_MUX_bfv_9_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_2_0_ (
            .carryinitin(\b2v_inst36.un2_count_1_cry_8 ),
            .carryinitout(bfn_9_2_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(b2v_inst20_un4_counter_7),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\b2v_inst20.counter_1_cry_8 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\b2v_inst20.counter_1_cry_16 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(\b2v_inst20.counter_1_cry_24 ),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_1_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_2_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(\b2v_inst16.un4_count_1_cry_8 ),
            .carryinitout(bfn_1_3_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\b2v_inst11.un3_count_off_1_cry_8 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_4_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_1_0_));
    defparam IN_MUX_bfv_4_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_2_0_));
    defparam IN_MUX_bfv_4_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_3_0_));
    defparam IN_MUX_bfv_4_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_4_0_));
    defparam IN_MUX_bfv_5_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_4_0_));
    defparam IN_MUX_bfv_5_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_5_0_));
    defparam IN_MUX_bfv_5_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_6_0_));
    defparam IN_MUX_bfv_4_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_6_0_));
    defparam IN_MUX_bfv_9_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_4_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_7_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_2_0_));
    defparam IN_MUX_bfv_7_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_3_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_6_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_2_0_));
    defparam IN_MUX_bfv_6_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_1_0_));
    defparam IN_MUX_bfv_5_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_1_0_));
    defparam IN_MUX_bfv_5_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_2_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(\b2v_inst11.un1_count_cry_8 ),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(\b2v_inst11.un1_count_clk_2_cry_8_cZ0 ),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_2_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_6_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(\b2v_inst200.un2_count_1_cry_7 ),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(\b2v_inst200.un2_count_1_cry_15 ),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_7_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_5_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(\b2v_inst11.un85_clk_100khz_cry_7 ),
            .carryinitout(bfn_7_6_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(\b2v_inst11.un85_clk_100khz_cry_15_cZ0 ),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_6_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_13_0_));
    defparam IN_MUX_bfv_6_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_14_0_ (
            .carryinitin(\b2v_inst11.un1_dutycycle_94_cry_7_cZ0 ),
            .carryinitout(bfn_6_14_0_));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(\b2v_inst11.un1_dutycycle_53_cry_7_cZ0 ),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(\b2v_inst11.un1_dutycycle_53_cry_15 ),
            .carryinitout(bfn_5_9_0_));
    ICE_GB \b2v_inst200.count_en_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__17362),
            .GLOBALBUFFEROUTPUT(\b2v_inst200.count_en_g ));
    ICE_GB \b2v_inst16.delayed_vddq_pwrgd_en_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__27625),
            .GLOBALBUFFEROUTPUT(b2v_inst16_delayed_vddq_pwrgd_en_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \b2v_inst16.count_RNI_3_LC_1_1_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_3_LC_1_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_3_LC_1_1_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst16.count_RNI_3_LC_1_1_0  (
            .in0(N__14491),
            .in1(N__14446),
            .in2(N__14476),
            .in3(N__14515),
            .lcout(\b2v_inst16.un13_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIF7UJ1_3_LC_1_1_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIF7UJ1_3_LC_1_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIF7UJ1_3_LC_1_1_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNIF7UJ1_3_LC_1_1_1  (
            .in0(N__14425),
            .in1(N__14502),
            .in2(_gnd_net_),
            .in3(N__30624),
            .lcout(\b2v_inst16.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_3_LC_1_1_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_3_LC_1_1_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_3_LC_1_1_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_3_LC_1_1_2  (
            .in0(N__14503),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34638),
            .ce(N__30629),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIHAVJ1_4_LC_1_1_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIHAVJ1_4_LC_1_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIHAVJ1_4_LC_1_1_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNIHAVJ1_4_LC_1_1_3  (
            .in0(N__15259),
            .in1(N__15270),
            .in2(_gnd_net_),
            .in3(N__30625),
            .lcout(\b2v_inst16.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIJD0K1_5_LC_1_1_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIJD0K1_5_LC_1_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIJD0K1_5_LC_1_1_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNIJD0K1_5_LC_1_1_5  (
            .in0(N__14419),
            .in1(N__14460),
            .in2(_gnd_net_),
            .in3(N__30626),
            .lcout(\b2v_inst16.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_5_LC_1_1_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_5_LC_1_1_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_5_LC_1_1_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_5_LC_1_1_6  (
            .in0(N__14461),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34638),
            .ce(N__30629),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNINJ2K1_7_LC_1_1_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNINJ2K1_7_LC_1_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNINJ2K1_7_LC_1_1_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNINJ2K1_7_LC_1_1_7  (
            .in0(N__15277),
            .in1(N__15288),
            .in2(_gnd_net_),
            .in3(N__30627),
            .lcout(\b2v_inst16.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_1_c_LC_1_2_0 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_1_c_LC_1_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_1_c_LC_1_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_1_c_LC_1_2_0  (
            .in0(_gnd_net_),
            .in1(N__15380),
            .in2(N__15226),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_2_0_),
            .carryout(\b2v_inst16.un4_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_1_2_1 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_1_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_1_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_1_2_1  (
            .in0(_gnd_net_),
            .in1(N__15192),
            .in2(_gnd_net_),
            .in3(N__14518),
            .lcout(\b2v_inst16.count_rst_7 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_1 ),
            .carryout(\b2v_inst16.un4_count_1_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_2_2 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_2_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_2_2  (
            .in0(N__20340),
            .in1(N__14514),
            .in2(_gnd_net_),
            .in3(N__14494),
            .lcout(\b2v_inst16.count_rst_8 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_2_cZ0 ),
            .carryout(\b2v_inst16.un4_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_1_2_3 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_1_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_1_2_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_1_2_3  (
            .in0(N__20343),
            .in1(N__14490),
            .in2(_gnd_net_),
            .in3(N__14479),
            .lcout(\b2v_inst16.count_rst_9 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_3 ),
            .carryout(\b2v_inst16.un4_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_1_2_4 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_1_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_1_2_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_1_2_4  (
            .in0(N__20341),
            .in1(N__14472),
            .in2(_gnd_net_),
            .in3(N__14452),
            .lcout(\b2v_inst16.count_rst_10 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_4 ),
            .carryout(\b2v_inst16.un4_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_1_2_5 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_1_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_1_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_1_2_5  (
            .in0(_gnd_net_),
            .in1(N__15171),
            .in2(_gnd_net_),
            .in3(N__14449),
            .lcout(\b2v_inst16.count_rst_11 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_5 ),
            .carryout(\b2v_inst16.un4_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_2_6 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_2_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_2_6  (
            .in0(N__20342),
            .in1(N__14445),
            .in2(_gnd_net_),
            .in3(N__14434),
            .lcout(\b2v_inst16.count_rst_12 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_6 ),
            .carryout(\b2v_inst16.un4_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_1_2_7 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_1_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_1_2_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_1_2_7  (
            .in0(N__20344),
            .in1(N__30198),
            .in2(_gnd_net_),
            .in3(N__14431),
            .lcout(\b2v_inst16.count_rst_13 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_7 ),
            .carryout(\b2v_inst16.un4_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_3_0 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_3_0 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_3_0  (
            .in0(N__20346),
            .in1(_gnd_net_),
            .in2(N__30150),
            .in3(N__14428),
            .lcout(\b2v_inst16.count_rst_14 ),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(\b2v_inst16.un4_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_1_3_1 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_1_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_1_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_1_3_1  (
            .in0(_gnd_net_),
            .in1(N__17319),
            .in2(_gnd_net_),
            .in3(N__14554),
            .lcout(\b2v_inst16.count_rst ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_9 ),
            .carryout(\b2v_inst16.un4_count_1_cry_10_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_10_c_RNIDGU31_LC_1_3_2 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_10_c_RNIDGU31_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_10_c_RNIDGU31_LC_1_3_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_10_c_RNIDGU31_LC_1_3_2  (
            .in0(N__20345),
            .in1(N__15240),
            .in2(_gnd_net_),
            .in3(N__14551),
            .lcout(\b2v_inst16.count_rst_0 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_10_cZ0 ),
            .carryout(\b2v_inst16.un4_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_1_3_3 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_1_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst16.un4_count_1_cry_11_c_RNIRRL3_LC_1_3_3  (
            .in0(_gnd_net_),
            .in1(N__15150),
            .in2(_gnd_net_),
            .in3(N__14548),
            .lcout(\b2v_inst16.count_rst_1 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_11 ),
            .carryout(\b2v_inst16.un4_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_1_3_4 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_1_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_1_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_1_3_4  (
            .in0(_gnd_net_),
            .in1(N__15388),
            .in2(_gnd_net_),
            .in3(N__14545),
            .lcout(\b2v_inst16.count_rst_2 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_12 ),
            .carryout(\b2v_inst16.un4_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_1_3_5 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_1_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_1_3_5  (
            .in0(_gnd_net_),
            .in1(N__15300),
            .in2(_gnd_net_),
            .in3(N__14542),
            .lcout(\b2v_inst16.count_rst_3 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_13 ),
            .carryout(\b2v_inst16.un4_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_1_3_6 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_1_3_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_1_3_6  (
            .in0(N__15346),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14539),
            .lcout(\b2v_inst16.count_rst_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_14_LC_1_3_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_14_LC_1_3_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_14_LC_1_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_14_LC_1_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15313),
            .lcout(\b2v_inst16.count_4_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34626),
            .ce(N__30622),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNID4TJ1_2_LC_1_4_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNID4TJ1_2_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNID4TJ1_2_LC_1_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNID4TJ1_2_LC_1_4_0  (
            .in0(N__14524),
            .in1(N__14535),
            .in2(_gnd_net_),
            .in3(N__30630),
            .lcout(\b2v_inst16.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_2_LC_1_4_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_2_LC_1_4_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_2_LC_1_4_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_2_LC_1_4_1  (
            .in0(N__14536),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34622),
            .ce(N__30628),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIFJV31_12_LC_1_4_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIFJV31_12_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIFJV31_12_LC_1_4_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNIFJV31_12_LC_1_4_2  (
            .in0(N__14599),
            .in1(N__14607),
            .in2(_gnd_net_),
            .in3(N__30633),
            .lcout(\b2v_inst16.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_12_LC_1_4_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_12_LC_1_4_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_12_LC_1_4_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_12_LC_1_4_3  (
            .in0(N__14608),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34622),
            .ce(N__30628),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIJM901_11_LC_1_4_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIJM901_11_LC_1_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIJM901_11_LC_1_4_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNIJM901_11_LC_1_4_4  (
            .in0(N__14584),
            .in1(N__14592),
            .in2(_gnd_net_),
            .in3(N__30632),
            .lcout(\b2v_inst16.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_11_LC_1_4_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_11_LC_1_4_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_11_LC_1_4_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_11_LC_1_4_5  (
            .in0(N__14593),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34622),
            .ce(N__30628),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNILG1K1_6_LC_1_4_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNILG1K1_6_LC_1_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNILG1K1_6_LC_1_4_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst16.count_RNILG1K1_6_LC_1_4_6  (
            .in0(N__14577),
            .in1(N__14566),
            .in2(_gnd_net_),
            .in3(N__30631),
            .lcout(\b2v_inst16.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_6_LC_1_4_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_6_LC_1_4_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_6_LC_1_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_6_LC_1_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14578),
            .lcout(\b2v_inst16.count_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34622),
            .ce(N__30628),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_6_LC_1_5_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_6_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_6_LC_1_5_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst200.count_RNI_6_LC_1_5_0  (
            .in0(N__15948),
            .in1(N__15843),
            .in2(N__15813),
            .in3(N__15891),
            .lcout(),
            .ltout(\b2v_inst200.un25_clk_100khz_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIC03N_3_0_LC_1_5_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIC03N_3_0_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIC03N_3_0_LC_1_5_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst200.count_RNIC03N_3_0_LC_1_5_1  (
            .in0(N__14656),
            .in1(N__14674),
            .in2(N__14560),
            .in3(N__15433),
            .lcout(\b2v_inst200.count_RNIC03N_3Z0Z_0 ),
            .ltout(\b2v_inst200.count_RNIC03N_3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_0_LC_1_5_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_0_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_0_LC_1_5_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst200.count_RNI_0_LC_1_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14557),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_RNI_0_0 ),
            .ltout(\b2v_inst200.count_RNI_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI96451_6_LC_1_5_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI96451_6_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI96451_6_LC_1_5_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \b2v_inst200.count_RNI96451_6_LC_1_5_3  (
            .in0(N__14668),
            .in1(N__15937),
            .in2(N__14635),
            .in3(N__15719),
            .lcout(\b2v_inst200.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI1QM71_11_LC_1_5_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI1QM71_11_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI1QM71_11_LC_1_5_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \b2v_inst200.count_RNI1QM71_11_LC_1_5_4  (
            .in0(N__15796),
            .in1(N__14632),
            .in2(N__33604),
            .in3(N__15721),
            .lcout(\b2v_inst200.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_11_LC_1_5_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_11_LC_1_5_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_11_LC_1_5_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst200.count_11_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(N__15795),
            .in2(_gnd_net_),
            .in3(N__33591),
            .lcout(\b2v_inst200.count_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34617),
            .ce(N__15659),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_10_LC_1_5_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_10_LC_1_5_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_10_LC_1_5_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst200.count_10_LC_1_5_6  (
            .in0(N__33590),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15828),
            .lcout(\b2v_inst200.count_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34617),
            .ce(N__15659),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIOMPC1_10_LC_1_5_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIOMPC1_10_LC_1_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIOMPC1_10_LC_1_5_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \b2v_inst200.count_RNIOMPC1_10_LC_1_5_7  (
            .in0(N__14626),
            .in1(N__33586),
            .in2(N__15832),
            .in3(N__15720),
            .lcout(\b2v_inst200.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIDC651_8_LC_1_6_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIDC651_8_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIDC651_8_LC_1_6_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \b2v_inst200.count_RNIDC651_8_LC_1_6_0  (
            .in0(N__14620),
            .in1(N__33592),
            .in2(N__15880),
            .in3(N__15718),
            .lcout(\b2v_inst200.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_8_LC_1_6_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_8_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_8_LC_1_6_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst200.count_8_LC_1_6_1  (
            .in0(N__33594),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15876),
            .lcout(\b2v_inst200.count_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34615),
            .ce(N__15658),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI73Q71_14_LC_1_6_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI73Q71_14_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI73Q71_14_LC_1_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNI73Q71_14_LC_1_6_2  (
            .in0(N__14662),
            .in1(N__16074),
            .in2(_gnd_net_),
            .in3(N__15716),
            .lcout(\b2v_inst200.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_0_LC_1_6_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_0_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_0_LC_1_6_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst200.count_0_LC_1_6_3  (
            .in0(N__33593),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15607),
            .lcout(\b2v_inst200.count_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34615),
            .ce(N__15658),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIC03N_0_LC_1_6_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIC03N_0_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIC03N_0_LC_1_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNIC03N_0_LC_1_6_4  (
            .in0(N__14614),
            .in1(N__15595),
            .in2(_gnd_net_),
            .in3(N__15717),
            .lcout(\b2v_inst200.countZ0Z_0 ),
            .ltout(\b2v_inst200.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIC03N_1_0_LC_1_6_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIC03N_1_0_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIC03N_1_0_LC_1_6_5 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \b2v_inst200.count_RNIC03N_1_0_LC_1_6_5  (
            .in0(_gnd_net_),
            .in1(N__14698),
            .in2(N__14677),
            .in3(N__16087),
            .lcout(\b2v_inst200.un25_clk_100khz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_6_LC_1_6_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_6_LC_1_6_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_6_LC_1_6_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst200.count_6_LC_1_6_6  (
            .in0(N__15936),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33595),
            .lcout(\b2v_inst200.count_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34615),
            .ce(N__15658),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_14_LC_1_6_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_14_LC_1_6_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_14_LC_1_6_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_14_LC_1_6_7  (
            .in0(N__16075),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34615),
            .ce(N__15658),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_3_LC_1_7_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_3_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_3_LC_1_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst200.count_RNI_3_LC_1_7_0  (
            .in0(N__15481),
            .in1(N__15922),
            .in2(N__15508),
            .in3(N__15532),
            .lcout(\b2v_inst200.un25_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI3T051_3_LC_1_7_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI3T051_3_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI3T051_3_LC_1_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNI3T051_3_LC_1_7_1  (
            .in0(N__14647),
            .in1(N__15519),
            .in2(_gnd_net_),
            .in3(N__15708),
            .lcout(\b2v_inst200.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_3_LC_1_7_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_3_LC_1_7_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_3_LC_1_7_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_3_LC_1_7_2  (
            .in0(N__15520),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34611),
            .ce(N__15657),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI50251_4_LC_1_7_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI50251_4_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI50251_4_LC_1_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst200.count_RNI50251_4_LC_1_7_3  (
            .in0(N__15492),
            .in1(N__14641),
            .in2(_gnd_net_),
            .in3(N__15709),
            .lcout(\b2v_inst200.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_4_LC_1_7_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_4_LC_1_7_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_4_LC_1_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_4_LC_1_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15493),
            .lcout(\b2v_inst200.count_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34611),
            .ce(N__15657),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI73351_5_LC_1_7_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI73351_5_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI73351_5_LC_1_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNI73351_5_LC_1_7_5  (
            .in0(N__14713),
            .in1(N__15468),
            .in2(_gnd_net_),
            .in3(N__15710),
            .lcout(\b2v_inst200.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_5_LC_1_7_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_5_LC_1_7_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_5_LC_1_7_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_5_LC_1_7_6  (
            .in0(N__15469),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34611),
            .ce(N__15657),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIB9551_7_LC_1_7_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIB9551_7_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIB9551_7_LC_1_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNIB9551_7_LC_1_7_7  (
            .in0(N__15445),
            .in1(N__15906),
            .in2(_gnd_net_),
            .in3(N__15711),
            .lcout(\b2v_inst200.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_9_LC_1_8_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_9_LC_1_8_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_9_LC_1_8_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_9_LC_1_8_0  (
            .in0(N__15859),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34609),
            .ce(N__15656),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIFF751_9_LC_1_8_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIFF751_9_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIFF751_9_LC_1_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNIFF751_9_LC_1_8_1  (
            .in0(N__14707),
            .in1(N__15858),
            .in2(_gnd_net_),
            .in3(N__15712),
            .lcout(\b2v_inst200.countZ0Z_9 ),
            .ltout(\b2v_inst200.countZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_9_LC_1_8_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_9_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_9_LC_1_8_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst200.count_RNI_9_LC_1_8_2  (
            .in0(N__15781),
            .in1(N__15757),
            .in2(N__14701),
            .in3(N__16063),
            .lcout(\b2v_inst200.un25_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI3TN71_12_LC_1_8_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI3TN71_12_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI3TN71_12_LC_1_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst200.count_RNI3TN71_12_LC_1_8_3  (
            .in0(N__15768),
            .in1(N__14689),
            .in2(_gnd_net_),
            .in3(N__15713),
            .lcout(\b2v_inst200.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_12_LC_1_8_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_12_LC_1_8_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_12_LC_1_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_12_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15769),
            .lcout(\b2v_inst200.count_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34609),
            .ce(N__15656),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI50P71_13_LC_1_8_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI50P71_13_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI50P71_13_LC_1_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNI50P71_13_LC_1_8_5  (
            .in0(N__14683),
            .in1(N__15744),
            .in2(_gnd_net_),
            .in3(N__15714),
            .lcout(\b2v_inst200.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_13_LC_1_8_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_13_LC_1_8_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_13_LC_1_8_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_13_LC_1_8_6  (
            .in0(N__15745),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34609),
            .ce(N__15656),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI96R71_15_LC_1_8_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI96R71_15_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI96R71_15_LC_1_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNI96R71_15_LC_1_8_7  (
            .in0(N__15457),
            .in1(N__16047),
            .in2(_gnd_net_),
            .in3(N__15715),
            .lcout(\b2v_inst200.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_LC_1_9_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_LC_1_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_1_c_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(N__16430),
            .in2(N__16696),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_1_9_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_1_9_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_1_9_1  (
            .in0(N__16606),
            .in1(N__16270),
            .in2(_gnd_net_),
            .in3(N__14737),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_1 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_1_9_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_1_9_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_1_9_2  (
            .in0(N__16600),
            .in1(N__16253),
            .in2(_gnd_net_),
            .in3(N__14734),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_2 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_1_9_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_1_9_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_1_9_3  (
            .in0(N__16603),
            .in1(_gnd_net_),
            .in2(N__16297),
            .in3(N__14731),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_3 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_1_9_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_1_9_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_1_9_4  (
            .in0(N__16601),
            .in1(_gnd_net_),
            .in2(N__16402),
            .in3(N__14728),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_4 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_1_9_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_1_9_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_1_9_5  (
            .in0(N__16604),
            .in1(_gnd_net_),
            .in2(N__16318),
            .in3(N__14725),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_5 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_1_9_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_1_9_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_1_9_6  (
            .in0(N__16602),
            .in1(_gnd_net_),
            .in2(N__16237),
            .in3(N__14722),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_6 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_1_9_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_1_9_7 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_1_9_7  (
            .in0(N__16605),
            .in1(_gnd_net_),
            .in2(N__16339),
            .in3(N__14719),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_7_cZ0 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_1_10_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_1_10_0 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_1_10_0  (
            .in0(N__16593),
            .in1(_gnd_net_),
            .in2(N__16717),
            .in3(N__14716),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_9_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_1_10_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_1_10_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16192),
            .in3(N__14773),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_9_cZ0 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_10_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_1_10_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_1_10_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16183),
            .in3(N__14770),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AAZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_10_cZ0 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_1_10_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_1_10_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16489),
            .in3(N__14767),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BAZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_11 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_1_10_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_1_10_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_1_10_4  (
            .in0(N__16594),
            .in1(_gnd_net_),
            .in2(N__16117),
            .in3(N__14764),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CAZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_12 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_1_10_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_1_10_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_1_10_5  (
            .in0(N__16618),
            .in1(_gnd_net_),
            .in2(N__16147),
            .in3(N__14761),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DAZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_13 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_1_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_1_10_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_1_10_6  (
            .in0(N__16595),
            .in1(N__16164),
            .in2(_gnd_net_),
            .in3(N__14758),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI0JFF5_5_LC_1_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI0JFF5_5_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI0JFF5_5_LC_1_11_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_clk_RNI0JFF5_5_LC_1_11_0  (
            .in0(N__14743),
            .in1(N__17480),
            .in2(_gnd_net_),
            .in3(N__14754),
            .lcout(\b2v_inst11.count_clkZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_5_LC_1_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_5_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_5_LC_1_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_5_LC_1_11_1  (
            .in0(N__14755),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34610),
            .ce(N__17542),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI281F5_15_LC_1_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI281F5_15_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI281F5_15_LC_1_11_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_clk_RNI281F5_15_LC_1_11_2  (
            .in0(N__14857),
            .in1(N__17483),
            .in2(_gnd_net_),
            .in3(N__14868),
            .lcout(\b2v_inst11.count_clkZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_15_LC_1_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_15_LC_1_11_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_15_LC_1_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_15_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14872),
            .lcout(\b2v_inst11.count_clk_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34610),
            .ce(N__17542),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI2MGF5_6_LC_1_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI2MGF5_6_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI2MGF5_6_LC_1_11_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_clk_RNI2MGF5_6_LC_1_11_4  (
            .in0(N__14839),
            .in1(N__17481),
            .in2(_gnd_net_),
            .in3(N__14850),
            .lcout(\b2v_inst11.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_6_LC_1_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_6_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_6_LC_1_11_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_6_LC_1_11_5  (
            .in0(N__14851),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34610),
            .ce(N__17542),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI6SIF5_8_LC_1_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI6SIF5_8_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI6SIF5_8_LC_1_11_6 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \b2v_inst11.count_clk_RNI6SIF5_8_LC_1_11_6  (
            .in0(N__14818),
            .in1(N__17482),
            .in2(N__14833),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clkZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_8_LC_1_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_8_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_8_LC_1_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_8_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14832),
            .lcout(\b2v_inst11.count_clk_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34610),
            .ce(N__17542),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI4PHF5_7_LC_1_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI4PHF5_7_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI4PHF5_7_LC_1_12_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_clk_RNI4PHF5_7_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__14797),
            .in2(N__14812),
            .in3(N__17524),
            .lcout(\b2v_inst11.count_clkZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_7_LC_1_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_7_LC_1_12_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_7_LC_1_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_7_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14811),
            .lcout(\b2v_inst11.count_clk_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34614),
            .ce(N__17537),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI8VJF5_9_LC_1_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI8VJF5_9_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI8VJF5_9_LC_1_12_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_clk_RNI8VJF5_9_LC_1_12_2  (
            .in0(N__14779),
            .in1(N__17525),
            .in2(_gnd_net_),
            .in3(N__14790),
            .lcout(\b2v_inst11.count_clkZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_9_LC_1_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_9_LC_1_12_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_9_LC_1_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_9_LC_1_12_3  (
            .in0(N__14791),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34614),
            .ce(N__17537),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIUFEF5_4_LC_1_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIUFEF5_4_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIUFEF5_4_LC_1_12_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_clk_RNIUFEF5_4_LC_1_12_4  (
            .in0(N__14896),
            .in1(N__17523),
            .in2(_gnd_net_),
            .in3(N__14907),
            .lcout(\b2v_inst11.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_4_LC_1_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_4_LC_1_12_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_4_LC_1_12_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_4_LC_1_12_5  (
            .in0(N__14908),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34614),
            .ce(N__17537),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNINJ641_7_LC_1_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNINJ641_7_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNINJ641_7_LC_1_12_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst11.count_clk_RNINJ641_7_LC_1_12_6  (
            .in0(N__24328),
            .in1(N__23043),
            .in2(_gnd_net_),
            .in3(N__16641),
            .lcout(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNICG51A_6_LC_1_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNICG51A_6_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNICG51A_6_LC_1_12_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_off_RNICG51A_6_LC_1_12_7  (
            .in0(N__16752),
            .in1(N__18138),
            .in2(_gnd_net_),
            .in3(N__16923),
            .lcout(\b2v_inst11.un3_count_off_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_5_LC_1_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_5_LC_1_13_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_5_LC_1_13_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_5_LC_1_13_0  (
            .in0(N__14935),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19562),
            .lcout(\b2v_inst11.count_off_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34616),
            .ce(N__18153),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI4411A_2_LC_1_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI4411A_2_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI4411A_2_LC_1_13_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_off_RNI4411A_2_LC_1_13_1  (
            .in0(N__14883),
            .in1(N__18130),
            .in2(_gnd_net_),
            .in3(N__14890),
            .lcout(\b2v_inst11.un3_count_off_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_2_LC_1_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_2_LC_1_13_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_2_LC_1_13_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_2_LC_1_13_2  (
            .in0(N__14968),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19561),
            .lcout(\b2v_inst11.count_offZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34616),
            .ce(N__18153),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIIQOD2_LC_1_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIIQOD2_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIIQOD2_LC_1_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_1_c_RNIIQOD2_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__19541),
            .in2(_gnd_net_),
            .in3(N__14967),
            .lcout(\b2v_inst11.count_off_1_2 ),
            .ltout(\b2v_inst11.count_off_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI4411A_0_2_LC_1_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI4411A_0_2_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI4411A_0_2_LC_1_13_4 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \b2v_inst11.count_off_RNI4411A_0_2_LC_1_13_4  (
            .in0(N__18154),
            .in1(N__14884),
            .in2(N__14875),
            .in3(N__14949),
            .lcout(\b2v_inst11.un34_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNICG51A_0_6_LC_1_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNICG51A_0_6_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNICG51A_0_6_LC_1_13_5 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \b2v_inst11.count_off_RNICG51A_0_6_LC_1_13_5  (
            .in0(N__16753),
            .in1(N__17911),
            .in2(N__16930),
            .in3(N__18155),
            .lcout(),
            .ltout(\b2v_inst11.un34_clk_100khz_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI4FF481_2_LC_1_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI4FF481_2_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI4FF481_2_LC_1_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.count_off_RNI4FF481_2_LC_1_13_6  (
            .in0(N__15088),
            .in1(N__17023),
            .in2(N__14989),
            .in3(N__14986),
            .lcout(\b2v_inst11.un34_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIAD41A_5_LC_1_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIAD41A_5_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIAD41A_5_LC_1_13_7 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \b2v_inst11.count_off_RNIAD41A_5_LC_1_13_7  (
            .in0(N__14980),
            .in1(N__18131),
            .in2(N__19581),
            .in3(N__14934),
            .lcout(\b2v_inst11.count_offZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_LC_1_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_LC_1_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_1_c_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__17863),
            .in2(N__17910),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\b2v_inst11.un3_count_off_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_1_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_1_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__14974),
            .in2(_gnd_net_),
            .in3(N__14959),
            .lcout(\b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_1 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_1_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_1_14_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15121),
            .in3(N__14956),
            .lcout(\b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_2_cZ0 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_3_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_1_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_1_14_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15109),
            .in3(N__14953),
            .lcout(\b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_3_cZ0 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_4_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_1_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_1_14_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14950),
            .in3(N__14926),
            .lcout(\b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_4_cZ0 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_1_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_1_14_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14923),
            .in3(N__14911),
            .lcout(\b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_5 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_1_14_6 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_1_14_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16990),
            .in3(N__15016),
            .lcout(\b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_6 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_1_14_7 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_1_14_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17038),
            .in3(N__15013),
            .lcout(\b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_7 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_1_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_1_15_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16948),
            .in3(N__15010),
            .lcout(\b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\b2v_inst11.un3_count_off_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_1_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_1_15_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17800),
            .in3(N__15007),
            .lcout(\b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_9 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_1_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_1_15_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16510),
            .in3(N__15004),
            .lcout(\b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_10 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_1_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_1_15_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16786),
            .in3(N__15001),
            .lcout(\b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_11 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_1_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_1_15_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16870),
            .in3(N__14998),
            .lcout(\b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_12 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_1_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_1_15_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16854),
            .in3(N__14995),
            .lcout(\b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_13 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_1_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_1_15_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_1_15_6  (
            .in0(N__16876),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14992),
            .lcout(\b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI8V45A_13_LC_1_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI8V45A_13_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI8V45A_13_LC_1_15_7 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \b2v_inst11.count_off_RNI8V45A_13_LC_1_15_7  (
            .in0(N__19580),
            .in1(N__18137),
            .in2(N__18175),
            .in3(N__17772),
            .lcout(\b2v_inst11.count_offZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIJSPD2_LC_1_16_0 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIJSPD2_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIJSPD2_LC_1_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_2_c_RNIJSPD2_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__19572),
            .in2(_gnd_net_),
            .in3(N__15078),
            .lcout(\b2v_inst11.count_off_1_3 ),
            .ltout(\b2v_inst11.count_off_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI6721A_3_LC_1_16_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI6721A_3_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI6721A_3_LC_1_16_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_off_RNI6721A_3_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__15066),
            .in2(N__15124),
            .in3(N__18132),
            .lcout(\b2v_inst11.un3_count_off_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI8A31A_4_LC_1_16_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI8A31A_4_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI8A31A_4_LC_1_16_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst11.count_off_RNI8A31A_4_LC_1_16_2  (
            .in0(N__18133),
            .in1(N__19573),
            .in2(N__15046),
            .in3(N__15057),
            .lcout(\b2v_inst11.count_offZ0Z_4 ),
            .ltout(\b2v_inst11.count_offZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI6721A_0_3_LC_1_16_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI6721A_0_3_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI6721A_0_3_LC_1_16_3 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \b2v_inst11.count_off_RNI6721A_0_3_LC_1_16_3  (
            .in0(N__15097),
            .in1(N__15067),
            .in2(N__15091),
            .in3(N__18136),
            .lcout(\b2v_inst11.un34_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_3_LC_1_16_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_3_LC_1_16_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_3_LC_1_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_3_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(N__19575),
            .in2(_gnd_net_),
            .in3(N__15079),
            .lcout(\b2v_inst11.count_offZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34630),
            .ce(N__18135),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_4_LC_1_16_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_4_LC_1_16_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_4_LC_1_16_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \b2v_inst11.count_off_4_LC_1_16_5  (
            .in0(N__15058),
            .in1(_gnd_net_),
            .in2(N__19582),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34630),
            .ce(N__18135),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_14_LC_1_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_14_LC_1_16_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_14_LC_1_16_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.count_off_14_LC_1_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15028),
            .in3(N__19579),
            .lcout(\b2v_inst11.count_off_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34630),
            .ce(N__18135),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIA265A_14_LC_1_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIA265A_14_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIA265A_14_LC_1_16_7 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \b2v_inst11.count_off_RNIA265A_14_LC_1_16_7  (
            .in0(N__19574),
            .in1(N__18134),
            .in2(N__15037),
            .in3(N__15024),
            .lcout(\b2v_inst11.count_offZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_7_LC_2_1_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_7_LC_2_1_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_7_LC_2_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_7_LC_2_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15289),
            .lcout(\b2v_inst16.count_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34647),
            .ce(N__30623),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_4_LC_2_1_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_4_LC_2_1_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_4_LC_2_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_4_LC_2_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15271),
            .lcout(\b2v_inst16.count_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34647),
            .ce(N__30623),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_1_LC_2_2_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_1_LC_2_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_1_LC_2_2_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst16.count_RNI_1_LC_2_2_0  (
            .in0(_gnd_net_),
            .in1(N__15222),
            .in2(_gnd_net_),
            .in3(N__15377),
            .lcout(\b2v_inst16.count_rst_6 ),
            .ltout(\b2v_inst16.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI2J651_0_1_LC_2_2_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI2J651_0_1_LC_2_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI2J651_0_1_LC_2_2_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst16.count_RNI2J651_0_1_LC_2_2_1  (
            .in0(_gnd_net_),
            .in1(N__15204),
            .in2(N__15253),
            .in3(N__30609),
            .lcout(\b2v_inst16.un4_count_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI2J651_1_LC_2_2_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI2J651_1_LC_2_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI2J651_1_LC_2_2_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \b2v_inst16.count_RNI2J651_1_LC_2_2_2  (
            .in0(N__15205),
            .in1(_gnd_net_),
            .in2(N__30643),
            .in3(N__15250),
            .lcout(),
            .ltout(\b2v_inst16.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIL9G52_1_LC_2_2_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIL9G52_1_LC_2_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIL9G52_1_LC_2_2_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst16.count_RNIL9G52_1_LC_2_2_3  (
            .in0(N__15244),
            .in1(N__30199),
            .in2(N__15229),
            .in3(N__30151),
            .lcout(\b2v_inst16.un13_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_1_LC_2_2_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_1_LC_2_2_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_1_LC_2_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst16.count_1_LC_2_2_4  (
            .in0(_gnd_net_),
            .in1(N__15221),
            .in2(_gnd_net_),
            .in3(N__15379),
            .lcout(\b2v_inst16.count_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34640),
            .ce(N__30639),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_10_LC_2_2_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_10_LC_2_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_10_LC_2_2_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst16.count_RNI_10_LC_2_2_5  (
            .in0(N__15196),
            .in1(N__17320),
            .in2(N__15175),
            .in3(N__15154),
            .lcout(),
            .ltout(\b2v_inst16.un13_clk_100khz_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIL9G52_0_1_LC_2_2_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIL9G52_0_1_LC_2_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIL9G52_0_1_LC_2_2_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \b2v_inst16.count_RNIL9G52_0_1_LC_2_2_6  (
            .in0(N__15139),
            .in1(N__15133),
            .in2(N__15127),
            .in3(N__15352),
            .lcout(\b2v_inst16.un13_clk_100khz_i ),
            .ltout(\b2v_inst16.un13_clk_100khz_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_0_LC_2_2_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_0_LC_2_2_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_0_LC_2_2_7 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \b2v_inst16.count_0_LC_2_2_7  (
            .in0(N__15378),
            .in1(_gnd_net_),
            .in2(N__15415),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34640),
            .ce(N__30639),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_13_LC_2_3_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_13_LC_2_3_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_13_LC_2_3_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_13_LC_2_3_0  (
            .in0(N__15397),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34632),
            .ce(N__30598),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_0_LC_2_3_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_0_LC_2_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_0_LC_2_3_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst16.count_RNI_0_LC_2_3_1  (
            .in0(N__20339),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15382),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI1I651_0_LC_2_3_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI1I651_0_LC_2_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI1I651_0_LC_2_3_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst16.count_RNI1I651_0_LC_2_3_2  (
            .in0(_gnd_net_),
            .in1(N__15412),
            .in2(N__15406),
            .in3(N__30571),
            .lcout(\b2v_inst16.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIHM041_13_LC_2_3_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIHM041_13_LC_2_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIHM041_13_LC_2_3_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst16.count_RNIHM041_13_LC_2_3_3  (
            .in0(N__30572),
            .in1(N__15403),
            .in2(_gnd_net_),
            .in3(N__15396),
            .lcout(\b2v_inst16.countZ0Z_13 ),
            .ltout(\b2v_inst16.countZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_15_LC_2_3_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_15_LC_2_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_15_LC_2_3_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst16.count_RNI_15_LC_2_3_4  (
            .in0(N__15381),
            .in1(N__15301),
            .in2(N__15355),
            .in3(N__15345),
            .lcout(\b2v_inst16.un13_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNILS241_15_LC_2_3_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNILS241_15_LC_2_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNILS241_15_LC_2_3_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst16.count_RNILS241_15_LC_2_3_5  (
            .in0(N__30574),
            .in1(N__15325),
            .in2(_gnd_net_),
            .in3(N__15333),
            .lcout(\b2v_inst16.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_15_LC_2_3_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_15_LC_2_3_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_15_LC_2_3_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_15_LC_2_3_6  (
            .in0(N__15334),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34632),
            .ce(N__30598),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIJP141_14_LC_2_3_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIJP141_14_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIJP141_14_LC_2_3_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst16.count_RNIJP141_14_LC_2_3_7  (
            .in0(N__30573),
            .in1(N__15319),
            .in2(_gnd_net_),
            .in3(N__15312),
            .lcout(\b2v_inst16.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_15_LC_2_4_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_15_LC_2_4_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_15_LC_2_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_15_LC_2_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16051),
            .lcout(\b2v_inst200.count_2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34628),
            .ce(N__15661),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_2_LC_2_4_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_2_LC_2_4_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_2_LC_2_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_2_LC_2_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15550),
            .lcout(\b2v_inst200.count_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34628),
            .ce(N__15661),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_7_LC_2_4_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_7_LC_2_4_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_7_LC_2_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_7_LC_2_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15910),
            .lcout(\b2v_inst200.count_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34628),
            .ce(N__15661),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_17_LC_2_5_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_17_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_17_LC_2_5_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \b2v_inst200.count_RNI_17_LC_2_5_0  (
            .in0(N__16026),
            .in1(N__15562),
            .in2(N__15589),
            .in3(N__15996),
            .lcout(\b2v_inst200.un25_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIB9S71_16_LC_2_5_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIB9S71_16_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIB9S71_16_LC_2_5_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNIB9S71_16_LC_2_5_1  (
            .in0(N__15427),
            .in1(N__16015),
            .in2(_gnd_net_),
            .in3(N__15707),
            .lcout(\b2v_inst200.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_16_LC_2_5_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_16_LC_2_5_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_16_LC_2_5_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_16_LC_2_5_2  (
            .in0(N__16014),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34623),
            .ce(N__15660),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIDCT71_17_LC_2_5_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIDCT71_17_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIDCT71_17_LC_2_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNIDCT71_17_LC_2_5_3  (
            .in0(N__15421),
            .in1(N__15981),
            .in2(_gnd_net_),
            .in3(N__15705),
            .lcout(\b2v_inst200.countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_17_LC_2_5_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_17_LC_2_5_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_17_LC_2_5_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_17_LC_2_5_4  (
            .in0(N__15982),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34623),
            .ce(N__15660),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIP16E1_1_LC_2_5_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIP16E1_1_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIP16E1_1_LC_2_5_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNIP16E1_1_LC_2_5_5  (
            .in0(N__15733),
            .in1(N__15573),
            .in2(_gnd_net_),
            .in3(N__15706),
            .lcout(\b2v_inst200.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_1_LC_2_5_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_1_LC_2_5_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_1_LC_2_5_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_1_LC_2_5_6  (
            .in0(N__15574),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34623),
            .ce(N__15660),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI1QV41_2_LC_2_5_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI1QV41_2_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI1QV41_2_LC_2_5_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNI1QV41_2_LC_2_5_7  (
            .in0(N__15727),
            .in1(N__15549),
            .in2(_gnd_net_),
            .in3(N__15704),
            .lcout(\b2v_inst200.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIC03N_0_0_LC_2_6_0 .C_ON=1'b1;
    defparam \b2v_inst200.count_RNIC03N_0_0_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIC03N_0_0_LC_2_6_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst200.count_RNIC03N_0_0_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(N__15606),
            .in2(_gnd_net_),
            .in3(N__33585),
            .lcout(\b2v_inst200.count_1_0 ),
            .ltout(),
            .carryin(bfn_2_6_0_),
            .carryout(\b2v_inst200.un2_count_1_cry_1_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIC03N_5_0_LC_2_6_1 .C_ON=1'b1;
    defparam \b2v_inst200.count_RNIC03N_5_0_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIC03N_5_0_LC_2_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.count_RNIC03N_5_0_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(N__15585),
            .in2(_gnd_net_),
            .in3(N__15565),
            .lcout(\b2v_inst200.count_RNIC03N_5Z0Z_0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_1_cy ),
            .carryout(\b2v_inst200.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_2_6_2 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_2_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_2_6_2  (
            .in0(_gnd_net_),
            .in1(N__15561),
            .in2(_gnd_net_),
            .in3(N__15535),
            .lcout(\b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_1 ),
            .carryout(\b2v_inst200.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_2_6_3 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_2_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_2_6_3  (
            .in0(_gnd_net_),
            .in1(N__15531),
            .in2(_gnd_net_),
            .in3(N__15511),
            .lcout(\b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_2 ),
            .carryout(\b2v_inst200.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_2_6_4 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_2_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_2_6_4  (
            .in0(_gnd_net_),
            .in1(N__15504),
            .in2(_gnd_net_),
            .in3(N__15484),
            .lcout(\b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_3 ),
            .carryout(\b2v_inst200.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_2_6_5 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_2_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_2_6_5  (
            .in0(_gnd_net_),
            .in1(N__15480),
            .in2(_gnd_net_),
            .in3(N__15460),
            .lcout(\b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_4 ),
            .carryout(\b2v_inst200.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_2_6_6 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_2_6_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_2_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15952),
            .in3(N__15925),
            .lcout(\b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_5 ),
            .carryout(\b2v_inst200.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_2_6_7 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_2_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_2_6_7  (
            .in0(_gnd_net_),
            .in1(N__15921),
            .in2(_gnd_net_),
            .in3(N__15895),
            .lcout(\b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_6 ),
            .carryout(\b2v_inst200.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_2_7_0 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_2_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_2_7_0  (
            .in0(_gnd_net_),
            .in1(N__15892),
            .in2(_gnd_net_),
            .in3(N__15868),
            .lcout(\b2v_inst200.un2_count_1_cry_7_c_RNIP33EZ0 ),
            .ltout(),
            .carryin(bfn_2_7_0_),
            .carryout(\b2v_inst200.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_2_7_1 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_2_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(N__15865),
            .in2(_gnd_net_),
            .in3(N__15850),
            .lcout(\b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_8 ),
            .carryout(\b2v_inst200.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_2_7_2 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_2_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(N__15847),
            .in2(_gnd_net_),
            .in3(N__15817),
            .lcout(\b2v_inst200.un2_count_1_cry_9_c_RNIR75EZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_9 ),
            .carryout(\b2v_inst200.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_2_7_3 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_2_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_2_7_3  (
            .in0(_gnd_net_),
            .in1(N__15814),
            .in2(_gnd_net_),
            .in3(N__15784),
            .lcout(\b2v_inst200.un2_count_1_cry_10_c_RNI3AZ0Z29 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_10 ),
            .carryout(\b2v_inst200.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_2_7_4 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_2_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_2_7_4  (
            .in0(_gnd_net_),
            .in1(N__15780),
            .in2(_gnd_net_),
            .in3(N__15760),
            .lcout(\b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_11 ),
            .carryout(\b2v_inst200.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_2_7_5 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_2_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_2_7_5  (
            .in0(_gnd_net_),
            .in1(N__15756),
            .in2(_gnd_net_),
            .in3(N__15736),
            .lcout(\b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_12 ),
            .carryout(\b2v_inst200.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_2_7_6 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_2_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_2_7_6  (
            .in0(_gnd_net_),
            .in1(N__16086),
            .in2(_gnd_net_),
            .in3(N__16066),
            .lcout(\b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_13 ),
            .carryout(\b2v_inst200.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_14_c_RNI7I69_LC_2_7_7 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_14_c_RNI7I69_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_14_c_RNI7I69_LC_2_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_14_c_RNI7I69_LC_2_7_7  (
            .in0(_gnd_net_),
            .in1(N__16062),
            .in2(_gnd_net_),
            .in3(N__16036),
            .lcout(\b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_14 ),
            .carryout(\b2v_inst200.un2_count_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_2_8_0 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_2_8_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_2_8_0  (
            .in0(N__33608),
            .in1(N__16033),
            .in2(_gnd_net_),
            .in3(N__16003),
            .lcout(\b2v_inst200.count_1_16 ),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(\b2v_inst200.un2_count_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_2_8_1 .C_ON=1'b0;
    defparam \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_2_8_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_2_8_1  (
            .in0(N__16000),
            .in1(N__33609),
            .in2(_gnd_net_),
            .in3(N__15985),
            .lcout(\b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIQRSE5_11_LC_2_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIQRSE5_11_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIQRSE5_11_LC_2_9_0 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \b2v_inst11.count_clk_RNIQRSE5_11_LC_2_9_0  (
            .in0(N__15961),
            .in1(N__16610),
            .in2(N__17499),
            .in3(N__15969),
            .lcout(\b2v_inst11.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_10_LC_2_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_10_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_10_LC_2_9_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \b2v_inst11.count_clk_10_LC_2_9_1  (
            .in0(N__16613),
            .in1(N__16201),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34608),
            .ce(N__17511),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_11_LC_2_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_11_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_11_LC_2_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_clk_11_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(N__16612),
            .in2(_gnd_net_),
            .in3(N__15970),
            .lcout(\b2v_inst11.count_clk_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34608),
            .ce(N__17511),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIS1M95_0_LC_2_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIS1M95_0_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIS1M95_0_LC_2_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_clk_RNIS1M95_0_LC_2_9_3  (
            .in0(N__16450),
            .in1(N__16213),
            .in2(_gnd_net_),
            .in3(N__17466),
            .lcout(\b2v_inst11.count_clkZ0Z_0 ),
            .ltout(\b2v_inst11.count_clkZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_0_LC_2_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_0_LC_2_9_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_0_LC_2_9_4 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \b2v_inst11.count_clk_0_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15955),
            .in3(N__16611),
            .lcout(\b2v_inst11.count_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34608),
            .ce(N__17511),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIHFHA5_10_LC_2_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIHFHA5_10_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIHFHA5_10_LC_2_9_5 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \b2v_inst11.count_clk_RNIHFHA5_10_LC_2_9_5  (
            .in0(N__16207),
            .in1(N__17467),
            .in2(N__16617),
            .in3(N__16200),
            .lcout(\b2v_inst11.count_clkZ0Z_10 ),
            .ltout(\b2v_inst11.count_clkZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_15_LC_2_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_15_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_15_LC_2_9_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst11.count_clk_RNI_15_LC_2_9_6  (
            .in0(N__16488),
            .in1(N__16182),
            .in2(N__16168),
            .in3(N__16165),
            .lcout(),
            .ltout(\b2v_inst11.un2_count_clk_17_0_o2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_13_LC_2_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_13_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_13_LC_2_9_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst11.count_clk_RNI_13_LC_2_9_7  (
            .in0(N__16431),
            .in1(N__16146),
            .in2(N__16150),
            .in3(N__16116),
            .lcout(\b2v_inst11.N_172 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI050F5_14_LC_2_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI050F5_14_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI050F5_14_LC_2_10_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_clk_RNI050F5_14_LC_2_10_0  (
            .in0(N__17485),
            .in1(N__16093),
            .in2(_gnd_net_),
            .in3(N__16101),
            .lcout(\b2v_inst11.count_clkZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_13_LC_2_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_13_LC_2_10_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_13_LC_2_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_13_LC_2_10_1  (
            .in0(N__16126),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34612),
            .ce(N__17527),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIU1VE5_13_LC_2_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIU1VE5_13_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIU1VE5_13_LC_2_10_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_clk_RNIU1VE5_13_LC_2_10_2  (
            .in0(N__17484),
            .in1(N__16132),
            .in2(_gnd_net_),
            .in3(N__16125),
            .lcout(\b2v_inst11.count_clkZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_14_LC_2_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_14_LC_2_10_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_14_LC_2_10_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_14_LC_2_10_3  (
            .in0(N__16102),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34612),
            .ce(N__17527),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIR4RV4_1_LC_2_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIR4RV4_1_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIR4RV4_1_LC_2_10_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst11.func_state_RNIR4RV4_1_LC_2_10_4  (
            .in0(N__22846),
            .in1(N__27587),
            .in2(N__16498),
            .in3(N__17929),
            .lcout(\b2v_inst11.count_clk_en ),
            .ltout(\b2v_inst11.count_clk_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIQ9CF5_2_LC_2_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIQ9CF5_2_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIQ9CF5_2_LC_2_10_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \b2v_inst11.count_clk_RNIQ9CF5_2_LC_2_10_5  (
            .in0(N__16366),
            .in1(_gnd_net_),
            .in2(N__16369),
            .in3(N__16357),
            .lcout(\b2v_inst11.count_clkZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_2_LC_2_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_2_LC_2_10_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_2_LC_2_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_2_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16365),
            .lcout(\b2v_inst11.count_clk_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34612),
            .ce(N__17527),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNISCDF5_3_LC_2_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNISCDF5_3_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNISCDF5_3_LC_2_10_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \b2v_inst11.count_clk_RNISCDF5_3_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(N__17554),
            .in2(N__17500),
            .in3(N__17565),
            .lcout(\b2v_inst11.count_clkZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_7_LC_2_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_7_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_7_LC_2_11_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst11.count_clk_RNI_7_LC_2_11_0  (
            .in0(N__16233),
            .in1(N__16348),
            .in2(_gnd_net_),
            .in3(N__16377),
            .lcout(\b2v_inst11.N_421 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_3_LC_2_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_3_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_3_LC_2_11_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_3_LC_2_11_1  (
            .in0(N__16313),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16255),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_2_LC_2_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_2_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_2_LC_2_11_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_2_LC_2_11_2  (
            .in0(N__16334),
            .in1(N__16289),
            .in2(N__16351),
            .in3(N__16269),
            .lcout(\b2v_inst11.N_373 ),
            .ltout(\b2v_inst11.N_373_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_5_LC_2_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_5_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_5_LC_2_11_3 .LUT_INIT=16'b0011111111111111;
    LogicCell40 \b2v_inst11.count_clk_RNI_5_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__16397),
            .in2(N__16342),
            .in3(N__16232),
            .lcout(\b2v_inst11.count_clk_RNIZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_2_LC_2_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_2_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_2_LC_2_11_4 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \b2v_inst11.count_clk_RNI_2_LC_2_11_4  (
            .in0(N__16335),
            .in1(N__16314),
            .in2(N__16296),
            .in3(N__16268),
            .lcout(),
            .ltout(\b2v_inst11.un2_count_clk_17_0_o3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_3_LC_2_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_3_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_3_LC_2_11_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \b2v_inst11.count_clk_RNI_3_LC_2_11_5  (
            .in0(N__16378),
            .in1(N__16254),
            .in2(N__16240),
            .in3(N__16231),
            .lcout(\b2v_inst11.count_clk_RNIZ0Z_3 ),
            .ltout(\b2v_inst11.count_clk_RNIZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNINJ641_3_LC_2_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNINJ641_3_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNINJ641_3_LC_2_11_6 .LUT_INIT=16'b0000001100000011;
    LogicCell40 \b2v_inst11.count_clk_RNINJ641_3_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__27318),
            .in2(N__16501),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un1_clk_100khz_32_and_i_o2_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIOEM52_1_LC_2_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIOEM52_1_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIOEM52_1_LC_2_11_7 .LUT_INIT=16'b1010100011111100;
    LogicCell40 \b2v_inst11.func_state_RNIOEM52_1_LC_2_11_7  (
            .in0(N__27317),
            .in1(N__29672),
            .in2(N__28751),
            .in3(N__22238),
            .lcout(\b2v_inst11.count_clk_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNISUTE5_12_LC_2_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNISUTE5_12_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNISUTE5_12_LC_2_12_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst11.count_clk_RNISUTE5_12_LC_2_12_0  (
            .in0(N__17495),
            .in1(N__16456),
            .in2(N__16599),
            .in3(N__16467),
            .lcout(\b2v_inst11.count_clkZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_12_LC_2_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_12_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_12_LC_2_12_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.count_clk_12_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16471),
            .in3(N__16565),
            .lcout(\b2v_inst11.count_clk_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34618),
            .ce(N__17538),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_1_LC_2_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_1_LC_2_12_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_1_LC_2_12_2 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \b2v_inst11.count_clk_1_LC_2_12_2  (
            .in0(N__16691),
            .in1(N__16440),
            .in2(_gnd_net_),
            .in3(N__16543),
            .lcout(\b2v_inst11.count_clk_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34618),
            .ce(N__17538),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_0_LC_2_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_0_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_0_LC_2_12_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_0_LC_2_12_3  (
            .in0(N__16439),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16564),
            .lcout(\b2v_inst11.count_clk_RNI_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_LC_2_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_LC_2_12_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_LC_2_12_4  (
            .in0(N__16692),
            .in1(N__16441),
            .in2(_gnd_net_),
            .in3(N__16542),
            .lcout(),
            .ltout(\b2v_inst11.count_clk_RNIZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIT2M95_1_LC_2_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIT2M95_1_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIT2M95_1_LC_2_12_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_clk_RNIT2M95_1_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__16414),
            .in2(N__16408),
            .in3(N__17494),
            .lcout(\b2v_inst11.count_clkZ0Z_1 ),
            .ltout(\b2v_inst11.count_clkZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_1_LC_2_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_1_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_1_LC_2_12_6 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \b2v_inst11.count_clk_RNI_1_LC_2_12_6  (
            .in0(N__16663),
            .in1(N__16713),
            .in2(N__16405),
            .in3(N__16398),
            .lcout(\b2v_inst11.N_187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_1_LC_2_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_1_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_1_LC_2_12_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_1_LC_2_12_7  (
            .in0(N__16712),
            .in1(N__16690),
            .in2(N__16672),
            .in3(N__16662),
            .lcout(\b2v_inst11.count_clk_RNI_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIF6NL_0_LC_2_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIF6NL_0_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIF6NL_0_LC_2_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.func_state_RNIF6NL_0_LC_2_13_0  (
            .in0(N__29365),
            .in1(N__28459),
            .in2(N__23131),
            .in3(N__23342),
            .lcout(\b2v_inst11.N_328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIF6NL_0_0_LC_2_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIF6NL_0_0_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIF6NL_0_0_LC_2_13_1 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \b2v_inst11.func_state_RNIF6NL_0_0_LC_2_13_1  (
            .in0(N__23341),
            .in1(N__29364),
            .in2(N__16651),
            .in3(N__23127),
            .lcout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIVU5C_1_LC_2_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIVU5C_1_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIVU5C_1_LC_2_13_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst11.count_clk_RNIVU5C_1_LC_2_13_2  (
            .in0(N__24868),
            .in1(N__28572),
            .in2(N__19637),
            .in3(N__23340),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIE5T11_1_1_LC_2_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIE5T11_1_1_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIE5T11_1_1_LC_2_13_3 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \b2v_inst11.func_state_RNIE5T11_1_1_LC_2_13_3  (
            .in0(N__21597),
            .in1(N__29363),
            .in2(N__16630),
            .in3(N__28096),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNICC5V2_1_LC_2_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNICC5V2_1_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNICC5V2_1_LC_2_13_4 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \b2v_inst11.func_state_RNICC5V2_1_LC_2_13_4  (
            .in0(N__16627),
            .in1(N__22929),
            .in2(N__16621),
            .in3(N__28457),
            .lcout(\b2v_inst11.func_state_RNICC5V2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIF0H71_1_LC_2_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIF0H71_1_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIF0H71_1_LC_2_13_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \b2v_inst11.func_state_RNIF0H71_1_LC_2_13_7  (
            .in0(N__28458),
            .in1(_gnd_net_),
            .in2(N__22933),
            .in3(N__23343),
            .lcout(\b2v_inst11.N_327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNI2O8H2_LC_2_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNI2O8H2_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNI2O8H2_LC_2_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_10_c_RNI2O8H2_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__19568),
            .in2(_gnd_net_),
            .in3(N__16824),
            .lcout(\b2v_inst11.count_off_1_11 ),
            .ltout(\b2v_inst11.count_off_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI4P25A_11_LC_2_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI4P25A_11_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI4P25A_11_LC_2_14_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_off_RNI4P25A_11_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__16770),
            .in2(N__16513),
            .in3(N__18100),
            .lcout(\b2v_inst11.un3_count_off_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_11_LC_2_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_11_LC_2_14_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_11_LC_2_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_11_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__19571),
            .in2(_gnd_net_),
            .in3(N__16825),
            .lcout(\b2v_inst11.count_offZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34627),
            .ce(N__18151),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIIP81A_0_9_LC_2_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIIP81A_0_9_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIIP81A_0_9_LC_2_14_3 .LUT_INIT=16'b0000000001000111;
    LogicCell40 \b2v_inst11.count_off_RNIIP81A_0_9_LC_2_14_3  (
            .in0(N__16723),
            .in1(N__18102),
            .in2(N__16963),
            .in3(N__17799),
            .lcout(),
            .ltout(\b2v_inst11.un34_clk_100khz_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIQ1RAS1_9_LC_2_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIQ1RAS1_9_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIQ1RAS1_9_LC_2_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.count_off_RNIQ1RAS1_9_LC_2_14_4  (
            .in0(N__16816),
            .in1(N__16759),
            .in2(N__16810),
            .in3(N__16834),
            .lcout(\b2v_inst11.count_off_RNIQ1RAS1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_12_LC_2_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_12_LC_2_14_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_12_LC_2_14_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \b2v_inst11.count_off_12_LC_2_14_5  (
            .in0(N__19570),
            .in1(_gnd_net_),
            .in2(N__16798),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34627),
            .ce(N__18151),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI6S35A_12_LC_2_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI6S35A_12_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI6S35A_12_LC_2_14_6 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst11.count_off_RNI6S35A_12_LC_2_14_6  (
            .in0(N__18101),
            .in1(N__19569),
            .in2(N__16807),
            .in3(N__16794),
            .lcout(\b2v_inst11.count_offZ0Z_12 ),
            .ltout(\b2v_inst11.count_offZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI4P25A_0_11_LC_2_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI4P25A_0_11_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI4P25A_0_11_LC_2_14_7 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \b2v_inst11.count_off_RNI4P25A_0_11_LC_2_14_7  (
            .in0(N__16777),
            .in1(N__16771),
            .in2(N__16762),
            .in3(N__18152),
            .lcout(\b2v_inst11.un34_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_6_LC_2_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_6_LC_2_15_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_6_LC_2_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_6_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__19519),
            .in2(_gnd_net_),
            .in3(N__16939),
            .lcout(\b2v_inst11.count_offZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34631),
            .ce(N__18156),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_9_LC_2_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_9_LC_2_15_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_9_LC_2_15_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \b2v_inst11.count_off_9_LC_2_15_1  (
            .in0(N__19518),
            .in1(_gnd_net_),
            .in2(N__16735),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_offZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34631),
            .ce(N__18156),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNIP80E2_LC_2_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNIP80E2_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNIP80E2_LC_2_15_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_8_c_RNIP80E2_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__19517),
            .in2(_gnd_net_),
            .in3(N__16731),
            .lcout(\b2v_inst11.count_off_1_9 ),
            .ltout(\b2v_inst11.count_off_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIIP81A_9_LC_2_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIIP81A_9_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIIP81A_9_LC_2_15_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst11.count_off_RNIIP81A_9_LC_2_15_3  (
            .in0(N__18143),
            .in1(_gnd_net_),
            .in2(N__16966),
            .in3(N__16962),
            .lcout(\b2v_inst11.un3_count_off_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNIM2TD2_LC_2_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNIM2TD2_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNIM2TD2_LC_2_15_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_5_c_RNIM2TD2_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__19515),
            .in2(_gnd_net_),
            .in3(N__16938),
            .lcout(\b2v_inst11.count_off_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_7_LC_2_15_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_7_LC_2_15_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_7_LC_2_15_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.count_off_7_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19563),
            .in3(N__16906),
            .lcout(\b2v_inst11.count_offZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34631),
            .ce(N__18156),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNIN4UD2_LC_2_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNIN4UD2_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNIN4UD2_LC_2_15_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_6_c_RNIN4UD2_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__19516),
            .in2(_gnd_net_),
            .in3(N__16905),
            .lcout(\b2v_inst11.count_off_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI01TT1_7_LC_2_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI01TT1_7_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI01TT1_7_LC_2_15_7 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \b2v_inst11.dutycycle_RNI01TT1_7_LC_2_15_7  (
            .in0(N__27034),
            .in1(N__26234),
            .in2(_gnd_net_),
            .in3(N__26253),
            .lcout(\b2v_inst11.dutycycle_RNI01TT1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_15_LC_2_16_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_15_LC_2_16_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_15_LC_2_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_15_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(N__19566),
            .in2(_gnd_net_),
            .in3(N__16887),
            .lcout(\b2v_inst11.count_off_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34639),
            .ce(N__18158),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIC575A_15_LC_2_16_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIC575A_15_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIC575A_15_LC_2_16_2 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \b2v_inst11.count_off_RNIC575A_15_LC_2_16_2  (
            .in0(N__19567),
            .in1(N__16894),
            .in2(N__18163),
            .in3(N__16888),
            .lcout(\b2v_inst11.count_offZ0Z_15 ),
            .ltout(\b2v_inst11.count_offZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_15_LC_2_16_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_15_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_15_LC_2_16_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.count_off_RNI_15_LC_2_16_3  (
            .in0(N__16869),
            .in1(N__16855),
            .in2(N__16837),
            .in3(N__17862),
            .lcout(\b2v_inst11.un34_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_8_LC_2_16_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_8_LC_2_16_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_8_LC_2_16_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \b2v_inst11.count_off_8_LC_2_16_4  (
            .in0(N__19565),
            .in1(_gnd_net_),
            .in2(N__17053),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34639),
            .ce(N__18158),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIGM71A_8_LC_2_16_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIGM71A_8_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIGM71A_8_LC_2_16_5 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \b2v_inst11.count_off_RNIGM71A_8_LC_2_16_5  (
            .in0(N__17059),
            .in1(N__19564),
            .in2(N__18157),
            .in3(N__17049),
            .lcout(\b2v_inst11.count_offZ0Z_8 ),
            .ltout(\b2v_inst11.count_offZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIEJ61A_0_7_LC_2_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIEJ61A_0_7_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIEJ61A_0_7_LC_2_16_6 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \b2v_inst11.count_off_RNIEJ61A_0_7_LC_2_16_6  (
            .in0(N__18162),
            .in1(N__17002),
            .in2(N__17026),
            .in3(N__17011),
            .lcout(\b2v_inst11.un34_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIEJ61A_7_LC_2_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIEJ61A_7_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIEJ61A_7_LC_2_16_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_off_RNIEJ61A_7_LC_2_16_7  (
            .in0(N__17010),
            .in1(N__18139),
            .in2(_gnd_net_),
            .in3(N__17001),
            .lcout(\b2v_inst11.un3_count_off_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_4_1_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_4_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_4_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_4_1_0  (
            .in0(_gnd_net_),
            .in1(N__18790),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_1_0_),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_4_1_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_4_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_4_1_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_4_1_1  (
            .in0(_gnd_net_),
            .in1(N__18327),
            .in2(N__20191),
            .in3(N__16978),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_4_1_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_4_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_4_1_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_4_1_2  (
            .in0(_gnd_net_),
            .in1(N__17110),
            .in2(N__18331),
            .in3(N__16975),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_4_1_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_4_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_4_1_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_4_1_3  (
            .in0(_gnd_net_),
            .in1(N__17954),
            .in2(N__17101),
            .in3(N__16972),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_4_1_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_4_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_4_1_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_4_1_4  (
            .in0(_gnd_net_),
            .in1(N__17089),
            .in2(N__17959),
            .in3(N__16969),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_4_1_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_4_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_4_1_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_4_1_5  (
            .in0(N__19999),
            .in1(N__18326),
            .in2(N__17080),
            .in3(N__17119),
            .lcout(\b2v_inst11.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_4_1_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_4_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_4_1_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_4_1_6  (
            .in0(N__17068),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17116),
            .lcout(\b2v_inst11.mult1_un96_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un96_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_4_1_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_4_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_4_1_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_4_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17113),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_2_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_2_0  (
            .in0(_gnd_net_),
            .in1(N__20212),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_2_0_),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_2_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_2_1  (
            .in0(_gnd_net_),
            .in1(N__17183),
            .in2(N__18385),
            .in3(N__17104),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_2_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_2_2  (
            .in0(_gnd_net_),
            .in1(N__17173),
            .in2(N__17188),
            .in3(N__17092),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_2_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_2_3  (
            .in0(_gnd_net_),
            .in1(N__21824),
            .in2(N__17164),
            .in3(N__17083),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_2_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_2_4  (
            .in0(_gnd_net_),
            .in1(N__17152),
            .in2(N__21831),
            .in3(N__17071),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_2_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_2_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_2_5  (
            .in0(N__17952),
            .in1(N__17187),
            .in2(N__17143),
            .in3(N__17062),
            .lcout(\b2v_inst11.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_2_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_2_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_2_6  (
            .in0(N__17131),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17191),
            .lcout(\b2v_inst11.mult1_un89_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_2_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_2_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21823),
            .lcout(\b2v_inst11.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_4_3_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_4_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_4_3_0  (
            .in0(_gnd_net_),
            .in1(N__18766),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_3_0_),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_4_3_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_4_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_4_3_1  (
            .in0(_gnd_net_),
            .in1(N__17201),
            .in2(N__18376),
            .in3(N__17167),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_4_3_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_4_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_4_3_2  (
            .in0(_gnd_net_),
            .in1(N__17263),
            .in2(N__17206),
            .in3(N__17155),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_4_3_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_4_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_4_3_3  (
            .in0(_gnd_net_),
            .in1(N__20069),
            .in2(N__17254),
            .in3(N__17146),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_4_3_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_4_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_4_3_4  (
            .in0(_gnd_net_),
            .in1(N__17242),
            .in2(N__20076),
            .in3(N__17134),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_4_3_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_4_3_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_4_3_5  (
            .in0(N__21822),
            .in1(N__17205),
            .in2(N__17233),
            .in3(N__17125),
            .lcout(\b2v_inst11.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_4_3_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_4_3_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_4_3_6  (
            .in0(N__17221),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17122),
            .lcout(\b2v_inst11.mult1_un82_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_3_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_3_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_3_7  (
            .in0(N__17953),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un85_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_4_4_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_4_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(N__18745),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_4_0_),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_4_4_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_4_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_4_4_1  (
            .in0(_gnd_net_),
            .in1(N__18404),
            .in2(N__19897),
            .in3(N__17257),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_4_4_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_4_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_4_4_2  (
            .in0(_gnd_net_),
            .in1(N__18466),
            .in2(N__18409),
            .in3(N__17245),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_4_4_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_4_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_4_4_3  (
            .in0(_gnd_net_),
            .in1(N__20384),
            .in2(N__18457),
            .in3(N__17236),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_4_4_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_4_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_4_4_4  (
            .in0(_gnd_net_),
            .in1(N__18445),
            .in2(N__20389),
            .in3(N__17224),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_4_4_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_4_4_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_4_4_5  (
            .in0(N__20068),
            .in1(N__18408),
            .in2(N__18436),
            .in3(N__17215),
            .lcout(\b2v_inst11.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_4_4_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_4_4_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_4_4_6  (
            .in0(N__18424),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17212),
            .lcout(\b2v_inst11.mult1_un75_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un75_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_4_4_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_4_4_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_4_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17209),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_4_5_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_4_5_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_4_5_2  (
            .in0(_gnd_net_),
            .in1(N__18934),
            .in2(N__18865),
            .in3(N__18898),
            .lcout(\b2v_inst11.mult1_un40_sum_i_5 ),
            .ltout(\b2v_inst11.mult1_un40_sum_i_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_4_5_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_4_5_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17323),
            .in3(N__18633),
            .lcout(\b2v_inst11.mult1_un47_sum_s_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI4M8F1_10_LC_4_5_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI4M8F1_10_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI4M8F1_10_LC_4_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNI4M8F1_10_LC_4_5_6  (
            .in0(N__17281),
            .in1(N__17295),
            .in2(_gnd_net_),
            .in3(N__30567),
            .lcout(\b2v_inst16.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_10_LC_4_5_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_10_LC_4_5_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_10_LC_4_5_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_10_LC_4_5_7  (
            .in0(N__17296),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34634),
            .ce(N__30605),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_6_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18955),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_6_0_),
            .carryout(\b2v_inst11.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_6_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_6_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17350),
            .in3(N__17275),
            .lcout(\b2v_inst11.mult1_un47_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un47_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un47_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_6_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_6_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17332),
            .in3(N__17272),
            .lcout(\b2v_inst11.mult1_un47_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un47_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un47_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_6_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_6_3  (
            .in0(_gnd_net_),
            .in1(N__20118),
            .in2(N__17341),
            .in3(N__17269),
            .lcout(\b2v_inst11.mult1_un47_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un47_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un47_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_4_6_4 .C_ON=1'b0;
    defparam \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_4_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_4_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17266),
            .lcout(\b2v_inst11.mult1_un47_sum_cry_5_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_6_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_6_5 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_6_5  (
            .in0(N__18500),
            .in1(N__18501),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un47_sum_l_fx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_4_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_4_6_6 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_4_6_6  (
            .in0(N__18671),
            .in1(N__18672),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un47_sum_l_fx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_en_LC_4_6_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_en_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_en_LC_4_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst200.count_en_LC_4_6_7  (
            .in0(_gnd_net_),
            .in1(N__33717),
            .in2(_gnd_net_),
            .in3(N__33082),
            .lcout(\b2v_inst200.count_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_4_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_4_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18925),
            .lcout(\b2v_inst11.un1_dutycycle_53_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_4_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_4_7_1 .LUT_INIT=16'b1111101000000101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_4_7_1  (
            .in0(N__18927),
            .in1(_gnd_net_),
            .in2(N__18897),
            .in3(N__18858),
            .lcout(\b2v_inst11.mult1_un40_sum_i_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18951),
            .lcout(\b2v_inst11.mult1_un47_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_4_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_4_7_5 .LUT_INIT=16'b1010010110100101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_4_7_5  (
            .in0(N__18926),
            .in1(_gnd_net_),
            .in2(N__18896),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un47_sum_s_4_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_4_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_4_8_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_4_8_0  (
            .in0(N__18783),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNI_0_LC_4_8_2 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI_0_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI_0_LC_4_8_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst36.curr_state_RNI_0_LC_4_8_2  (
            .in0(N__30403),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.N_2925_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_3_LC_4_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_3_LC_4_8_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_3_LC_4_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_3_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17572),
            .lcout(\b2v_inst11.count_clk_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34620),
            .ce(N__17526),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI3JFN6_13_LC_4_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI3JFN6_13_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI3JFN6_13_LC_4_9_0 .LUT_INIT=16'b0111010100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI3JFN6_13_LC_4_9_0  (
            .in0(N__27759),
            .in1(N__22253),
            .in2(N__17401),
            .in3(N__27596),
            .lcout(\b2v_inst11.dutycycle_en_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIAI7C4_13_LC_4_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIAI7C4_13_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIAI7C4_13_LC_4_9_1 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \b2v_inst11.dutycycle_RNIAI7C4_13_LC_4_9_1  (
            .in0(N__21313),
            .in1(N__22586),
            .in2(_gnd_net_),
            .in3(N__22396),
            .lcout(\b2v_inst11.N_150_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIAI7C4_14_LC_4_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIAI7C4_14_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIAI7C4_14_LC_4_9_2 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNIAI7C4_14_LC_4_9_2  (
            .in0(N__22587),
            .in1(_gnd_net_),
            .in2(N__22402),
            .in3(N__21244),
            .lcout(),
            .ltout(\b2v_inst11.N_152_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI3JFN6_14_LC_4_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI3JFN6_14_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI3JFN6_14_LC_4_9_3 .LUT_INIT=16'b0010000010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI3JFN6_14_LC_4_9_3  (
            .in0(N__27597),
            .in1(N__22255),
            .in2(N__17392),
            .in3(N__27760),
            .lcout(\b2v_inst11.dutycycle_en_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI4UUA8_15_LC_4_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI4UUA8_15_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI4UUA8_15_LC_4_9_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI4UUA8_15_LC_4_9_4  (
            .in0(N__27292),
            .in1(N__17373),
            .in2(N__21106),
            .in3(N__17383),
            .lcout(\b2v_inst11.dutycycleZ0Z_12 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIAI7C4_15_LC_4_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIAI7C4_15_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIAI7C4_15_LC_4_9_5 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \b2v_inst11.dutycycle_RNIAI7C4_15_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(N__22588),
            .in2(N__17389),
            .in3(N__22400),
            .lcout(),
            .ltout(\b2v_inst11.N_155_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI3JFN6_15_LC_4_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI3JFN6_15_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI3JFN6_15_LC_4_9_6 .LUT_INIT=16'b0111010100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI3JFN6_15_LC_4_9_6  (
            .in0(N__27758),
            .in1(N__22254),
            .in2(N__17386),
            .in3(N__27595),
            .lcout(\b2v_inst11.dutycycle_en_12 ),
            .ltout(\b2v_inst11.dutycycle_en_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_15_LC_4_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_15_LC_4_9_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_15_LC_4_9_7 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \b2v_inst11.dutycycle_15_LC_4_9_7  (
            .in0(N__21105),
            .in1(N__17374),
            .in2(N__17377),
            .in3(N__27316),
            .lcout(\b2v_inst11.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34613),
            .ce(),
            .sr(N__24232));
    defparam \b2v_inst11.dutycycle_13_LC_4_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_13_LC_4_10_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_13_LC_4_10_0 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \b2v_inst11.dutycycle_13_LC_4_10_0  (
            .in0(N__17605),
            .in1(N__21265),
            .in2(N__17596),
            .in3(N__27315),
            .lcout(\b2v_inst11.dutycycleZ1Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34619),
            .ce(),
            .sr(N__24227));
    defparam \b2v_inst11.dutycycle_RNI_2_12_LC_4_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_12_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_12_LC_4_10_1 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_12_LC_4_10_1  (
            .in0(N__21434),
            .in1(N__19339),
            .in2(_gnd_net_),
            .in3(N__22359),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_2Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_10_9_LC_4_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_10_9_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_10_9_LC_4_10_2 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_10_9_LC_4_10_2  (
            .in0(N__19340),
            .in1(N__19011),
            .in2(N__17611),
            .in3(N__21014),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_10Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_13_LC_4_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_13_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_13_LC_4_10_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_13_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(N__21246),
            .in2(N__17608),
            .in3(N__21306),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI0OSA8_13_LC_4_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI0OSA8_13_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI0OSA8_13_LC_4_10_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \b2v_inst11.dutycycle_RNI0OSA8_13_LC_4_10_4  (
            .in0(N__17604),
            .in1(N__21264),
            .in2(N__17595),
            .in3(N__27314),
            .lcout(\b2v_inst11.dutycycleZ0Z_9 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_13_LC_4_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_13_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_13_LC_4_10_5 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_13_LC_4_10_5  (
            .in0(N__21433),
            .in1(_gnd_net_),
            .in2(N__17581),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_0Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_10_LC_4_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_10_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_10_LC_4_10_6 .LUT_INIT=16'b0000001100001011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_10_LC_4_10_6  (
            .in0(N__22360),
            .in1(N__19345),
            .in2(N__17578),
            .in3(N__19177),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_10 ),
            .ltout(\b2v_inst11.dutycycle_RNI_1Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_14_LC_4_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_14_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_14_LC_4_10_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_14_LC_4_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17575),
            .in3(N__21245),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIHTFQ_8_LC_4_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIHTFQ_8_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIHTFQ_8_LC_4_11_0 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIHTFQ_8_LC_4_11_0  (
            .in0(N__17672),
            .in1(N__26954),
            .in2(_gnd_net_),
            .in3(N__26879),
            .lcout(\b2v_inst11.dutycycle_RNIHTFQZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIJU083_8_LC_4_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIJU083_8_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIJU083_8_LC_4_11_1 .LUT_INIT=16'b1111111101001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIJU083_8_LC_4_11_1  (
            .in0(N__22593),
            .in1(N__28117),
            .in2(N__22783),
            .in3(N__22240),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNIJU083Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNITG8K7_8_LC_4_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNITG8K7_8_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNITG8K7_8_LC_4_11_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \b2v_inst11.dutycycle_RNITG8K7_8_LC_4_11_2  (
            .in0(N__27312),
            .in1(_gnd_net_),
            .in2(N__17695),
            .in3(N__17647),
            .lcout(\b2v_inst11.N_108_f0 ),
            .ltout(\b2v_inst11.N_108_f0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_8_LC_4_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_8_LC_4_11_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_8_LC_4_11_3 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \b2v_inst11.dutycycle_8_LC_4_11_3  (
            .in0(N__17680),
            .in1(N__27780),
            .in2(N__17692),
            .in3(N__17674),
            .lcout(\b2v_inst11.dutycycleZ1Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34624),
            .ce(),
            .sr(N__24231));
    defparam \b2v_inst11.dutycycle_RNI2NK31_8_LC_4_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI2NK31_8_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI2NK31_8_LC_4_11_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI2NK31_8_LC_4_11_4  (
            .in0(N__17673),
            .in1(N__26955),
            .in2(N__21034),
            .in3(N__26880),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI2NK31Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIA8B23_8_LC_4_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIA8B23_8_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIA8B23_8_LC_4_11_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNIA8B23_8_LC_4_11_5  (
            .in0(_gnd_net_),
            .in1(N__17689),
            .in2(N__17683),
            .in3(N__27313),
            .lcout(\b2v_inst11.dutycycle_e_1_8 ),
            .ltout(\b2v_inst11.dutycycle_e_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI9QKHC_8_LC_4_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI9QKHC_8_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI9QKHC_8_LC_4_11_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI9QKHC_8_LC_4_11_6  (
            .in0(N__17671),
            .in1(N__17659),
            .in2(N__17653),
            .in3(N__27778),
            .lcout(\b2v_inst11.dutycycleZ0Z_1 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIJU083_0_8_LC_4_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIJU083_0_8_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIJU083_0_8_LC_4_11_7 .LUT_INIT=16'b1111111100111111;
    LogicCell40 \b2v_inst11.dutycycle_RNIJU083_0_8_LC_4_11_7  (
            .in0(_gnd_net_),
            .in1(N__22592),
            .in2(N__17650),
            .in3(N__22239),
            .lcout(\b2v_inst11.dutycycle_RNIJU083_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIM6F44_0_LC_4_12_0 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIM6F44_0_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIM6F44_0_LC_4_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_RNIM6F44_0_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33778),
            .lcout(delayed_vccin_vccinaux_ok_RNIM6F44_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_9_LC_4_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_9_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_9_LC_4_12_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_9_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__21013),
            .in2(_gnd_net_),
            .in3(N__22361),
            .lcout(\b2v_inst11.un1_dutycycle_53_41_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_12_LC_4_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_12_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_12_LC_4_12_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_12_LC_4_12_2  (
            .in0(N__21417),
            .in1(N__19337),
            .in2(N__24382),
            .in3(N__19432),
            .lcout(\b2v_inst11.g0_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_1_1_LC_4_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_1_1_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_1_1_LC_4_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.func_state_RNI_1_1_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28455),
            .lcout(\b2v_inst11.func_state_RNI_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIT4D71_1_LC_4_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIT4D71_1_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIT4D71_1_LC_4_12_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst11.func_state_RNIT4D71_1_LC_4_12_4  (
            .in0(N__28456),
            .in1(N__17986),
            .in2(N__29362),
            .in3(N__26964),
            .lcout(),
            .ltout(\b2v_inst11.N_289_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIFIVO1_LC_4_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIFIVO1_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIFIVO1_LC_4_12_5 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIFIVO1_LC_4_12_5  (
            .in0(N__28292),
            .in1(N__20776),
            .in2(N__17707),
            .in3(N__21591),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_1_0_iv_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI666T2_LC_4_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI666T2_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI666T2_LC_4_12_6 .LUT_INIT=16'b1111000111111111;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI666T2_LC_4_12_6  (
            .in0(N__28291),
            .in1(N__28708),
            .in2(N__17704),
            .in3(N__29099),
            .lcout(\b2v_inst11.N_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_12_LC_4_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_12_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_12_LC_4_12_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_12_LC_4_12_7  (
            .in0(N__19431),
            .in1(N__18580),
            .in2(N__19344),
            .in3(N__21416),
            .lcout(\b2v_inst11.m15_e_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_12_LC_4_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_12_LC_4_13_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_12_LC_4_13_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \b2v_inst11.dutycycle_12_LC_4_13_0  (
            .in0(N__27296),
            .in1(N__17761),
            .in2(N__17755),
            .in3(N__21355),
            .lcout(\b2v_inst11.dutycycleZ1Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34633),
            .ce(),
            .sr(N__24238));
    defparam \b2v_inst11.dutycycle_RNINJ641_11_LC_4_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNINJ641_11_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNINJ641_11_LC_4_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNINJ641_11_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__19318),
            .in2(_gnd_net_),
            .in3(N__27294),
            .lcout(),
            .ltout(\b2v_inst11.N_302_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIGKEF3_11_LC_4_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIGKEF3_11_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIGKEF3_11_LC_4_13_2 .LUT_INIT=16'b0101011100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNIGKEF3_11_LC_4_13_2  (
            .in0(N__27779),
            .in1(N__17734),
            .in2(N__17701),
            .in3(N__27599),
            .lcout(\b2v_inst11.dutycycle_RNIGKEF3Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNINJ641_12_LC_4_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNINJ641_12_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNINJ641_12_LC_4_13_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNINJ641_12_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__27295),
            .in2(_gnd_net_),
            .in3(N__21415),
            .lcout(),
            .ltout(\b2v_inst11.N_301_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIGKEF3_12_LC_4_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIGKEF3_12_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIGKEF3_12_LC_4_13_4 .LUT_INIT=16'b0010001000101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIGKEF3_12_LC_4_13_4  (
            .in0(N__27598),
            .in1(N__27777),
            .in2(N__17698),
            .in3(N__17733),
            .lcout(\b2v_inst11.dutycycle_RNIGKEF3Z0Z_12 ),
            .ltout(\b2v_inst11.dutycycle_RNIGKEF3Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIBMQ25_12_LC_4_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIBMQ25_12_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIBMQ25_12_LC_4_13_5 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \b2v_inst11.dutycycle_RNIBMQ25_12_LC_4_13_5  (
            .in0(N__21354),
            .in1(N__17751),
            .in2(N__17743),
            .in3(N__27293),
            .lcout(\b2v_inst11.dutycycleZ0Z_10 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_12_LC_4_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_12_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_12_LC_4_13_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_12_LC_4_13_6  (
            .in0(N__19319),
            .in1(_gnd_net_),
            .in2(N__17740),
            .in3(N__19015),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_56_a0_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_13_LC_4_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_13_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_13_LC_4_13_7 .LUT_INIT=16'b1111111101010000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_13_LC_4_13_7  (
            .in0(N__19084),
            .in1(N__21335),
            .in2(N__17737),
            .in3(N__19246),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIAI7C4_2_LC_4_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIAI7C4_2_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIAI7C4_2_LC_4_14_0 .LUT_INIT=16'b1010111110001111;
    LogicCell40 \b2v_inst11.dutycycle_RNIAI7C4_2_LC_4_14_0  (
            .in0(N__19357),
            .in1(N__27304),
            .in2(N__22603),
            .in3(N__19402),
            .lcout(\b2v_inst11.N_232_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_1_LC_4_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_1_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_1_LC_4_14_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_1_LC_4_14_1  (
            .in0(N__23375),
            .in1(N__29112),
            .in2(N__23286),
            .in3(N__29236),
            .lcout(),
            .ltout(\b2v_inst11.un1_func_state25_6_0_o_N_325_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_4_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_4_14_2 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_4_14_2  (
            .in0(N__17719),
            .in1(N__28462),
            .in2(N__17725),
            .in3(N__19605),
            .lcout(),
            .ltout(\b2v_inst11.un1_func_state25_6_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_en_LC_4_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_en_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_en_LC_4_14_3 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \b2v_inst11.count_off_en_LC_4_14_3  (
            .in0(N__27619),
            .in1(N__21505),
            .in2(N__17722),
            .in3(N__17713),
            .lcout(\b2v_inst11.count_off_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_LC_4_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_LC_4_14_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_LC_4_14_4  (
            .in0(N__25086),
            .in1(N__28461),
            .in2(N__19396),
            .in3(N__23374),
            .lcout(\b2v_inst11.un1_func_state25_6_0_o_N_323_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_0_LC_4_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_0_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_0_LC_4_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_0_LC_4_14_5  (
            .in0(N__22875),
            .in1(N__29111),
            .in2(N__23285),
            .in3(N__19641),
            .lcout(\b2v_inst11.un1_func_state25_6_0_o_N_324_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINJ641_1_LC_4_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINJ641_1_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINJ641_1_LC_4_14_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.func_state_RNINJ641_1_LC_4_14_6  (
            .in0(N__23054),
            .in1(N__28460),
            .in2(N__23382),
            .in3(N__24313),
            .lcout(\b2v_inst11.N_322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI51SU9_1_LC_4_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI51SU9_1_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI51SU9_1_LC_4_15_0 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \b2v_inst11.count_off_RNI51SU9_1_LC_4_15_0  (
            .in0(N__17869),
            .in1(N__19468),
            .in2(N__18077),
            .in3(N__17878),
            .lcout(\b2v_inst11.count_offZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI40SU9_0_LC_4_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI40SU9_0_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI40SU9_0_LC_4_15_1 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \b2v_inst11.count_off_RNI40SU9_0_LC_4_15_1  (
            .in0(N__19467),
            .in1(N__17827),
            .in2(N__17852),
            .in3(N__18033),
            .lcout(\b2v_inst11.count_offZ0Z_0 ),
            .ltout(\b2v_inst11.count_offZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_1_LC_4_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_1_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_1_LC_4_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.count_off_RNI_1_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17914),
            .in3(N__17897),
            .lcout(\b2v_inst11.count_off_RNIZ0Z_1 ),
            .ltout(\b2v_inst11.count_off_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_1_LC_4_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_1_LC_4_15_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_1_LC_4_15_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \b2v_inst11.count_off_1_LC_4_15_3  (
            .in0(N__19471),
            .in1(_gnd_net_),
            .in2(N__17872),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34648),
            .ce(N__18037),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_0_LC_4_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_0_LC_4_15_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_0_LC_4_15_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst11.count_off_0_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__17845),
            .in2(_gnd_net_),
            .in3(N__19472),
            .lcout(\b2v_inst11.count_off_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34648),
            .ce(N__18037),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_10_LC_4_15_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_10_LC_4_15_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_10_LC_4_15_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_10_LC_4_15_5  (
            .in0(N__19469),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17811),
            .lcout(\b2v_inst11.count_off_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34648),
            .ce(N__18037),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIRAR1A_10_LC_4_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIRAR1A_10_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIRAR1A_10_LC_4_15_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst11.count_off_RNIRAR1A_10_LC_4_15_6  (
            .in0(N__18038),
            .in1(N__17821),
            .in2(N__17815),
            .in3(N__19466),
            .lcout(\b2v_inst11.count_offZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_13_LC_4_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_13_LC_4_15_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_13_LC_4_15_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_13_LC_4_15_7  (
            .in0(N__19470),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17776),
            .lcout(\b2v_inst11.count_off_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34648),
            .ce(N__18037),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIVU5C_0_LC_4_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIVU5C_0_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIVU5C_0_LC_4_16_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.func_state_RNIVU5C_0_LC_4_16_7  (
            .in0(N__28488),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24316),
            .lcout(\b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_1_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_1_0  (
            .in0(_gnd_net_),
            .in1(N__18826),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_1_0_),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_1_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_1_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_1_1  (
            .in0(_gnd_net_),
            .in1(N__18185),
            .in2(N__18367),
            .in3(N__17977),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_1_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_1_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_1_2  (
            .in0(_gnd_net_),
            .in1(N__18298),
            .in2(N__18190),
            .in3(N__17974),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_1_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_1_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_1_3  (
            .in0(_gnd_net_),
            .in1(N__18351),
            .in2(N__18283),
            .in3(N__17971),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_1_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_1_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_1_4  (
            .in0(_gnd_net_),
            .in1(N__18262),
            .in2(N__18355),
            .in3(N__17968),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_1_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_1_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_1_5  (
            .in0(N__20148),
            .in1(N__18189),
            .in2(N__18247),
            .in3(N__17965),
            .lcout(\b2v_inst11.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_1_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_1_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_1_6  (
            .in0(N__18211),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17962),
            .lcout(\b2v_inst11.mult1_un110_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_1_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_1_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17958),
            .lcout(\b2v_inst11.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_5_2_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_5_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_5_2_0  (
            .in0(_gnd_net_),
            .in1(N__18808),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_2_0_),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_5_2_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_5_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_5_2_1  (
            .in0(_gnd_net_),
            .in1(N__18230),
            .in2(N__18316),
            .in3(N__18292),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_5_2_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_5_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_5_2_2  (
            .in0(_gnd_net_),
            .in1(N__18289),
            .in2(N__18235),
            .in3(N__18274),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_5_2_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_5_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_5_2_3  (
            .in0(_gnd_net_),
            .in1(N__20000),
            .in2(N__18271),
            .in3(N__18256),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_5_2_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_5_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_5_2_4  (
            .in0(_gnd_net_),
            .in1(N__18253),
            .in2(N__20007),
            .in3(N__18238),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_5_2_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_5_2_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_5_2_5  (
            .in0(N__18349),
            .in1(N__18234),
            .in2(N__18220),
            .in3(N__18205),
            .lcout(\b2v_inst11.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_5_2_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_5_2_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_5_2_6  (
            .in0(N__18202),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18196),
            .lcout(\b2v_inst11.mult1_un103_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un103_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_5_2_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_5_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_5_2_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_5_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18193),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_5_3_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_5_3_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(N__19728),
            .in2(_gnd_net_),
            .in3(N__20272),
            .lcout(\b2v_inst11.mult1_un131_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_3_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_3_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18825),
            .lcout(\b2v_inst11.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_3_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_3_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_5_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20271),
            .lcout(\b2v_inst11.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_5_3_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_5_3_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_5_3_3  (
            .in0(N__20273),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19944),
            .lcout(\b2v_inst11.mult1_un131_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_3_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_3_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18762),
            .lcout(\b2v_inst11.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_3_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_3_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18741),
            .lcout(\b2v_inst11.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_3_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_3_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18807),
            .lcout(\b2v_inst11.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_3_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_3_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_5_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18350),
            .lcout(\b2v_inst11.un85_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_4_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_4_0  (
            .in0(_gnd_net_),
            .in1(N__19914),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_4_0_),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_2_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_4_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(N__20171),
            .in2(N__20398),
            .in3(N__18460),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_2_c ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_3_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_4_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_4_2  (
            .in0(_gnd_net_),
            .in1(N__18394),
            .in2(N__20176),
            .in3(N__18448),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_3_c ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_4_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_4_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_4_3  (
            .in0(_gnd_net_),
            .in1(N__18562),
            .in2(N__20050),
            .in3(N__18439),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_4_c ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_5_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_4_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_4_4  (
            .in0(_gnd_net_),
            .in1(N__18553),
            .in2(N__20049),
            .in3(N__18427),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_5_c ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_6_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_4_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_4_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_4_5  (
            .in0(N__20383),
            .in1(N__20175),
            .in2(N__18544),
            .in3(N__18418),
            .lcout(\b2v_inst11.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_6_c ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_4_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_4_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_4_6  (
            .in0(N__18532),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18415),
            .lcout(\b2v_inst11.mult1_un68_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un68_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_4_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_4_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18412),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_5_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_5_0  (
            .in0(_gnd_net_),
            .in1(N__20415),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_5_0_),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_5_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(N__20422),
            .in2(N__18597),
            .in3(N__18388),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_5_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(N__18593),
            .in2(N__18514),
            .in3(N__18556),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_5_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(N__18475),
            .in2(N__18619),
            .in3(N__18547),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_5_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(N__18618),
            .in2(N__18712),
            .in3(N__18535),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_5_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_5_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_5_5  (
            .in0(N__20038),
            .in1(N__18691),
            .in2(N__18598),
            .in3(N__18526),
            .lcout(\b2v_inst11.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_5_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_5_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18655),
            .in3(N__18523),
            .lcout(\b2v_inst11.mult1_un61_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_5_6_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_5_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20443),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_6_0_),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_5_6_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_5_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_5_6_1  (
            .in0(_gnd_net_),
            .in1(N__18520),
            .in2(_gnd_net_),
            .in3(N__18505),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_5_6_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_5_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__18502),
            .in2(N__18484),
            .in3(N__18469),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_5_6_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_5_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(N__20096),
            .in2(N__18721),
            .in3(N__18703),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_5_6_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_5_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_5_6_4  (
            .in0(_gnd_net_),
            .in1(N__20114),
            .in2(N__18700),
            .in3(N__18685),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_5_6_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_5_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_5_6_5  (
            .in0(N__18614),
            .in1(N__18682),
            .in2(N__18676),
            .in3(N__18646),
            .lcout(\b2v_inst11.mult1_un61_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_5_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_5_6_6 .LUT_INIT=16'b0000110011110011;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_5_6_6  (
            .in0(_gnd_net_),
            .in1(N__18643),
            .in2(N__18637),
            .in3(N__18622),
            .lcout(\b2v_inst11.mult1_un54_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un54_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_5_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_5_6_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18601),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_LC_5_7_0 .C_ON=1'b1;
    defparam \b2v_inst11.dutycycle_RNI_0_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_LC_5_7_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(N__24819),
            .in2(N__25597),
            .in3(N__25385),
            .lcout(\b2v_inst11.m15_e_2 ),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_0_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_5_7_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_5_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_5_7_1  (
            .in0(_gnd_net_),
            .in1(N__25594),
            .in2(N__20521),
            .in3(N__18568),
            .lcout(\b2v_inst11.mult1_un138_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_0_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_5_7_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_5_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(N__27428),
            .in2(N__20464),
            .in3(N__18565),
            .lcout(\b2v_inst11.mult1_un131_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_1_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_5_7_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_5_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(N__23992),
            .in2(N__27435),
            .in3(N__18832),
            .lcout(\b2v_inst11.mult1_un124_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_2_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_3_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_5_7_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_5_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_5_7_4  (
            .in0(_gnd_net_),
            .in1(N__22465),
            .in2(N__22453),
            .in3(N__18829),
            .lcout(\b2v_inst11.mult1_un117_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_3_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_4_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_5_7_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_5_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_5_7_5  (
            .in0(_gnd_net_),
            .in1(N__26766),
            .in2(N__22483),
            .in3(N__18811),
            .lcout(\b2v_inst11.mult1_un110_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_4_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_5_7_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_5_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_5_7_6  (
            .in0(_gnd_net_),
            .in1(N__20449),
            .in2(N__26779),
            .in3(N__18793),
            .lcout(\b2v_inst11.mult1_un103_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_5_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_6_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_5_7_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_5_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_5_7_7  (
            .in0(_gnd_net_),
            .in1(N__20455),
            .in2(N__22363),
            .in3(N__18772),
            .lcout(\b2v_inst11.mult1_un96_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_6_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_5_8_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_5_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(N__20892),
            .in2(N__19096),
            .in3(N__18769),
            .lcout(\b2v_inst11.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_5_8_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_5_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__21442),
            .in2(N__19192),
            .in3(N__18748),
            .lcout(\b2v_inst11.mult1_un82_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_8_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_9_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_5_8_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_5_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_5_8_2  (
            .in0(_gnd_net_),
            .in1(N__21324),
            .in2(N__19060),
            .in3(N__18727),
            .lcout(\b2v_inst11.mult1_un75_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_9_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_5_8_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_5_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_5_8_3  (
            .in0(_gnd_net_),
            .in1(N__21224),
            .in2(N__19036),
            .in3(N__18724),
            .lcout(\b2v_inst11.mult1_un68_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_10 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_5_8_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_5_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_5_8_4  (
            .in0(_gnd_net_),
            .in1(N__21140),
            .in2(N__19027),
            .in3(N__18985),
            .lcout(\b2v_inst11.mult1_un61_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_11 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_5_8_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_5_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_5_8_5  (
            .in0(_gnd_net_),
            .in1(N__21325),
            .in2(N__18982),
            .in3(N__18967),
            .lcout(\b2v_inst11.mult1_un54_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_12 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_5_8_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_5_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_5_8_6  (
            .in0(_gnd_net_),
            .in1(N__18964),
            .in2(N__21240),
            .in3(N__18937),
            .lcout(\b2v_inst11.mult1_un47_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_13 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_5_8_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_5_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_5_8_7  (
            .in0(_gnd_net_),
            .in1(N__18838),
            .in2(N__21154),
            .in3(N__18910),
            .lcout(\b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_14 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_5_9_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_5_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_5_9_0  (
            .in0(_gnd_net_),
            .in1(N__21155),
            .in2(N__18907),
            .in3(N__18871),
            .lcout(\b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\b2v_inst11.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.CO2_THRU_LUT4_0_LC_5_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.CO2_THRU_LUT4_0_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.CO2_THRU_LUT4_0_LC_5_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.CO2_THRU_LUT4_0_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18868),
            .lcout(\b2v_inst11.CO2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_15_LC_5_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_15_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_15_LC_5_9_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_15_LC_5_9_2  (
            .in0(N__21149),
            .in1(N__21223),
            .in2(_gnd_net_),
            .in3(N__18844),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_9_LC_5_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_9_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_9_LC_5_9_3 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_9_LC_5_9_3  (
            .in0(N__26232),
            .in1(N__22779),
            .in2(N__22362),
            .in3(N__21011),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_44_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_9_LC_5_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_9_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_9_LC_5_9_4 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_9_LC_5_9_4  (
            .in0(N__21012),
            .in1(N__18991),
            .in2(N__19042),
            .in3(N__20659),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_6Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_11_LC_5_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_11_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_11_LC_5_9_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_11_LC_5_9_5  (
            .in0(N__22354),
            .in1(N__21231),
            .in2(N__19039),
            .in3(N__20891),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_10_LC_5_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_10_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_10_LC_5_9_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_10_LC_5_9_6  (
            .in0(N__22778),
            .in1(N__28972),
            .in2(N__28036),
            .in3(N__22350),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_15_LC_5_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_15_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_15_LC_5_9_7 .LUT_INIT=16'b0011110011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_15_LC_5_9_7  (
            .in0(N__21156),
            .in1(N__18997),
            .in2(N__19213),
            .in3(N__20647),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_7_LC_5_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_7_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_7_LC_5_10_0 .LUT_INIT=16'b0100010000100010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_7_LC_5_10_0  (
            .in0(N__26213),
            .in1(N__22728),
            .in2(_gnd_net_),
            .in3(N__19142),
            .lcout(),
            .ltout(\b2v_inst11.un1_m7_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_4_LC_5_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_4_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_4_LC_5_10_1 .LUT_INIT=16'b0010010110110101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_4_LC_5_10_1  (
            .in0(N__22729),
            .in1(N__28014),
            .in2(N__19018),
            .in3(N__28934),
            .lcout(\b2v_inst11.un1_i3_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_11_LC_5_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_11_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_11_LC_5_10_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_11_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__20890),
            .in2(_gnd_net_),
            .in3(N__21436),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_4_LC_5_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_4_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_4_LC_5_10_3 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_4_LC_5_10_3  (
            .in0(N__28016),
            .in1(N__28936),
            .in2(N__19154),
            .in3(N__19338),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_4_LC_5_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_4_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_4_LC_5_10_4 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_4_LC_5_10_4  (
            .in0(N__26215),
            .in1(N__22734),
            .in2(N__28973),
            .in3(N__28018),
            .lcout(\b2v_inst11.un1_dutycycle_53_44_0_2_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_4_LC_5_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_4_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_4_LC_5_10_5 .LUT_INIT=16'b0000001110101011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_4_LC_5_10_5  (
            .in0(N__19143),
            .in1(N__28935),
            .in2(N__22771),
            .in3(N__26214),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_39_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_9_LC_5_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_9_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_9_LC_5_10_6 .LUT_INIT=16'b1110111000001110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_9_LC_5_10_6  (
            .in0(N__20996),
            .in1(N__22733),
            .in2(N__19078),
            .in3(N__28017),
            .lcout(\b2v_inst11.un1_dutycycle_53_39_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_LC_5_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_LC_5_10_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_LC_5_10_7  (
            .in0(N__22414),
            .in1(N__22761),
            .in2(N__19155),
            .in3(N__20674),
            .lcout(\b2v_inst11.N_357 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_9_LC_5_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_9_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_9_LC_5_11_0 .LUT_INIT=16'b0000010111001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_9_LC_5_11_0  (
            .in0(N__20592),
            .in1(N__22645),
            .in2(N__28032),
            .in3(N__20957),
            .lcout(\b2v_inst11.dutycycle_RNI_8Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNINJ641_9_LC_5_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNINJ641_9_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNINJ641_9_LC_5_11_1 .LUT_INIT=16'b0000000000011111;
    LogicCell40 \b2v_inst11.dutycycle_RNINJ641_9_LC_5_11_1  (
            .in0(N__27305),
            .in1(N__28107),
            .in2(N__19156),
            .in3(N__22241),
            .lcout(\b2v_inst11.dutycycle_eena_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_LC_5_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_LC_5_11_2 .LUT_INIT=16'b1110110011101110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_LC_5_11_2  (
            .in0(N__22776),
            .in1(N__26189),
            .in2(N__28974),
            .in3(N__19150),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_39_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_13_LC_5_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_13_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_13_LC_5_11_3 .LUT_INIT=16'b0011111111000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_13_LC_5_11_3  (
            .in0(N__21314),
            .in1(N__19075),
            .in2(N__19069),
            .in3(N__19066),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_9_LC_5_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_9_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_9_LC_5_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_9_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20956),
            .lcout(\b2v_inst11.dutycycle_RNI_5Z0Z_9 ),
            .ltout(\b2v_inst11.dutycycle_RNI_5Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_9_LC_5_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_9_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_9_LC_5_11_5 .LUT_INIT=16'b0011000001110111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_9_LC_5_11_5  (
            .in0(N__20958),
            .in1(N__28940),
            .in2(N__19048),
            .in3(N__22775),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_10_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_LC_5_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_LC_5_11_6 .LUT_INIT=16'b1100111010001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_LC_5_11_6  (
            .in0(N__28024),
            .in1(N__26188),
            .in2(N__19045),
            .in3(N__22764),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNIZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_12_LC_5_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_12_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_12_LC_5_11_7 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_12_LC_5_11_7  (
            .in0(N__20959),
            .in1(N__22777),
            .in2(N__19195),
            .in3(N__21440),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_4_LC_5_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_4_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_4_LC_5_12_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_4_LC_5_12_0  (
            .in0(N__28971),
            .in1(N__19162),
            .in2(_gnd_net_),
            .in3(N__19111),
            .lcout(),
            .ltout(\b2v_inst11.m18_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_11_9_LC_5_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_11_9_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_11_9_LC_5_12_1 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_11_9_LC_5_12_1  (
            .in0(N__19168),
            .in1(N__20994),
            .in2(N__19180),
            .in3(N__28011),
            .lcout(\b2v_inst11.dutycycle_RNI_11Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_7_LC_5_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_7_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_7_LC_5_12_2 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_7_LC_5_12_2  (
            .in0(N__19141),
            .in1(N__26203),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_7_LC_5_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_7_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_7_LC_5_12_3 .LUT_INIT=16'b0101010101011101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_7_LC_5_12_3  (
            .in0(N__22725),
            .in1(N__19140),
            .in2(N__26230),
            .in3(N__28010),
            .lcout(\b2v_inst11.dutycycle_RNI_5Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_7_LC_5_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_7_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_7_LC_5_12_4 .LUT_INIT=16'b0010001011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_7_LC_5_12_4  (
            .in0(N__19139),
            .in1(N__26199),
            .in2(_gnd_net_),
            .in3(N__22726),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_7_LC_5_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_7_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_7_LC_5_12_5 .LUT_INIT=16'b1010100101101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_7_LC_5_12_5  (
            .in0(N__19201),
            .in1(N__19105),
            .in2(N__26231),
            .in3(N__28012),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_11_LC_5_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_11_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_11_LC_5_12_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_11_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19099),
            .in3(N__20880),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_9_LC_5_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_9_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_9_LC_5_12_7 .LUT_INIT=16'b1100110010001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_9_LC_5_12_7  (
            .in0(N__22727),
            .in1(N__20995),
            .in2(N__22615),
            .in3(N__22348),
            .lcout(\b2v_inst11.un1_dutycycle_53_13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_11_LC_5_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_11_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_11_LC_5_13_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_11_LC_5_13_0  (
            .in0(N__20876),
            .in1(N__21409),
            .in2(_gnd_net_),
            .in3(N__22345),
            .lcout(\b2v_inst11.G_6_i_a4_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_11_LC_5_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_11_LC_5_13_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_11_LC_5_13_1 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \b2v_inst11.dutycycle_11_LC_5_13_1  (
            .in0(N__19228),
            .in1(N__19239),
            .in2(N__21457),
            .in3(N__27303),
            .lcout(\b2v_inst11.dutycycleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34641),
            .ce(),
            .sr(N__24237));
    defparam \b2v_inst11.dutycycle_RNI_0_11_LC_5_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_11_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_11_LC_5_13_2 .LUT_INIT=16'b1111010100110101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_11_LC_5_13_2  (
            .in0(N__20875),
            .in1(N__19328),
            .in2(N__21441),
            .in3(N__22346),
            .lcout(),
            .ltout(\b2v_inst11.G_6_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_9_9_LC_5_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_9_9_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_9_9_LC_5_13_3 .LUT_INIT=16'b0000001000001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_9_9_LC_5_13_3  (
            .in0(N__20998),
            .in1(N__19270),
            .in2(N__19255),
            .in3(N__19252),
            .lcout(\b2v_inst11.un1_dutycycle_53_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI9JP25_11_LC_5_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI9JP25_11_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI9JP25_11_LC_5_13_4 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI9JP25_11_LC_5_13_4  (
            .in0(N__27302),
            .in1(N__21453),
            .in2(N__19240),
            .in3(N__19227),
            .lcout(\b2v_inst11.dutycycleZ0Z_7 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_11_LC_5_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_11_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_11_LC_5_13_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_11_LC_5_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19219),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_11 ),
            .ltout(\b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_9_LC_5_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_9_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_9_LC_5_13_6 .LUT_INIT=16'b1110111100001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_9_LC_5_13_6  (
            .in0(N__22774),
            .in1(N__20997),
            .in2(N__19216),
            .in3(N__22347),
            .lcout(\b2v_inst11.un1_dutycycle_53_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_11_LC_5_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_11_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_11_LC_5_13_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_11_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(N__22773),
            .in2(_gnd_net_),
            .in3(N__20874),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_0_LC_5_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_0_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_0_LC_5_14_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_0_LC_5_14_0  (
            .in0(N__25571),
            .in1(N__25364),
            .in2(N__28028),
            .in3(N__24512),
            .lcout(\b2v_inst11.g2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_12_LC_5_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_12_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_12_LC_5_14_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_12_LC_5_14_1  (
            .in0(N__19333),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21394),
            .lcout(\b2v_inst11.N_354 ),
            .ltout(\b2v_inst11.N_354_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_2_LC_5_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_2_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_2_LC_5_14_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_2_LC_5_14_2  (
            .in0(N__27417),
            .in1(_gnd_net_),
            .in2(N__19348),
            .in3(N__19429),
            .lcout(\b2v_inst11.N_360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_2_1_LC_5_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_2_1_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_2_1_LC_5_14_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.func_state_RNI_2_1_LC_5_14_3  (
            .in0(N__24511),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_3046_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_12_LC_5_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_12_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_12_LC_5_14_4 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_12_LC_5_14_4  (
            .in0(N__21395),
            .in1(N__19332),
            .in2(_gnd_net_),
            .in3(N__19430),
            .lcout(),
            .ltout(\b2v_inst11.g3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_0_LC_5_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_0_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_0_LC_5_14_5 .LUT_INIT=16'b1100110011111101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_0_LC_5_14_5  (
            .in0(N__19279),
            .in1(N__28832),
            .in2(N__19273),
            .in3(N__28141),
            .lcout(\b2v_inst11.g2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_4_LC_5_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_4_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_4_LC_5_14_6 .LUT_INIT=16'b0001000100010011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_4_LC_5_14_6  (
            .in0(N__26219),
            .in1(N__22772),
            .in2(N__28996),
            .in3(N__27999),
            .lcout(\b2v_inst11.N_14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNINJ641_0_5_LC_5_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNINJ641_0_5_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNINJ641_0_5_LC_5_14_7 .LUT_INIT=16'b1111000111111111;
    LogicCell40 \b2v_inst11.dutycycle_RNINJ641_0_5_LC_5_14_7  (
            .in0(N__28829),
            .in1(N__19264),
            .in2(N__27322),
            .in3(N__24314),
            .lcout(\b2v_inst11.dutycycle_RNINJ641_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_5_LC_5_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_5_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_5_LC_5_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_5_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__21492),
            .in2(_gnd_net_),
            .in3(N__23176),
            .lcout(\b2v_inst11.dutycycle_RNI_6Z0Z_5 ),
            .ltout(\b2v_inst11.dutycycle_RNI_6Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINJ641_2_1_LC_5_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINJ641_2_1_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINJ641_2_1_LC_5_15_1 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \b2v_inst11.func_state_RNINJ641_2_1_LC_5_15_1  (
            .in0(N__29239),
            .in1(N__21073),
            .in2(N__19258),
            .in3(N__21600),
            .lcout(\b2v_inst11.func_state_1_m2s2_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_3_1_LC_5_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_3_1_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_3_1_LC_5_15_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.func_state_RNI_3_1_LC_5_15_2  (
            .in0(N__21601),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24317),
            .lcout(\b2v_inst11.func_state_RNI_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIT4D71_1_LC_5_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIT4D71_1_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIT4D71_1_LC_5_15_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst11.count_clk_RNIT4D71_1_LC_5_15_3  (
            .in0(N__28559),
            .in1(N__24092),
            .in2(N__23428),
            .in3(N__19642),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIKOJB2_0_LC_5_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIKOJB2_0_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIKOJB2_0_LC_5_15_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \b2v_inst11.func_state_RNIKOJB2_0_LC_5_15_4  (
            .in0(N__22882),
            .in1(N__23242),
            .in2(N__19609),
            .in3(N__19606),
            .lcout(\b2v_inst11.N_122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_5_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_5_15_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_5_15_6  (
            .in0(N__28668),
            .in1(N__28253),
            .in2(_gnd_net_),
            .in3(N__28560),
            .lcout(\b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_LC_5_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_LC_5_15_7 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_LC_5_15_7  (
            .in0(N__21082),
            .in1(N__28142),
            .in2(N__27427),
            .in3(N__19428),
            .lcout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_0_0_LC_5_16_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_0_0_LC_5_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_0_0_LC_5_16_4 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a2_0_0_LC_5_16_4  (
            .in0(N__28219),
            .in1(N__28549),
            .in2(_gnd_net_),
            .in3(N__24301),
            .lcout(\b2v_inst11.un1_func_state25_6_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIC5UE2_1_LC_5_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIC5UE2_1_LC_5_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIC5UE2_1_LC_5_16_6 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \b2v_inst11.func_state_RNIC5UE2_1_LC_5_16_6  (
            .in0(N__19384),
            .in1(N__28548),
            .in2(N__24097),
            .in3(N__23376),
            .lcout(),
            .ltout(\b2v_inst11.func_state_1_m0_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIIVR84_0_LC_5_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIIVR84_0_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIIVR84_0_LC_5_16_7 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst11.func_state_RNIIVR84_0_LC_5_16_7  (
            .in0(N__23377),
            .in1(N__19372),
            .in2(N__19360),
            .in3(N__21475),
            .lcout(\b2v_inst11.func_state_1_m0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_1_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_1_0  (
            .in0(_gnd_net_),
            .in1(N__19858),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_1_0_),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_1_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_1_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_1_1  (
            .in0(_gnd_net_),
            .in1(N__19757),
            .in2(N__19714),
            .in3(N__19702),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_1_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_1_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_1_2  (
            .in0(_gnd_net_),
            .in1(N__19699),
            .in2(N__19762),
            .in3(N__19693),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_1_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_1_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_1_3  (
            .in0(_gnd_net_),
            .in1(N__20149),
            .in2(N__19690),
            .in3(N__19681),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_1_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_1_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_1_4  (
            .in0(_gnd_net_),
            .in1(N__19678),
            .in2(N__20157),
            .in3(N__19672),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_1_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_1_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_1_5  (
            .in0(N__19876),
            .in1(N__19761),
            .in2(N__19669),
            .in3(N__19660),
            .lcout(\b2v_inst11.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_1_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_1_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_1_6  (
            .in0(N__19657),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19651),
            .lcout(\b2v_inst11.mult1_un117_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un117_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_1_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_1_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19648),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_6_2_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_6_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_6_2_0  (
            .in0(_gnd_net_),
            .in1(N__20236),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_2_0_),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_6_2_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_6_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_6_2_1  (
            .in0(_gnd_net_),
            .in1(N__19793),
            .in2(N__19840),
            .in3(N__19645),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_6_2_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_6_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_6_2_2  (
            .in0(_gnd_net_),
            .in1(N__19828),
            .in2(N__19798),
            .in3(N__19822),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_6_2_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_6_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_6_2_3  (
            .in0(_gnd_net_),
            .in1(N__19877),
            .in2(N__19819),
            .in3(N__19810),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_6_2_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_6_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_6_2_4  (
            .in0(_gnd_net_),
            .in1(N__19807),
            .in2(N__19884),
            .in3(N__19801),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_6_2_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_6_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_6_2_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_6_2_5  (
            .in0(N__20263),
            .in1(N__19797),
            .in2(N__19783),
            .in3(N__19774),
            .lcout(\b2v_inst11.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_6_2_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_6_2_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_6_2_6  (
            .in0(N__19771),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19765),
            .lcout(\b2v_inst11.mult1_un124_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_6_2_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_6_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_6_2_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_6_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20153),
            .lcout(\b2v_inst11.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_6_3_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_6_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_6_3_0  (
            .in0(_gnd_net_),
            .in1(N__21744),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_6_3_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_6_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_6_3_1  (
            .in0(_gnd_net_),
            .in1(N__20218),
            .in2(N__19747),
            .in3(N__19738),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_6_3_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_6_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_6_3_2  (
            .in0(_gnd_net_),
            .in1(N__19735),
            .in2(N__19729),
            .in3(N__19981),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_6_3_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_6_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_6_3_3  (
            .in0(_gnd_net_),
            .in1(N__20264),
            .in2(N__19978),
            .in3(N__19966),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_6_3_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_6_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_6_3_4  (
            .in0(_gnd_net_),
            .in1(N__19963),
            .in2(N__20274),
            .in3(N__19957),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_6_3_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_6_3_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_6_3_5  (
            .in0(N__21796),
            .in1(N__19954),
            .in2(N__19948),
            .in3(N__19930),
            .lcout(\b2v_inst11.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_6_3_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_6_3_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_6_3_6  (
            .in0(_gnd_net_),
            .in1(N__19927),
            .in2(_gnd_net_),
            .in3(N__19921),
            .lcout(\b2v_inst11.mult1_un131_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un131_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_6_3_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_6_3_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_6_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19918),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_4_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19915),
            .lcout(\b2v_inst11.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_4_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19885),
            .lcout(\b2v_inst11.un85_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_4_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_4_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19854),
            .lcout(\b2v_inst11.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_6_4_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_6_4_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_6_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20275),
            .lcout(\b2v_inst11.un85_clk_100khz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_4_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_4_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20232),
            .lcout(\b2v_inst11.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_6_4_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_6_4_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_6_4_6  (
            .in0(N__20208),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_4_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_4_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20045),
            .lcout(\b2v_inst11.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_6_5_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_6_5_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20161),
            .lcout(\b2v_inst11.un85_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_6_5_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_5_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_5_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_6_5_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_6_5_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_6_5_2  (
            .in0(N__20080),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un85_clk_100khz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_6_5_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_6_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_6_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20037),
            .lcout(\b2v_inst11.mult1_un61_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_6_5_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_6_5_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_6_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20011),
            .lcout(\b2v_inst11.un85_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_5_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20442),
            .lcout(\b2v_inst11.mult1_un54_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_5_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_5_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20416),
            .lcout(\b2v_inst11.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_6_5_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_6_5_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_6_5_7  (
            .in0(N__20388),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un85_clk_100khz_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.delayed_vddq_pwrgd_LC_6_6_0 .C_ON=1'b0;
    defparam \b2v_inst16.delayed_vddq_pwrgd_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.delayed_vddq_pwrgd_LC_6_6_0 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \b2v_inst16.delayed_vddq_pwrgd_LC_6_6_0  (
            .in0(N__20629),
            .in1(N__20543),
            .in2(_gnd_net_),
            .in3(N__25077),
            .lcout(\b2v_inst16.delayed_vddq_pwrgdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34643),
            .ce(N__33684),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIPRCE_1_LC_6_6_1 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIPRCE_1_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIPRCE_1_LC_6_6_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \b2v_inst16.curr_state_RNIPRCE_1_LC_6_6_1  (
            .in0(N__20540),
            .in1(N__20358),
            .in2(N__20305),
            .in3(N__34058),
            .lcout(\b2v_inst16.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst16.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNI7SG01_1_LC_6_6_2 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNI7SG01_1_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNI7SG01_1_LC_6_6_2 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \b2v_inst16.curr_state_RNI7SG01_1_LC_6_6_2  (
            .in0(N__20628),
            .in1(_gnd_net_),
            .in2(N__20365),
            .in3(N__25073),
            .lcout(),
            .ltout(\b2v_inst16.curr_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_1_LC_6_6_3 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_1_LC_6_6_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.curr_state_1_LC_6_6_3 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \b2v_inst16.curr_state_1_LC_6_6_3  (
            .in0(N__20542),
            .in1(N__20554),
            .in2(N__20362),
            .in3(N__20359),
            .lcout(\b2v_inst16.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34643),
            .ce(N__33684),
            .sr(_gnd_net_));
    defparam \b2v_inst16.delayed_vddq_pwrgd_RNIJ10L1_LC_6_6_4 .C_ON=1'b0;
    defparam \b2v_inst16.delayed_vddq_pwrgd_RNIJ10L1_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.delayed_vddq_pwrgd_RNIJ10L1_LC_6_6_4 .LUT_INIT=16'b1110010011111111;
    LogicCell40 \b2v_inst16.delayed_vddq_pwrgd_RNIJ10L1_LC_6_6_4  (
            .in0(N__33715),
            .in1(N__20296),
            .in2(N__20548),
            .in3(N__25078),
            .lcout(b2v_inst16_un2_vpp_en_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_0_LC_6_6_5 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_0_LC_6_6_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.curr_state_0_LC_6_6_5 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \b2v_inst16.curr_state_0_LC_6_6_5  (
            .in0(N__20541),
            .in1(_gnd_net_),
            .in2(N__25085),
            .in3(N__20627),
            .lcout(\b2v_inst16.curr_state_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34643),
            .ce(N__33684),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNO_0_1_LC_6_6_6 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNO_0_1_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNO_0_1_LC_6_6_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst16.curr_state_RNO_0_1_LC_6_6_6  (
            .in0(N__34059),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20560),
            .lcout(\b2v_inst16.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIKEBL_1_LC_6_6_7 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIKEBL_1_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIKEBL_1_LC_6_6_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst16.curr_state_RNIKEBL_1_LC_6_6_7  (
            .in0(N__20544),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33714),
            .lcout(\b2v_inst16.count_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_0_LC_6_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_0_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_0_LC_6_7_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_0_LC_6_7_0  (
            .in0(N__28990),
            .in1(N__25595),
            .in2(_gnd_net_),
            .in3(N__25389),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_6_7_2 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_6_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(N__33081),
            .in2(_gnd_net_),
            .in3(N__20509),
            .lcout(\b2v_inst200.m11_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.DSW_PWROK_RNIUDI9_LC_6_7_4 .C_ON=1'b0;
    defparam \b2v_inst36.DSW_PWROK_RNIUDI9_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.DSW_PWROK_RNIUDI9_LC_6_7_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst36.DSW_PWROK_RNIUDI9_LC_6_7_4  (
            .in0(N__34060),
            .in1(N__22156),
            .in2(_gnd_net_),
            .in3(N__29998),
            .lcout(V105A_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_LC_6_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_LC_6_7_7 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_LC_6_7_7  (
            .in0(N__25390),
            .in1(N__26765),
            .in2(N__27436),
            .in3(N__28991),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_10_LC_6_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_10_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_10_LC_6_8_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_10_LC_6_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20572),
            .in3(N__22355),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_5_LC_6_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_5_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_5_LC_6_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_5_LC_6_8_7  (
            .in0(N__20596),
            .in1(N__21015),
            .in2(N__26782),
            .in3(N__28019),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_14_LC_6_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_14_LC_6_9_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_14_LC_6_9_1 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst11.dutycycle_14_LC_6_9_1  (
            .in0(N__27307),
            .in1(N__20701),
            .in2(N__21186),
            .in3(N__20692),
            .lcout(\b2v_inst11.dutycycleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34621),
            .ce(),
            .sr(N__24163));
    defparam \b2v_inst11.dutycycle_RNI2RTA8_14_LC_6_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI2RTA8_14_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI2RTA8_14_LC_6_9_2 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \b2v_inst11.dutycycle_RNI2RTA8_14_LC_6_9_2  (
            .in0(N__20700),
            .in1(N__20691),
            .in2(N__21187),
            .in3(N__27306),
            .lcout(\b2v_inst11.dutycycleZ0Z_13 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_15_LC_6_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_15_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_15_LC_6_9_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_15_LC_6_9_3  (
            .in0(N__21336),
            .in1(N__22309),
            .in2(N__20677),
            .in3(N__21153),
            .lcout(\b2v_inst11.un2_count_clk_17_0_a2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_10_LC_6_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_10_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_10_LC_6_9_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_10_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(N__22786),
            .in2(_gnd_net_),
            .in3(N__22308),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_50_a4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_7_LC_6_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_7_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_7_LC_6_9_6 .LUT_INIT=16'b0000000010101011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_7_LC_6_9_6  (
            .in0(N__26223),
            .in1(N__20668),
            .in2(N__20662),
            .in3(N__20658),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o2_LC_6_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o2_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o2_LC_6_10_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \b2v_inst11.un1_count_clk_1_sqmuxa_0_o2_LC_6_10_0  (
            .in0(N__28747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28307),
            .lcout(\b2v_inst11.N_158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst17.un4_vccio_en_0_a3_LC_6_10_3 .C_ON=1'b0;
    defparam \b2v_inst17.un4_vccio_en_0_a3_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst17.un4_vccio_en_0_a3_LC_6_10_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst17.un4_vccio_en_0_a3_LC_6_10_3  (
            .in0(N__20641),
            .in1(N__20626),
            .in2(_gnd_net_),
            .in3(N__29652),
            .lcout(VCCIO_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_10_LC_6_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_10_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_10_LC_6_10_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_10_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__26212),
            .in2(_gnd_net_),
            .in3(N__22287),
            .lcout(\b2v_inst11.un1_dutycycle_53_axb_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_LC_6_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_LC_6_10_5 .LUT_INIT=16'b1111100011100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_LC_6_10_5  (
            .in0(N__26211),
            .in1(N__22784),
            .in2(N__28962),
            .in3(N__24779),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_3 ),
            .ltout(\b2v_inst11.dutycycle_RNIZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_9_LC_6_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_9_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_9_LC_6_10_6 .LUT_INIT=16'b1011110101000010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_9_LC_6_10_6  (
            .in0(N__28015),
            .in1(N__20976),
            .in2(N__20581),
            .in3(N__20578),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI03R98_4_LC_6_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI03R98_4_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI03R98_4_LC_6_11_0 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI03R98_4_LC_6_11_0  (
            .in0(N__27231),
            .in1(N__21064),
            .in2(N__20733),
            .in3(N__20742),
            .lcout(\b2v_inst11.dutycycleZ0Z_8 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIAI7C4_4_LC_6_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIAI7C4_4_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIAI7C4_4_LC_6_11_1 .LUT_INIT=16'b0101111101001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIAI7C4_4_LC_6_11_1  (
            .in0(N__22585),
            .in1(N__27234),
            .in2(N__20761),
            .in3(N__28118),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNIAI7C4Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI3JFN6_4_LC_6_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI3JFN6_4_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI3JFN6_4_LC_6_11_2 .LUT_INIT=16'b0010001000101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI3JFN6_4_LC_6_11_2  (
            .in0(N__27618),
            .in1(N__27751),
            .in2(N__20758),
            .in3(N__22242),
            .lcout(\b2v_inst11.dutycycle_RNI3JFN6Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI3JFN6_0_LC_6_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI3JFN6_0_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI3JFN6_0_LC_6_11_3 .LUT_INIT=16'b1011001100000000;
    LogicCell40 \b2v_inst11.func_state_RNI3JFN6_0_LC_6_11_3  (
            .in0(N__22584),
            .in1(N__27750),
            .in2(N__20755),
            .in3(N__27617),
            .lcout(\b2v_inst11.func_state_RNI3JFN6Z0Z_0 ),
            .ltout(\b2v_inst11.func_state_RNI3JFN6Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_9_LC_6_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_9_LC_6_11_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_9_LC_6_11_4 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \b2v_inst11.dutycycle_9_LC_6_11_4  (
            .in0(N__27233),
            .in1(N__20910),
            .in2(N__20746),
            .in3(N__20719),
            .lcout(\b2v_inst11.dutycycleZ1Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34635),
            .ce(),
            .sr(N__24162));
    defparam \b2v_inst11.dutycycle_4_LC_6_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_4_LC_6_11_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_4_LC_6_11_6 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \b2v_inst11.dutycycle_4_LC_6_11_6  (
            .in0(N__27232),
            .in1(N__21063),
            .in2(N__20734),
            .in3(N__20743),
            .lcout(\b2v_inst11.dutycycleZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34635),
            .ce(),
            .sr(N__24162));
    defparam \b2v_inst11.dutycycle_RNIAI0A8_9_LC_6_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIAI0A8_9_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIAI0A8_9_LC_6_11_7 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \b2v_inst11.dutycycle_RNIAI0A8_9_LC_6_11_7  (
            .in0(N__20718),
            .in1(N__20710),
            .in2(N__20914),
            .in3(N__27230),
            .lcout(\b2v_inst11.dutycycleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI0KJ31_7_LC_6_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI0KJ31_7_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI0KJ31_7_LC_6_12_0 .LUT_INIT=16'b0011010101010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI0KJ31_7_LC_6_12_0  (
            .in0(N__20799),
            .in1(N__21043),
            .in2(N__26881),
            .in3(N__26960),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI0KJ31Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI74A23_7_LC_6_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI74A23_7_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI74A23_7_LC_6_12_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \b2v_inst11.dutycycle_RNI74A23_7_LC_6_12_1  (
            .in0(N__27275),
            .in1(_gnd_net_),
            .in2(N__20704),
            .in3(N__20785),
            .lcout(\b2v_inst11.dutycycle_RNI74A23Z0Z_7 ),
            .ltout(\b2v_inst11.dutycycle_RNI74A23Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIF271B_7_LC_6_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIF271B_7_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIF271B_7_LC_6_12_2 .LUT_INIT=16'b0010111000001111;
    LogicCell40 \b2v_inst11.dutycycle_RNIF271B_7_LC_6_12_2  (
            .in0(N__20797),
            .in1(N__20839),
            .in2(N__20842),
            .in3(N__27752),
            .lcout(\b2v_inst11.dutycycleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI7UR36_0_LC_6_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI7UR36_0_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI7UR36_0_LC_6_12_3 .LUT_INIT=16'b0000000000011111;
    LogicCell40 \b2v_inst11.func_state_RNI7UR36_0_LC_6_12_3  (
            .in0(N__27274),
            .in1(N__28140),
            .in2(N__20809),
            .in3(N__22227),
            .lcout(\b2v_inst11.dutycycle_e_1_7 ),
            .ltout(\b2v_inst11.dutycycle_e_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_7_LC_6_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_7_LC_6_12_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_7_LC_6_12_4 .LUT_INIT=16'b0011101000110011;
    LogicCell40 \b2v_inst11.dutycycle_7_LC_6_12_4  (
            .in0(N__20800),
            .in1(N__20833),
            .in2(N__20827),
            .in3(N__27753),
            .lcout(\b2v_inst11.dutycycleZ1Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34642),
            .ce(),
            .sr(N__24210));
    defparam \b2v_inst11.dutycycle_RNI25OT3_7_LC_6_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI25OT3_7_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI25OT3_7_LC_6_12_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.dutycycle_RNI25OT3_7_LC_6_12_5  (
            .in0(N__24484),
            .in1(N__20824),
            .in2(_gnd_net_),
            .in3(N__26680),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI25OT3Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIGALV4_0_LC_6_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIGALV4_0_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIGALV4_0_LC_6_12_6 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \b2v_inst11.func_state_RNIGALV4_0_LC_6_12_6  (
            .in0(N__23290),
            .in1(N__26210),
            .in2(N__20812),
            .in3(N__23121),
            .lcout(\b2v_inst11.func_state_RNIGALV4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIGSFQ_7_LC_6_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIGSFQ_7_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIGSFQ_7_LC_6_12_7 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \b2v_inst11.dutycycle_RNIGSFQ_7_LC_6_12_7  (
            .in0(N__26959),
            .in1(N__20798),
            .in2(_gnd_net_),
            .in3(N__26873),
            .lcout(\b2v_inst11.dutycycle_RNIGSFQZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_0_LC_6_13_0 .C_ON=1'b1;
    defparam \b2v_inst11.dutycycle_RNI_2_0_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_0_LC_6_13_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_0_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(N__25548),
            .in2(_gnd_net_),
            .in3(N__25383),
            .lcout(\b2v_inst11.g0_2_3 ),
            .ltout(),
            .carryin(bfn_6_13_0_),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_0_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_6_13_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_6_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(N__29217),
            .in2(N__25392),
            .in3(N__20779),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_0_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDU8_LC_6_13_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDU8_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDU8_LC_6_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDU8_LC_6_13_2  (
            .in0(_gnd_net_),
            .in1(N__29237),
            .in2(N__27413),
            .in3(N__20764),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_1_c_RNIBDUZ0Z8 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_1 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_6_13_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_6_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_6_13_3  (
            .in0(_gnd_net_),
            .in1(N__29216),
            .in2(N__24816),
            .in3(N__21067),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_2 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_6_13_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_6_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_6_13_4  (
            .in0(_gnd_net_),
            .in1(N__29238),
            .in2(N__28992),
            .in3(N__21052),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_3 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNI578D1_LC_6_13_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNI578D1_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNI578D1_LC_6_13_5 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_4_c_RNI578D1_LC_6_13_5  (
            .in0(N__27235),
            .in1(N__29222),
            .in2(N__26781),
            .in3(N__21049),
            .lcout(\b2v_inst11.g1_4_0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_4 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNI_LC_6_13_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNI_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNI_LC_6_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_5_c_RNI_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(N__27956),
            .in2(N__29250),
            .in3(N__21046),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_5_c_RNIZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_5_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_6_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_6_13_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_6_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_6_13_7  (
            .in0(_gnd_net_),
            .in1(N__29221),
            .in2(N__26224),
            .in3(N__21037),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_6_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHP49_LC_6_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHP49_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHP49_LC_6_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHP49_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(N__22785),
            .in2(N__29247),
            .in3(N__21019),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHPZ0Z49 ),
            .ltout(),
            .carryin(bfn_6_14_0_),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIR59_LC_6_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIR59_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIR59_LC_6_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIR59_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(N__29214),
            .in2(N__21016),
            .in3(N__20899),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_8_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_9_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJT69_LC_6_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJT69_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJT69_LC_6_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJT69_LC_6_14_2  (
            .in0(_gnd_net_),
            .in1(N__22349),
            .in2(N__29248),
            .in3(N__20896),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJTZ0Z69 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_9_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNP5_LC_6_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNP5_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNP5_LC_6_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNP5_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(N__29200),
            .in2(N__20893),
            .in3(N__21445),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNPZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_10 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQ5_LC_6_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQ5_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQ5_LC_6_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQ5_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(N__21435),
            .in2(N__29246),
            .in3(N__21340),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_11 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_6_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_6_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_6_14_5  (
            .in0(_gnd_net_),
            .in1(N__29201),
            .in2(N__21337),
            .in3(N__21250),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_12 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_6_14_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_6_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(N__21247),
            .in2(N__29249),
            .in3(N__21166),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_13 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_6_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_6_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_6_14_7  (
            .in0(N__21163),
            .in1(N__29215),
            .in2(_gnd_net_),
            .in3(N__21109),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_5_LC_6_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_5_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_5_LC_6_15_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_5_LC_6_15_0  (
            .in0(N__25346),
            .in1(N__26780),
            .in2(N__25570),
            .in3(N__27912),
            .lcout(\b2v_inst11.dutycycle_RNI_5Z0Z_5 ),
            .ltout(\b2v_inst11.dutycycle_RNI_5Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_0_LC_6_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_0_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_0_LC_6_15_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst11.func_state_RNI_0_LC_6_15_1  (
            .in0(N__23110),
            .in1(N__24279),
            .in2(N__21085),
            .in3(N__23204),
            .lcout(\b2v_inst11.N_156 ),
            .ltout(\b2v_inst11.N_156_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_2_LC_6_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_2_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_2_LC_6_15_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_2_LC_6_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21076),
            .in3(N__23174),
            .lcout(\b2v_inst11.N_418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINJ641_1_1_LC_6_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINJ641_1_1_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINJ641_1_1_LC_6_15_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst11.func_state_RNINJ641_1_1_LC_6_15_3  (
            .in0(N__24722),
            .in1(N__23238),
            .in2(_gnd_net_),
            .in3(N__24278),
            .lcout(\b2v_inst11.N_331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_6_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_6_15_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_6_15_4  (
            .in0(N__23205),
            .in1(N__29235),
            .in2(N__23056),
            .in3(N__23175),
            .lcout(\b2v_inst11.un1_func_state25_6_0_o_N_307_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_1_LC_6_15_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_1_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_1_LC_6_15_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst11.func_state_RNI_1_LC_6_15_5  (
            .in0(_gnd_net_),
            .in1(N__28454),
            .in2(_gnd_net_),
            .in3(N__24277),
            .lcout(\b2v_inst11.N_169 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIQQRO_5_LC_6_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIQQRO_5_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIQQRO_5_LC_6_15_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.dutycycle_RNIQQRO_5_LC_6_15_6  (
            .in0(N__21493),
            .in1(N__24854),
            .in2(N__23184),
            .in3(N__25065),
            .lcout(),
            .ltout(\b2v_inst11.N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI8PGM6_5_LC_6_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI8PGM6_5_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI8PGM6_5_LC_6_15_7 .LUT_INIT=16'b0101010101011101;
    LogicCell40 \b2v_inst11.dutycycle_RNI8PGM6_5_LC_6_15_7  (
            .in0(N__27776),
            .in1(N__29023),
            .in2(N__21481),
            .in3(N__23455),
            .lcout(\b2v_inst11.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_0_0_LC_6_16_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_0_0_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_0_0_LC_6_16_0 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \b2v_inst11.func_state_RNI_0_0_LC_6_16_0  (
            .in0(_gnd_net_),
            .in1(N__23109),
            .in2(N__23206),
            .in3(N__23183),
            .lcout(\b2v_inst11.func_state_RNI_0Z0Z_0 ),
            .ltout(\b2v_inst11.func_state_RNI_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINJ641_0_0_LC_6_16_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINJ641_0_0_LC_6_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINJ641_0_0_LC_6_16_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.func_state_RNINJ641_0_0_LC_6_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21478),
            .in3(N__24723),
            .lcout(\b2v_inst11.func_state_RNINJ641_0Z0Z_0 ),
            .ltout(\b2v_inst11.func_state_RNINJ641_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIQCBN4_9_LC_6_16_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIQCBN4_9_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIQCBN4_9_LC_6_16_2 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \b2v_inst11.count_off_RNIQCBN4_9_LC_6_16_2  (
            .in0(N__21463),
            .in1(N__27772),
            .in2(N__21469),
            .in3(N__23308),
            .lcout(\b2v_inst11.count_off_RNIQCBN4Z0Z_9 ),
            .ltout(\b2v_inst11.count_off_RNIQCBN4Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDINH9_0_LC_6_16_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDINH9_0_LC_6_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDINH9_0_LC_6_16_3 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \b2v_inst11.func_state_RNIDINH9_0_LC_6_16_3  (
            .in0(N__21547),
            .in1(N__21526),
            .in2(N__21466),
            .in3(N__25066),
            .lcout(\b2v_inst11.func_state_RNIDINH9Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI7J1P_1_LC_6_16_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI7J1P_1_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI7J1P_1_LC_6_16_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \b2v_inst11.func_state_RNI7J1P_1_LC_6_16_4  (
            .in0(N__28674),
            .in1(N__34006),
            .in2(N__28308),
            .in3(N__21598),
            .lcout(\b2v_inst11.N_333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIQBAL3_1_LC_6_16_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIQBAL3_1_LC_6_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIQBAL3_1_LC_6_16_5 .LUT_INIT=16'b1100111111101111;
    LogicCell40 \b2v_inst11.func_state_RNIQBAL3_1_LC_6_16_5  (
            .in0(N__21599),
            .in1(N__21553),
            .in2(N__27781),
            .in3(N__24096),
            .lcout(\b2v_inst11.N_73 ),
            .ltout(\b2v_inst11.N_73_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI673P9_0_LC_6_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI673P9_0_LC_6_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI673P9_0_LC_6_16_6 .LUT_INIT=16'b0000010001010100;
    LogicCell40 \b2v_inst11.func_state_RNI673P9_0_LC_6_16_6  (
            .in0(N__25067),
            .in1(N__21541),
            .in2(N__21535),
            .in3(N__21532),
            .lcout(\b2v_inst11.func_state_RNI673P9Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIPAG14_0_LC_6_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIPAG14_0_LC_6_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIPAG14_0_LC_6_16_7 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \b2v_inst11.func_state_RNIPAG14_0_LC_6_16_7  (
            .in0(N__23467),
            .in1(N__23212),
            .in2(N__23427),
            .in3(N__24724),
            .lcout(\b2v_inst11.func_state_1_m0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_7_2_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_7_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_7_2_0  (
            .in0(_gnd_net_),
            .in1(N__23953),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_2_0_),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_7_2_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_7_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_7_2_1  (
            .in0(_gnd_net_),
            .in1(N__21713),
            .in2(N__21757),
            .in3(N__21520),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_7_2_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_7_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_7_2_2  (
            .in0(_gnd_net_),
            .in1(N__21703),
            .in2(N__21718),
            .in3(N__21517),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_7_2_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_7_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_7_2_3  (
            .in0(_gnd_net_),
            .in1(N__21855),
            .in2(N__21685),
            .in3(N__21514),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_7_2_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_7_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_7_2_4  (
            .in0(_gnd_net_),
            .in1(N__21661),
            .in2(N__21859),
            .in3(N__21511),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_7_2_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_7_2_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_7_2_5  (
            .in0(N__23709),
            .in1(N__21717),
            .in2(N__21646),
            .in3(N__21508),
            .lcout(\b2v_inst11.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_7_2_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_7_2_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_7_2_6  (
            .in0(N__21610),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21721),
            .lcout(\b2v_inst11.mult1_un145_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_7_2_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_7_2_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_7_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21854),
            .lcout(\b2v_inst11.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_7_3_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_7_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_7_3_0  (
            .in0(_gnd_net_),
            .in1(N__21778),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_3_0_),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_7_3_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_7_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_7_3_1  (
            .in0(_gnd_net_),
            .in1(N__21994),
            .in2(N__21627),
            .in3(N__21697),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_7_3_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_7_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_7_3_2  (
            .in0(_gnd_net_),
            .in1(N__21623),
            .in2(N__21694),
            .in3(N__21676),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_7_3_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_7_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_7_3_3  (
            .in0(_gnd_net_),
            .in1(N__21797),
            .in2(N__21673),
            .in3(N__21655),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_7_3_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_7_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_7_3_4  (
            .in0(_gnd_net_),
            .in1(N__21652),
            .in2(N__21802),
            .in3(N__21637),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_7_3_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_7_3_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_7_3_5  (
            .in0(N__21853),
            .in1(N__21634),
            .in2(N__21628),
            .in3(N__21604),
            .lcout(\b2v_inst11.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_7_3_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_7_3_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_7_3_6  (
            .in0(N__21868),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21862),
            .lcout(\b2v_inst11.mult1_un138_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un138_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_7_3_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_7_3_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_7_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21838),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un85_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_7_4_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_7_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_7_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23718),
            .lcout(\b2v_inst11.un85_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_7_4_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_7_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_7_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23619),
            .lcout(\b2v_inst11.un85_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_4_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_4_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_4_2  (
            .in0(N__23949),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_7_4_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_7_4_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_7_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25465),
            .lcout(\b2v_inst11.un85_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_7_4_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_7_4_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_7_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21835),
            .lcout(\b2v_inst11.un85_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_7_4_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_7_4_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_7_4_5  (
            .in0(N__21801),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un85_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_4_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_4_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21774),
            .lcout(\b2v_inst11.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_7_4_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_7_4_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_7_4_7  (
            .in0(N__21745),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_7_5_0 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_7_5_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_7_5_0  (
            .in0(N__26536),
            .in1(N__25408),
            .in2(N__21988),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un1_count_cry_0_i ),
            .ltout(),
            .carryin(bfn_7_5_0_),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_7_5_1 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_7_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_7_5_1  (
            .in0(_gnd_net_),
            .in1(N__21964),
            .in2(N__21973),
            .in3(N__26563),
            .lcout(\b2v_inst11.N_5647_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_0 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_7_5_2 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_7_5_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_7_5_2  (
            .in0(N__25920),
            .in1(N__21958),
            .in2(N__21952),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5648_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_1 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_7_5_3 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_7_5_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_7_5_3  (
            .in0(N__25624),
            .in1(N__21943),
            .in2(N__21937),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5649_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_2 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_7_5_4 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_7_5_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_7_5_4  (
            .in0(_gnd_net_),
            .in1(N__21913),
            .in2(N__21925),
            .in3(N__26029),
            .lcout(\b2v_inst11.N_5650_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_3 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_7_5_5 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_7_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_7_5_5  (
            .in0(_gnd_net_),
            .in1(N__21898),
            .in2(N__21907),
            .in3(N__25987),
            .lcout(\b2v_inst11.N_5651_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_4 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_7_5_6 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_7_5_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_7_5_6  (
            .in0(N__25758),
            .in1(N__21892),
            .in2(N__21886),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5652_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_5 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_7_5_7 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_7_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_7_5_7  (
            .in0(_gnd_net_),
            .in1(N__22120),
            .in2(N__21877),
            .in3(N__25894),
            .lcout(\b2v_inst11.N_5653_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_6 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_7_6_0 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_7_6_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_7_6_0  (
            .in0(N__26407),
            .in1(N__22105),
            .in2(N__22114),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5654_i ),
            .ltout(),
            .carryin(bfn_7_6_0_),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_7_6_1 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_7_6_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_7_6_1  (
            .in0(N__26364),
            .in1(N__22099),
            .in2(N__22087),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5655_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_8 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_7_6_2 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_7_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__22069),
            .in2(N__22078),
            .in3(N__25819),
            .lcout(\b2v_inst11.N_5656_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_9 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_7_6_3 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_7_6_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_7_6_3  (
            .in0(N__25846),
            .in1(N__22063),
            .in2(N__22051),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5657_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_10 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_7_6_4 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_7_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(N__22030),
            .in2(N__22042),
            .in3(N__25787),
            .lcout(\b2v_inst11.N_5658_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_11 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_7_6_5 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_7_6_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_7_6_5  (
            .in0(N__26071),
            .in1(N__22024),
            .in2(N__22018),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5659_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_12 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_7_6_6 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_7_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(N__22000),
            .in2(N__22009),
            .in3(N__25731),
            .lcout(\b2v_inst11.N_5660_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_13 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_7_6_7 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_7_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_7_6_7  (
            .in0(_gnd_net_),
            .in1(N__22165),
            .in2(N__22174),
            .in3(N__25866),
            .lcout(\b2v_inst11.N_5661_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_14 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_15_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_7_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_7_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22159),
            .lcout(\b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_0_LC_7_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_0_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_0_LC_7_7_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst11.count_RNI_0_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__26531),
            .in2(_gnd_net_),
            .in3(N__26440),
            .lcout(\b2v_inst11.count_RNI_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_7_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_7_7_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_7_7_3  (
            .in0(N__25701),
            .in1(N__25656),
            .in2(_gnd_net_),
            .in3(N__26638),
            .lcout(\b2v_inst11.curr_state_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNI8TT2_0_LC_7_7_4 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI8TT2_0_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI8TT2_0_LC_7_7_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst36.curr_state_RNI8TT2_0_LC_7_7_4  (
            .in0(N__30402),
            .in1(N__30306),
            .in2(_gnd_net_),
            .in3(N__30358),
            .lcout(\b2v_inst36.curr_state_RNI8TT2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNICRLO_LC_7_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNICRLO_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNICRLO_LC_7_8_0 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_15_c_RNICRLO_LC_7_8_0  (
            .in0(N__25655),
            .in1(N__22126),
            .in2(N__26649),
            .in3(N__33718),
            .lcout(),
            .ltout(\b2v_inst11.pwm_out_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.pwm_out_RNIEV5S_LC_7_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_RNIEV5S_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.pwm_out_RNIEV5S_LC_7_8_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \b2v_inst11.pwm_out_RNIEV5S_LC_7_8_1  (
            .in0(_gnd_net_),
            .in1(N__26611),
            .in2(N__22147),
            .in3(N__25654),
            .lcout(PWRBTN_LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNIOCA3_0_0_LC_7_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_0_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_0_LC_7_8_2 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \b2v_inst11.curr_state_RNIOCA3_0_0_LC_7_8_2  (
            .in0(N__25653),
            .in1(_gnd_net_),
            .in2(N__34085),
            .in3(N__25700),
            .lcout(\b2v_inst11.pwm_out_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_0_LC_7_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_0_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.curr_state_0_LC_7_8_3 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \b2v_inst11.curr_state_0_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(N__26642),
            .in2(N__25702),
            .in3(N__25652),
            .lcout(\b2v_inst11.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34637),
            .ce(N__33679),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNIJK34_0_LC_7_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNIJK34_0_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNIJK34_0_LC_7_8_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.curr_state_RNIJK34_0_LC_7_8_5  (
            .in0(N__22432),
            .in1(N__34036),
            .in2(_gnd_net_),
            .in3(N__22426),
            .lcout(\b2v_inst11.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst11.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNIOCA3_0_LC_7_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_LC_7_8_6 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \b2v_inst11.curr_state_RNIOCA3_0_LC_7_8_6  (
            .in0(N__34037),
            .in1(_gnd_net_),
            .in2(N__22420),
            .in3(N__25696),
            .lcout(\b2v_inst11.count_0_sqmuxa_i ),
            .ltout(\b2v_inst11.count_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_0_LC_7_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_0_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_0_LC_7_8_7 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \b2v_inst11.count_0_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22417),
            .in3(N__26535),
            .lcout(\b2v_inst11.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34637),
            .ce(N__33679),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_4_LC_7_9_0 .C_ON=1'b0;
    defparam \b2v_inst20.counter_4_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_4_LC_7_9_0 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \b2v_inst20.counter_4_LC_7_9_0  (
            .in0(N__31005),
            .in1(N__30985),
            .in2(_gnd_net_),
            .in3(N__26878),
            .lcout(\b2v_inst20.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34625),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_3_LC_7_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_3_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_3_LC_7_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_3_LC_7_9_2  (
            .in0(N__26236),
            .in1(N__24818),
            .in2(N__25596),
            .in3(N__25391),
            .lcout(\b2v_inst11.g0_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIJU083_0_LC_7_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIJU083_0_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIJU083_0_LC_7_9_4 .LUT_INIT=16'b1010111010111111;
    LogicCell40 \b2v_inst11.func_state_RNIJU083_0_LC_7_9_4  (
            .in0(N__23251),
            .in1(N__24464),
            .in2(N__27090),
            .in3(N__27021),
            .lcout(\b2v_inst11.func_state_RNIJU083Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_3_LC_7_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_3_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_3_LC_7_9_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_3_LC_7_9_7  (
            .in0(N__24817),
            .in1(N__28994),
            .in2(_gnd_net_),
            .in3(N__26235),
            .lcout(\b2v_inst11.N_349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIAI7C4_10_LC_7_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIAI7C4_10_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIAI7C4_10_LC_7_10_0 .LUT_INIT=16'b0101010101000000;
    LogicCell40 \b2v_inst11.dutycycle_RNIAI7C4_10_LC_7_10_0  (
            .in0(N__22244),
            .in1(N__22310),
            .in2(N__22577),
            .in3(N__22401),
            .lcout(\b2v_inst11.dutycycle_RNIAI7C4Z0Z_10 ),
            .ltout(\b2v_inst11.dutycycle_RNIAI7C4Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIP8IN8_10_LC_7_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIP8IN8_10_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIP8IN8_10_LC_7_10_1 .LUT_INIT=16'b0011101100110001;
    LogicCell40 \b2v_inst11.dutycycle_RNIP8IN8_10_LC_7_10_1  (
            .in0(N__27693),
            .in1(N__22513),
            .in2(N__22366),
            .in3(N__22493),
            .lcout(\b2v_inst11.dutycycleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNINJ641_3_LC_7_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNINJ641_3_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNINJ641_3_LC_7_10_3 .LUT_INIT=16'b1111111100001110;
    LogicCell40 \b2v_inst11.dutycycle_RNINJ641_3_LC_7_10_3  (
            .in0(N__27257),
            .in1(N__28153),
            .in2(N__24812),
            .in3(N__22243),
            .lcout(),
            .ltout(\b2v_inst11.un1_clk_100khz_43_and_i_o2_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI3JFN6_3_LC_7_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI3JFN6_3_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI3JFN6_3_LC_7_10_4 .LUT_INIT=16'b0011101100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI3JFN6_3_LC_7_10_4  (
            .in0(N__22553),
            .in1(N__27692),
            .in2(N__22528),
            .in3(N__27535),
            .lcout(\b2v_inst11.dutycycle_e_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.N_221_i_LC_7_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.N_221_i_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.N_221_i_LC_7_10_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst11.N_221_i_LC_7_10_5  (
            .in0(N__29071),
            .in1(N__29314),
            .in2(N__34091),
            .in3(N__28591),
            .lcout(\b2v_inst11.N_221_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI4I3C2_10_LC_7_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI4I3C2_10_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI4I3C2_10_LC_7_10_6 .LUT_INIT=16'b1101110100001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI4I3C2_10_LC_7_10_6  (
            .in0(N__22525),
            .in1(N__27258),
            .in2(N__22498),
            .in3(N__27536),
            .lcout(\b2v_inst11.dutycycle_RNI4I3C2Z0Z_10 ),
            .ltout(\b2v_inst11.dutycycle_RNI4I3C2Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_10_LC_7_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_10_LC_7_10_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_10_LC_7_10_7 .LUT_INIT=16'b0000111110001101;
    LogicCell40 \b2v_inst11.dutycycle_10_LC_7_10_7  (
            .in0(N__27694),
            .in1(N__22497),
            .in2(N__22507),
            .in3(N__22504),
            .lcout(\b2v_inst11.dutycycleZ1Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34636),
            .ce(),
            .sr(N__24160));
    defparam \b2v_inst11.dutycycle_RNI_1_5_LC_7_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_5_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_5_LC_7_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_5_LC_7_11_0  (
            .in0(N__22763),
            .in1(N__22831),
            .in2(N__26757),
            .in3(N__28956),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_3_LC_7_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_3_LC_7_11_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_3_LC_7_11_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \b2v_inst11.dutycycle_3_LC_7_11_1  (
            .in0(N__27229),
            .in1(N__22800),
            .in2(N__22813),
            .in3(N__22825),
            .lcout(\b2v_inst11.dutycycleZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34644),
            .ce(),
            .sr(N__24161));
    defparam \b2v_inst11.dutycycle_RNI_4_3_LC_7_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_3_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_3_LC_7_11_2 .LUT_INIT=16'b0000001100111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_3_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__25379),
            .in2(N__24807),
            .in3(N__27987),
            .lcout(),
            .ltout(\b2v_inst11.d_i3_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_5_LC_7_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_5_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_5_LC_7_11_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_5_LC_7_11_3  (
            .in0(N__23977),
            .in1(N__22446),
            .in2(N__22468),
            .in3(N__26732),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_3_LC_7_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_3_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_3_LC_7_11_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_3_LC_7_11_4  (
            .in0(N__26180),
            .in1(_gnd_net_),
            .in2(N__24808),
            .in3(N__28955),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_3_LC_7_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_3_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_3_LC_7_11_5 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_3_LC_7_11_5  (
            .in0(N__28954),
            .in1(N__24782),
            .in2(_gnd_net_),
            .in3(N__26179),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIUVP98_3_LC_7_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIUVP98_3_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIUVP98_3_LC_7_11_6 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \b2v_inst11.dutycycle_RNIUVP98_3_LC_7_11_6  (
            .in0(N__22824),
            .in1(N__22809),
            .in2(N__22801),
            .in3(N__27228),
            .lcout(\b2v_inst11.dutycycleZ0Z_6 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_3_LC_7_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_3_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_3_LC_7_11_7 .LUT_INIT=16'b0001010101010111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_3_LC_7_11_7  (
            .in0(N__28953),
            .in1(N__26178),
            .in2(N__22789),
            .in3(N__22762),
            .lcout(\b2v_inst11.dutycycle_RNI_5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINJ641_0_1_LC_7_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINJ641_0_1_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINJ641_0_1_LC_7_12_0 .LUT_INIT=16'b1111111100011101;
    LogicCell40 \b2v_inst11.func_state_RNINJ641_0_1_LC_7_12_0  (
            .in0(N__27029),
            .in1(N__24482),
            .in2(N__27109),
            .in3(N__22912),
            .lcout(\b2v_inst11.func_state_RNINJ641_0Z0Z_1 ),
            .ltout(\b2v_inst11.func_state_RNINJ641_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNINJ641_2_LC_7_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNINJ641_2_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNINJ641_2_LC_7_12_1 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNINJ641_2_LC_7_12_1  (
            .in0(N__27389),
            .in1(N__24393),
            .in2(N__22636),
            .in3(N__24315),
            .lcout(\b2v_inst11.g0_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_1_LC_7_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_1_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_1_LC_7_12_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_0_o3_1_1_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__28739),
            .in2(_gnd_net_),
            .in3(N__28322),
            .lcout(\b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1 ),
            .ltout(\b2v_inst11.dutycycle_1_0_iv_0_o3_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_7_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_7_12_3 .LUT_INIT=16'b0010111101111111;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_7_12_3  (
            .in0(N__24483),
            .in1(N__27103),
            .in2(N__22633),
            .in3(N__27030),
            .lcout(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_6_LC_7_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_6_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_6_LC_7_12_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_6_LC_7_12_4  (
            .in0(N__22630),
            .in1(N__22624),
            .in2(N__28013),
            .in3(N__28168),
            .lcout(\b2v_inst11.un1_dutycycle_164_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_4_LC_7_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_4_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_4_LC_7_12_5 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_4_LC_7_12_5  (
            .in0(N__28930),
            .in1(N__26187),
            .in2(_gnd_net_),
            .in3(N__27965),
            .lcout(\b2v_inst11.g0_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_7_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_7_12_6 .LUT_INIT=16'b0010010111111111;
    LogicCell40 \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_LC_7_12_6  (
            .in0(N__28746),
            .in1(N__33994),
            .in2(N__28345),
            .in3(N__29085),
            .lcout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_oZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIF6NL_1_LC_7_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIF6NL_1_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIF6NL_1_LC_7_12_7 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \b2v_inst11.func_state_RNIF6NL_1_LC_7_12_7  (
            .in0(N__28740),
            .in1(_gnd_net_),
            .in2(N__28343),
            .in3(N__28395),
            .lcout(\b2v_inst11.un1_clk_100khz_2_i_o3_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_LC_7_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_1_LC_7_13_0 .LUT_INIT=16'b0111111100100000;
    LogicCell40 \b2v_inst11.dutycycle_1_LC_7_13_0  (
            .in0(N__27547),
            .in1(N__22900),
            .in2(N__24544),
            .in3(N__22894),
            .lcout(\b2v_inst11.dutycycleZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34653),
            .ce(),
            .sr(N__24187));
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNI1V3D1_LC_7_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNI1V3D1_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNI1V3D1_LC_7_13_1 .LUT_INIT=16'b1111101011110011;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_0_c_RNI1V3D1_LC_7_13_1  (
            .in0(N__23113),
            .in1(N__22906),
            .in2(N__23053),
            .in3(N__28405),
            .lcout(\b2v_inst11.dutycycle_1_0_1 ),
            .ltout(\b2v_inst11.dutycycle_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIP4GA6_1_LC_7_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIP4GA6_1_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIP4GA6_1_LC_7_13_2 .LUT_INIT=16'b0100111011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIP4GA6_1_LC_7_13_2  (
            .in0(N__27546),
            .in1(N__22893),
            .in2(N__22885),
            .in3(N__24537),
            .lcout(\b2v_inst11.dutycycle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_1_0_LC_7_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_1_0_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_1_0_LC_7_13_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.func_state_RNI_1_0_LC_7_13_3  (
            .in0(N__23112),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28404),
            .lcout(\b2v_inst11.func_state_RNI_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_0_1_LC_7_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_0_1_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_0_1_LC_7_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.func_state_RNI_0_1_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__28403),
            .in2(_gnd_net_),
            .in3(N__23422),
            .lcout(\b2v_inst11.func_state_RNI_0Z0Z_1 ),
            .ltout(\b2v_inst11.func_state_RNI_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_3_0_LC_7_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_3_0_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_3_0_LC_7_13_6 .LUT_INIT=16'b0000000100001111;
    LogicCell40 \b2v_inst11.func_state_RNI_3_0_LC_7_13_6  (
            .in0(N__23423),
            .in1(N__28429),
            .in2(N__22852),
            .in3(N__23111),
            .lcout(),
            .ltout(\b2v_inst11.un1_func_state25_4_i_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIOJI01_0_LC_7_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIOJI01_0_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIOJI01_0_LC_7_13_7 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \b2v_inst11.func_state_RNIOJI01_0_LC_7_13_7  (
            .in0(N__28577),
            .in1(_gnd_net_),
            .in2(N__22849),
            .in3(N__29660),
            .lcout(\b2v_inst11.N_321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_6_LC_7_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_6_LC_7_14_0 .SEQ_MODE=4'b1011;
    defparam \b2v_inst11.dutycycle_6_LC_7_14_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \b2v_inst11.dutycycle_6_LC_7_14_0  (
            .in0(N__22984),
            .in1(N__22990),
            .in2(N__27620),
            .in3(N__22972),
            .lcout(\b2v_inst11.dutycycle_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34659),
            .ce(),
            .sr(N__24214));
    defparam \b2v_inst11.func_state_RNINJ641_0_LC_7_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINJ641_0_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINJ641_0_LC_7_14_1 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \b2v_inst11.func_state_RNINJ641_0_LC_7_14_1  (
            .in0(N__25549),
            .in1(N__28413),
            .in2(N__23055),
            .in3(N__23114),
            .lcout(\b2v_inst11.dutycycle_1_0_0 ),
            .ltout(\b2v_inst11.dutycycle_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIEOI16_0_LC_7_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIEOI16_0_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIEOI16_0_LC_7_14_2 .LUT_INIT=16'b0111111100001000;
    LogicCell40 \b2v_inst11.dutycycle_RNIEOI16_0_LC_7_14_2  (
            .in0(N__27606),
            .in1(N__22960),
            .in2(N__23005),
            .in3(N__22941),
            .lcout(\b2v_inst11.dutycycleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIKOJB2_LC_7_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIKOJB2_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIKOJB2_LC_7_14_4 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIKOJB2_LC_7_14_4  (
            .in0(N__24109),
            .in1(N__27262),
            .in2(N__26965),
            .in3(N__23002),
            .lcout(\b2v_inst11.g1 ),
            .ltout(\b2v_inst11.g1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIBDKS9_6_LC_7_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIBDKS9_6_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIBDKS9_6_LC_7_14_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIBDKS9_6_LC_7_14_5  (
            .in0(N__27603),
            .in1(N__22983),
            .in2(N__22975),
            .in3(N__22971),
            .lcout(\b2v_inst11.dutycycleZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIEFS24_0_LC_7_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIEFS24_0_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIEFS24_0_LC_7_14_6 .LUT_INIT=16'b0101010111111101;
    LogicCell40 \b2v_inst11.dutycycle_RNIEFS24_0_LC_7_14_6  (
            .in0(N__27770),
            .in1(N__25550),
            .in2(N__29678),
            .in3(N__24835),
            .lcout(\b2v_inst11.dutycycle_eena ),
            .ltout(\b2v_inst11.dutycycle_eena_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_0_LC_7_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_0_LC_7_14_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_0_LC_7_14_7 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \b2v_inst11.dutycycle_0_LC_7_14_7  (
            .in0(N__22942),
            .in1(N__22951),
            .in2(N__22945),
            .in3(N__27610),
            .lcout(\b2v_inst11.dutycycleZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34659),
            .ce(),
            .sr(N__24214));
    defparam \b2v_inst11.count_clk_RNI_2_3_LC_7_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_2_3_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_2_3_LC_7_15_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.count_clk_RNI_2_3_LC_7_15_1  (
            .in0(N__29277),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28158),
            .lcout(N_19_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_9_LC_7_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_9_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_9_LC_7_15_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.count_off_RNI_9_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23383),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_RNIZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNITBKN1_1_LC_7_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNITBKN1_1_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNITBKN1_1_LC_7_15_3 .LUT_INIT=16'b1100110111001111;
    LogicCell40 \b2v_inst11.func_state_RNITBKN1_1_LC_7_15_3  (
            .in0(N__28678),
            .in1(N__24493),
            .in2(N__28290),
            .in3(N__28157),
            .lcout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1 ),
            .ltout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIBHHP2_0_LC_7_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIBHHP2_0_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIBHHP2_0_LC_7_15_4 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \b2v_inst11.func_state_RNIBHHP2_0_LC_7_15_4  (
            .in0(N__23284),
            .in1(_gnd_net_),
            .in2(N__23254),
            .in3(N__23108),
            .lcout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_4_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI2N9T2_1_LC_7_15_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI2N9T2_1_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI2N9T2_1_LC_7_15_5 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \b2v_inst11.func_state_RNI2N9T2_1_LC_7_15_5  (
            .in0(N__27771),
            .in1(N__23231),
            .in2(_gnd_net_),
            .in3(N__23062),
            .lcout(\b2v_inst11.func_state_1_m0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_0_LC_7_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_0_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_0_LC_7_15_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_0_LC_7_15_6  (
            .in0(N__27957),
            .in1(N__25551),
            .in2(N__24378),
            .in3(N__25318),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_0 ),
            .ltout(\b2v_inst11.dutycycle_RNI_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIF6NL_2_LC_7_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIF6NL_2_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIF6NL_2_LC_7_15_7 .LUT_INIT=16'b0011001101111111;
    LogicCell40 \b2v_inst11.dutycycle_RNIF6NL_2_LC_7_15_7  (
            .in0(N__23188),
            .in1(N__23143),
            .in2(N__23134),
            .in3(N__28159),
            .lcout(\b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIS50RB_0_LC_7_16_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIS50RB_0_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIS50RB_0_LC_7_16_0 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \b2v_inst11.func_state_RNIS50RB_0_LC_7_16_0  (
            .in0(N__27604),
            .in1(N__24690),
            .in2(N__23440),
            .in3(N__23448),
            .lcout(\b2v_inst11.func_stateZ0Z_0 ),
            .ltout(\b2v_inst11.func_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_2_0_LC_7_16_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_2_0_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_2_0_LC_7_16_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.func_state_RNI_2_0_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23068),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_3013_i ),
            .ltout(\b2v_inst11.N_3013_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIT4D71_9_LC_7_16_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIT4D71_9_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIT4D71_9_LC_7_16_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst11.count_off_RNIT4D71_9_LC_7_16_2  (
            .in0(N__23414),
            .in1(N__28576),
            .in2(N__23065),
            .in3(N__24082),
            .lcout(\b2v_inst11.N_330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI70K8_0_LC_7_16_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI70K8_0_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI70K8_0_LC_7_16_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.func_state_RNI70K8_0_LC_7_16_4  (
            .in0(N__28276),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23466),
            .lcout(\b2v_inst11.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_0_LC_7_16_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_0_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.func_state_0_LC_7_16_5 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \b2v_inst11.func_state_0_LC_7_16_5  (
            .in0(N__23449),
            .in1(N__23439),
            .in2(N__24694),
            .in3(N__27605),
            .lcout(\b2v_inst11.func_stateZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34669),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_0_9_LC_7_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_0_9_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_0_9_LC_7_16_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_RNI_0_9_LC_7_16_6  (
            .in0(N__23415),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29284),
            .lcout(),
            .ltout(\b2v_inst11.N_335_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNINJ641_9_LC_7_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNINJ641_9_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNINJ641_9_LC_7_16_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \b2v_inst11.count_off_RNINJ641_9_LC_7_16_7  (
            .in0(N__24291),
            .in1(N__24716),
            .in2(N__23386),
            .in3(N__23378),
            .lcout(\b2v_inst11.func_state_1_ss0_i_0_o2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI_2_LC_8_1_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI_2_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI_2_LC_8_1_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst36.count_RNI_2_LC_8_1_0  (
            .in0(N__29968),
            .in1(N__24918),
            .in2(N__25179),
            .in3(N__29909),
            .lcout(\b2v_inst36.un12_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_2_c_RNIBSB8_LC_8_1_1 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_2_c_RNIBSB8_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_2_c_RNIBSB8_LC_8_1_1 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_2_c_RNIBSB8_LC_8_1_1  (
            .in0(N__29883),
            .in1(N__32205),
            .in2(N__29914),
            .in3(N__32080),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIH5D01_3_LC_8_1_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIH5D01_3_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIH5D01_3_LC_8_1_2 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \b2v_inst36.count_RNIH5D01_3_LC_8_1_2  (
            .in0(N__31932),
            .in1(N__29872),
            .in2(N__23302),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIPHH01_7_LC_8_1_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIPHH01_7_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIPHH01_7_LC_8_1_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIPHH01_7_LC_8_1_3  (
            .in0(N__23296),
            .in1(N__31934),
            .in2(_gnd_net_),
            .in3(N__23488),
            .lcout(\b2v_inst36.countZ0Z_7 ),
            .ltout(\b2v_inst36.countZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_7_LC_8_1_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_7_LC_8_1_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_7_LC_8_1_4 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst36.count_7_LC_8_1_4  (
            .in0(N__32082),
            .in1(N__32208),
            .in2(N__23299),
            .in3(N__25156),
            .lcout(\b2v_inst36.count_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34682),
            .ce(N__31935),
            .sr(N__31827));
    defparam \b2v_inst36.un2_count_1_cry_4_c_RNID0E8_LC_8_1_5 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_4_c_RNID0E8_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_4_c_RNID0E8_LC_8_1_5 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_4_c_RNID0E8_LC_8_1_5  (
            .in0(N__24903),
            .in1(N__32206),
            .in2(N__24922),
            .in3(N__32081),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNILBF01_5_LC_8_1_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNILBF01_5_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNILBF01_5_LC_8_1_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst36.count_RNILBF01_5_LC_8_1_6  (
            .in0(N__31933),
            .in1(_gnd_net_),
            .in2(N__23500),
            .in3(N__23494),
            .lcout(\b2v_inst36.countZ0Z_5 ),
            .ltout(\b2v_inst36.countZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_5_LC_8_1_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_5_LC_8_1_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_5_LC_8_1_7 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst36.count_5_LC_8_1_7  (
            .in0(N__24904),
            .in1(N__32207),
            .in2(N__23497),
            .in3(N__32083),
            .lcout(\b2v_inst36.count_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34682),
            .ce(N__31935),
            .sr(N__31827));
    defparam \b2v_inst36.un2_count_1_cry_10_c_RNIQ3J1_LC_8_2_0 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_10_c_RNIQ3J1_LC_8_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_10_c_RNIQ3J1_LC_8_2_0 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_10_c_RNIQ3J1_LC_8_2_0  (
            .in0(N__32086),
            .in1(N__30084),
            .in2(N__29749),
            .in3(N__32197),
            .lcout(\b2v_inst36.count_rst_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_6_c_RNIF4G8_LC_8_2_1 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_6_c_RNIF4G8_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_6_c_RNIF4G8_LC_8_2_1 .LUT_INIT=16'b0000010000001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_6_c_RNIF4G8_LC_8_2_1  (
            .in0(N__25180),
            .in1(N__32193),
            .in2(N__32089),
            .in3(N__25152),
            .lcout(\b2v_inst36.count_rst_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_7_c_RNIG6H8_LC_8_2_2 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_7_c_RNIG6H8_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_7_c_RNIG6H8_LC_8_2_2 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_7_c_RNIG6H8_LC_8_2_2  (
            .in0(N__32084),
            .in1(N__29859),
            .in2(N__25138),
            .in3(N__32196),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIRKI01_8_LC_8_2_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIRKI01_8_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIRKI01_8_LC_8_2_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.count_RNIRKI01_8_LC_8_2_3  (
            .in0(_gnd_net_),
            .in1(N__23476),
            .in2(N__23482),
            .in3(N__31907),
            .lcout(\b2v_inst36.countZ0Z_8 ),
            .ltout(\b2v_inst36.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_8_LC_8_2_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_8_LC_8_2_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_8_LC_8_2_4 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \b2v_inst36.count_8_LC_8_2_4  (
            .in0(N__32087),
            .in1(N__25137),
            .in2(N__23479),
            .in3(N__32198),
            .lcout(\b2v_inst36.count_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34675),
            .ce(N__31976),
            .sr(N__31840));
    defparam \b2v_inst36.un2_count_1_cry_9_c_RNIIAJ8_LC_8_2_5 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_9_c_RNIIAJ8_LC_8_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_9_c_RNIIAJ8_LC_8_2_5 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_9_c_RNIIAJ8_LC_8_2_5  (
            .in0(N__25116),
            .in1(N__32194),
            .in2(N__29841),
            .in3(N__32085),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI6MB61_10_LC_8_2_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI6MB61_10_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI6MB61_10_LC_8_2_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst36.count_RNI6MB61_10_LC_8_2_6  (
            .in0(N__31908),
            .in1(_gnd_net_),
            .in2(N__23470),
            .in3(N__23575),
            .lcout(\b2v_inst36.countZ0Z_10 ),
            .ltout(\b2v_inst36.countZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_10_LC_8_2_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_10_LC_8_2_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_10_LC_8_2_7 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst36.count_10_LC_8_2_7  (
            .in0(N__25117),
            .in1(N__32195),
            .in2(N__23578),
            .in3(N__32088),
            .lcout(\b2v_inst36.count_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34675),
            .ce(N__31976),
            .sr(N__31840));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_8_3_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_8_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__27426),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_8_3_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_8_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(N__23684),
            .in2(N__23569),
            .in3(N__23557),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_8_3_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_8_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_8_3_2  (
            .in0(_gnd_net_),
            .in1(N__23554),
            .in2(N__23689),
            .in3(N__23548),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_8_3_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_8_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(N__23714),
            .in2(N__23545),
            .in3(N__23536),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_8_3_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_8_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_8_3_4  (
            .in0(_gnd_net_),
            .in1(N__23533),
            .in2(N__23719),
            .in3(N__23527),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_8_3_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_8_3_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_8_3_5  (
            .in0(N__23613),
            .in1(N__23688),
            .in2(N__23524),
            .in3(N__23512),
            .lcout(\b2v_inst11.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_8_3_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_8_3_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_8_3_6  (
            .in0(N__23509),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23503),
            .lcout(\b2v_inst11.mult1_un152_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_8_3_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_8_3_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_8_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23713),
            .lcout(\b2v_inst11.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_8_4_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_8_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_8_4_0  (
            .in0(_gnd_net_),
            .in1(N__25384),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_8_4_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_8_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_8_4_1  (
            .in0(_gnd_net_),
            .in1(N__23588),
            .in2(N__24343),
            .in3(N__23674),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_1 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_8_4_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_8_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(N__23671),
            .in2(N__23593),
            .in3(N__23665),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_8_4_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_8_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(N__23615),
            .in2(N__23662),
            .in3(N__23653),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_8_4_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_8_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_8_4_4  (
            .in0(_gnd_net_),
            .in1(N__23650),
            .in2(N__23620),
            .in3(N__23644),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_8_4_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_8_4_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_8_4_5  (
            .in0(N__25464),
            .in1(N__23592),
            .in2(N__23641),
            .in3(N__23632),
            .lcout(\b2v_inst11.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_8_4_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_8_4_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_8_4_6  (
            .in0(N__23629),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23623),
            .lcout(\b2v_inst11.mult1_un159_sum_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_8_4_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_8_4_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_8_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23614),
            .lcout(\b2v_inst11.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIQF4M_14_LC_8_5_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIQF4M_14_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIQF4M_14_LC_8_5_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNIQF4M_14_LC_8_5_0  (
            .in0(N__23743),
            .in1(N__34055),
            .in2(_gnd_net_),
            .in3(N__23847),
            .lcout(\b2v_inst11.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_14_LC_8_5_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_14_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_14_LC_8_5_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_14_LC_8_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23851),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34661),
            .ce(N__33687),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIS3FN_6_LC_8_5_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIS3FN_6_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIS3FN_6_LC_8_5_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNIS3FN_6_LC_8_5_2  (
            .in0(N__23737),
            .in1(N__34053),
            .in2(_gnd_net_),
            .in3(N__23775),
            .lcout(\b2v_inst11.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_6_LC_8_5_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_6_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_6_LC_8_5_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_6_LC_8_5_3  (
            .in0(N__23776),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34661),
            .ce(N__33687),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNISI5M_15_LC_8_5_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNISI5M_15_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNISI5M_15_LC_8_5_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNISI5M_15_LC_8_5_4  (
            .in0(N__23731),
            .in1(N__34056),
            .in2(_gnd_net_),
            .in3(N__23826),
            .lcout(\b2v_inst11.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_15_LC_8_5_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_15_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_15_LC_8_5_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_15_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23830),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34661),
            .ce(N__33687),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIU6GN_7_LC_8_5_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIU6GN_7_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIU6GN_7_LC_8_5_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNIU6GN_7_LC_8_5_6  (
            .in0(N__23725),
            .in1(N__34054),
            .in2(_gnd_net_),
            .in3(N__23763),
            .lcout(\b2v_inst11.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_7_LC_8_5_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_7_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_7_LC_8_5_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_7_LC_8_5_7  (
            .in0(N__23764),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34661),
            .ce(N__33687),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_1_c_LC_8_6_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_1_c_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_1_c_LC_8_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_count_cry_1_c_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__26517),
            .in2(N__26559),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\b2v_inst11.un1_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_8_6_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_8_6_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_8_6_1  (
            .in0(N__26479),
            .in1(_gnd_net_),
            .in2(N__25921),
            .in3(N__23788),
            .lcout(\b2v_inst11.un1_count_cry_1_c_RNIIIQDZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_1 ),
            .carryout(\b2v_inst11.un1_count_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_8_6_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_8_6_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_8_6_2  (
            .in0(N__26483),
            .in1(_gnd_net_),
            .in2(N__25620),
            .in3(N__23785),
            .lcout(\b2v_inst11.un1_count_cry_2_c_RNIJKRDZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_2 ),
            .carryout(\b2v_inst11.un1_count_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_8_6_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_8_6_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_8_6_3  (
            .in0(N__26480),
            .in1(_gnd_net_),
            .in2(N__26025),
            .in3(N__23782),
            .lcout(\b2v_inst11.un1_count_cry_3_c_RNIKMSDZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_3 ),
            .carryout(\b2v_inst11.un1_count_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_8_6_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_8_6_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_8_6_4  (
            .in0(N__26484),
            .in1(_gnd_net_),
            .in2(N__25983),
            .in3(N__23779),
            .lcout(\b2v_inst11.un1_count_cry_4_c_RNILOTDZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_4 ),
            .carryout(\b2v_inst11.un1_count_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_8_6_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_8_6_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_8_6_5  (
            .in0(N__26481),
            .in1(_gnd_net_),
            .in2(N__25759),
            .in3(N__23767),
            .lcout(\b2v_inst11.un1_count_cry_5_c_RNIMQUDZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_5 ),
            .carryout(\b2v_inst11.un1_count_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_8_6_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_8_6_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_8_6_6  (
            .in0(N__26485),
            .in1(_gnd_net_),
            .in2(N__25893),
            .in3(N__23755),
            .lcout(\b2v_inst11.un1_count_cry_6_c_RNINSVDZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_6 ),
            .carryout(\b2v_inst11.un1_count_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_8_6_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_8_6_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_8_6_7  (
            .in0(N__26482),
            .in1(N__26396),
            .in2(_gnd_net_),
            .in3(N__23752),
            .lcout(\b2v_inst11.un1_count_cry_7_c_RNIOU0EZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_7 ),
            .carryout(\b2v_inst11.un1_count_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_8_7_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_8_7_0 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_8_7_0  (
            .in0(N__26488),
            .in1(_gnd_net_),
            .in2(N__26354),
            .in3(N__23749),
            .lcout(\b2v_inst11.un1_count_cry_8_c_RNIP02EZ0 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\b2v_inst11.un1_count_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_8_7_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_8_7_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_8_7_1  (
            .in0(N__26462),
            .in1(_gnd_net_),
            .in2(N__25814),
            .in3(N__23746),
            .lcout(\b2v_inst11.un1_count_cry_9_c_RNIQ23EZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_9 ),
            .carryout(\b2v_inst11.un1_count_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_8_7_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_8_7_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_8_7_2  (
            .in0(N__26489),
            .in1(N__25835),
            .in2(_gnd_net_),
            .in3(N__23860),
            .lcout(\b2v_inst11.un1_count_cry_10_c_RNI24RZ0Z6 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_10 ),
            .carryout(\b2v_inst11.un1_count_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_8_7_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_8_7_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_8_7_3  (
            .in0(N__26463),
            .in1(_gnd_net_),
            .in2(N__25788),
            .in3(N__23857),
            .lcout(\b2v_inst11.un1_count_cry_11_c_RNI36SZ0Z6 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_11 ),
            .carryout(\b2v_inst11.un1_count_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_8_7_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_8_7_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_8_7_4  (
            .in0(N__26490),
            .in1(_gnd_net_),
            .in2(N__26070),
            .in3(N__23854),
            .lcout(\b2v_inst11.un1_count_cry_12_c_RNI48TZ0Z6 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_12 ),
            .carryout(\b2v_inst11.un1_count_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_8_7_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_8_7_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_8_7_5  (
            .in0(N__26464),
            .in1(_gnd_net_),
            .in2(N__25735),
            .in3(N__23836),
            .lcout(\b2v_inst11.un1_count_cry_13_c_RNI5AUZ0Z6 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_13 ),
            .carryout(\b2v_inst11.un1_count_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_8_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_8_7_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_8_7_6  (
            .in0(N__26491),
            .in1(N__25870),
            .in2(_gnd_net_),
            .in3(N__23833),
            .lcout(\b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIM92M_12_LC_8_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIM92M_12_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIM92M_12_LC_8_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNIM92M_12_LC_8_7_7  (
            .in0(N__23893),
            .in1(N__34057),
            .in2(_gnd_net_),
            .in3(N__23904),
            .lcout(\b2v_inst11.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIB49T_10_LC_8_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIB49T_10_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIB49T_10_LC_8_8_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_RNIB49T_10_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__23803),
            .in2(N__23815),
            .in3(N__34051),
            .lcout(\b2v_inst11.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_10_LC_8_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_10_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_10_LC_8_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_10_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23814),
            .lcout(\b2v_inst11.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34646),
            .ce(N__33682),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIK61M_11_LC_8_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIK61M_11_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIK61M_11_LC_8_8_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNIK61M_11_LC_8_8_2  (
            .in0(N__23929),
            .in1(N__34052),
            .in2(_gnd_net_),
            .in3(N__23796),
            .lcout(\b2v_inst11.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_11_LC_8_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_11_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_11_LC_8_8_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_11_LC_8_8_3  (
            .in0(N__23797),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34646),
            .ce(N__33682),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIKNAN_2_LC_8_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIKNAN_2_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIKNAN_2_LC_8_8_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNIKNAN_2_LC_8_8_4  (
            .in0(N__23911),
            .in1(N__34050),
            .in2(_gnd_net_),
            .in3(N__23922),
            .lcout(\b2v_inst11.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_2_LC_8_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_2_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_2_LC_8_8_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_2_LC_8_8_5  (
            .in0(N__23923),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34646),
            .ce(N__33682),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_12_LC_8_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_12_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_12_LC_8_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_12_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23905),
            .lcout(\b2v_inst11.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34646),
            .ce(N__33682),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_a2_0_LC_8_9_0 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_a2_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_a2_0_LC_8_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst5.curr_state_7_1_0__m6_i_a2_0_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__23874),
            .in2(_gnd_net_),
            .in3(N__32959),
            .lcout(G_2727),
            .ltout(G_2727_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_1_LC_8_9_1 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_1_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst5.curr_state_1_LC_8_9_1 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \b2v_inst5.curr_state_1_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23887),
            .in3(N__26668),
            .lcout(\b2v_inst5.curr_state_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34629),
            .ce(N__33680),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_LC_8_9_2 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst5.RSMRSTn_LC_8_9_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \b2v_inst5.RSMRSTn_LC_8_9_2  (
            .in0(N__34753),
            .in1(N__26306),
            .in2(_gnd_net_),
            .in3(N__23875),
            .lcout(RSMRSTn_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34629),
            .ce(N__33680),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNITB7B1_1_LC_8_9_3 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNITB7B1_1_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNITB7B1_1_LC_8_9_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \b2v_inst5.curr_state_RNITB7B1_1_LC_8_9_3  (
            .in0(N__23873),
            .in1(N__34065),
            .in2(N__26308),
            .in3(N__34756),
            .lcout(\b2v_inst5.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_o3_0_LC_8_9_4 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_o3_0_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_o3_0_LC_8_9_4 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \b2v_inst5.curr_state_7_1_0__m6_i_o3_0_LC_8_9_4  (
            .in0(N__34754),
            .in1(N__26301),
            .in2(_gnd_net_),
            .in3(N__23872),
            .lcout(N_229),
            .ltout(N_229_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNI76HI_1_LC_8_9_5 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNI76HI_1_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNI76HI_1_LC_8_9_5 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \b2v_inst5.curr_state_RNI76HI_1_LC_8_9_5  (
            .in0(N__26282),
            .in1(N__23884),
            .in2(N__23878),
            .in3(N__34064),
            .lcout(\b2v_inst5.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst5.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNI5VS71_1_LC_8_9_6 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNI5VS71_1_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNI5VS71_1_LC_8_9_6 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \b2v_inst5.curr_state_RNI5VS71_1_LC_8_9_6  (
            .in0(N__34755),
            .in1(_gnd_net_),
            .in2(N__23959),
            .in3(N__26305),
            .lcout(curr_state_RNI5VS71_0_1),
            .ltout(curr_state_RNI5VS71_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_0_LC_8_9_7 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_0_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst5.curr_state_0_LC_8_9_7 .LUT_INIT=16'b1111001011110010;
    LogicCell40 \b2v_inst5.curr_state_0_LC_8_9_7  (
            .in0(N__26283),
            .in1(N__26307),
            .in2(N__23956),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.curr_state_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34629),
            .ce(N__33680),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_3_LC_8_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_3_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_3_LC_8_10_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_3_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__25589),
            .in2(_gnd_net_),
            .in3(N__24795),
            .lcout(\b2v_inst11.mult1_un145_sum ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_fast_LC_8_10_1 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_fast_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.tmp_1_fast_LC_8_10_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst20.tmp_1_fast_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__24455),
            .in2(_gnd_net_),
            .in3(N__26866),
            .lcout(SYNTHESIZED_WIRE_47keep_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34645),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_0_c_RNO_LC_8_10_2 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_0_c_RNO_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_0_c_RNO_LC_8_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_0_c_RNO_LC_8_10_2  (
            .in0(N__31079),
            .in1(N__31001),
            .in2(N__31044),
            .in3(N__31108),
            .lcout(\b2v_inst20.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.G_146_LC_8_10_3 .C_ON=1'b0;
    defparam \b2v_inst36.G_146_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.G_146_LC_8_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst36.G_146_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__26925),
            .in2(_gnd_net_),
            .in3(N__26827),
            .lcout(b2v_inst16_delayed_vddq_pwrgd_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_RNI8DFE_LC_8_10_4 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_RNI8DFE_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.RSMRSTn_RNI8DFE_LC_8_10_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \b2v_inst5.RSMRSTn_RNI8DFE_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__27071),
            .in2(N__24468),
            .in3(N__27004),
            .lcout(RSMRSTn_RNI8DFE),
            .ltout(RSMRSTn_RNI8DFE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o2_LC_8_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o2_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o2_LC_8_10_5 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \b2v_inst11.func_state_0_sqmuxa_0_o2_LC_8_10_5  (
            .in0(N__29328),
            .in1(N__28597),
            .in2(N__23932),
            .in3(N__26924),
            .lcout(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o2_0_LC_8_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o2_0_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o2_0_LC_8_10_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \b2v_inst11.func_state_0_sqmuxa_0_o2_0_LC_8_10_6  (
            .in0(N__26926),
            .in1(N__27070),
            .in2(N__28753),
            .in3(N__28347),
            .lcout(\b2v_inst11.N_182 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIE5T11_2_1_LC_8_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIE5T11_2_1_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIE5T11_2_1_LC_8_11_0 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \b2v_inst11.func_state_RNIE5T11_2_1_LC_8_11_0  (
            .in0(N__28573),
            .in1(N__27091),
            .in2(N__29353),
            .in3(N__29273),
            .lcout(\b2v_inst11.g0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_5_LC_8_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_5_LC_8_11_1 .SEQ_MODE=4'b1011;
    defparam \b2v_inst11.dutycycle_5_LC_8_11_1 .LUT_INIT=16'b1010101011111100;
    LogicCell40 \b2v_inst11.dutycycle_5_LC_8_11_1  (
            .in0(N__24028),
            .in1(N__24018),
            .in2(N__24037),
            .in3(N__27451),
            .lcout(\b2v_inst11.dutycycle_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34649),
            .ce(),
            .sr(N__24164));
    defparam \b2v_inst11.func_state_RNIT4D71_0_1_LC_8_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIT4D71_0_1_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIT4D71_0_1_LC_8_11_2 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \b2v_inst11.func_state_RNIT4D71_0_1_LC_8_11_2  (
            .in0(N__24058),
            .in1(N__28574),
            .in2(_gnd_net_),
            .in3(N__29272),
            .lcout(\b2v_inst11.func_state_RNIT4D71_0Z0Z_1 ),
            .ltout(\b2v_inst11.func_state_RNIT4D71_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIIOE3D_5_LC_8_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIIOE3D_5_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIIOE3D_5_LC_8_11_3 .LUT_INIT=16'b1010101011111100;
    LogicCell40 \b2v_inst11.dutycycle_RNIIOE3D_5_LC_8_11_3  (
            .in0(N__24027),
            .in1(N__24019),
            .in2(N__24004),
            .in3(N__27450),
            .lcout(dutycycle_RNIIOE3D_0_5),
            .ltout(dutycycle_RNIIOE3D_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_5_LC_8_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_5_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_5_LC_8_11_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_5_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24001),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_5 ),
            .ltout(\b2v_inst11.dutycycle_RNI_4Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_LC_8_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_LC_8_11_5 .LUT_INIT=16'b0101010111110101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_LC_8_11_5  (
            .in0(N__25333),
            .in1(_gnd_net_),
            .in2(N__23998),
            .in3(N__28958),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_axb_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_2_LC_8_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_2_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_2_LC_8_11_6 .LUT_INIT=16'b0110100101101001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_2_LC_8_11_6  (
            .in0(N__27986),
            .in1(N__24781),
            .in2(N__23995),
            .in3(N__27409),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_3_LC_8_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_3_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_3_LC_8_11_7 .LUT_INIT=16'b0000000001100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_3_LC_8_11_7  (
            .in0(N__24780),
            .in1(N__27985),
            .in2(N__25360),
            .in3(N__28957),
            .lcout(\b2v_inst11.un1_i3_mux_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_4_LC_8_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_4_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_4_LC_8_12_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_4_LC_8_12_0  (
            .in0(N__28163),
            .in1(N__23971),
            .in2(_gnd_net_),
            .in3(N__28993),
            .lcout(\b2v_inst11.un1_dutycycle_inv_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_LC_8_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_LC_8_12_1 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_LC_8_12_1  (
            .in0(N__24526),
            .in1(N__24421),
            .in2(N__28020),
            .in3(N__28164),
            .lcout(\b2v_inst11.N_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNINJ641_5_LC_8_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNINJ641_5_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNINJ641_5_LC_8_12_2 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \b2v_inst11.dutycycle_RNINJ641_5_LC_8_12_2  (
            .in0(N__28744),
            .in1(N__29092),
            .in2(N__28344),
            .in3(N__24364),
            .lcout(),
            .ltout(\b2v_inst11.g1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIE7D82_2_LC_8_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIE7D82_2_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIE7D82_2_LC_8_12_3 .LUT_INIT=16'b1100110001110010;
    LogicCell40 \b2v_inst11.dutycycle_RNIE7D82_2_LC_8_12_3  (
            .in0(N__24412),
            .in1(N__24406),
            .in2(N__24397),
            .in3(N__24394),
            .lcout(\b2v_inst11.un1_dutycycle_172_m4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.SYNTHESIZED_WIRE_49_i_0_o3_0_LC_8_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.SYNTHESIZED_WIRE_49_i_0_o3_0_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.SYNTHESIZED_WIRE_49_i_0_o3_0_LC_8_12_4 .LUT_INIT=16'b0100111101111111;
    LogicCell40 \b2v_inst11.SYNTHESIZED_WIRE_49_i_0_o3_0_LC_8_12_4  (
            .in0(N__27092),
            .in1(N__26927),
            .in2(N__28752),
            .in3(N__27028),
            .lcout(SYNTHESIZED_WIRE_49_i_0_o3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_5_LC_8_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_5_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_5_LC_8_12_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_5_LC_8_12_5  (
            .in0(N__24365),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28828),
            .lcout(G_26_0_a5_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_12_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_12_6  (
            .in0(N__27408),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINJ641_1_0_LC_8_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINJ641_1_0_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINJ641_1_0_LC_8_12_7 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \b2v_inst11.func_state_RNINJ641_1_0_LC_8_12_7  (
            .in0(N__24324),
            .in1(N__27236),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(b2v_inst11_count_off_1_sqmuxa_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_2_LC_8_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_2_LC_8_13_0 .SEQ_MODE=4'b1011;
    defparam \b2v_inst11.dutycycle_2_LC_8_13_0 .LUT_INIT=16'b0111111100001000;
    LogicCell40 \b2v_inst11.dutycycle_2_LC_8_13_0  (
            .in0(N__27550),
            .in1(N__24586),
            .in2(N__24580),
            .in3(N__24553),
            .lcout(\b2v_inst11.dutycycleZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34660),
            .ce(),
            .sr(N__24236));
    defparam \b2v_inst11.func_state_RNI4IKJB_1_LC_8_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI4IKJB_1_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI4IKJB_1_LC_8_13_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \b2v_inst11.func_state_RNI4IKJB_1_LC_8_13_1  (
            .in0(N__24676),
            .in1(N__27548),
            .in2(N__24628),
            .in3(N__24651),
            .lcout(\b2v_inst11.func_state ),
            .ltout(\b2v_inst11.func_state_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIPKCK_2_LC_8_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIPKCK_2_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIPKCK_2_LC_8_13_2 .LUT_INIT=16'b0000010100010001;
    LogicCell40 \b2v_inst11.dutycycle_RNIPKCK_2_LC_8_13_2  (
            .in0(N__29634),
            .in1(N__29286),
            .in2(N__24592),
            .in3(N__27382),
            .lcout(),
            .ltout(\b2v_inst11.N_303_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNILQFE3_2_LC_8_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNILQFE3_2_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNILQFE3_2_LC_8_13_3 .LUT_INIT=16'b0011011100110011;
    LogicCell40 \b2v_inst11.dutycycle_RNILQFE3_2_LC_8_13_3  (
            .in0(N__24677),
            .in1(N__27754),
            .in2(N__24589),
            .in3(N__24874),
            .lcout(\b2v_inst11.dutycycle_eena_1 ),
            .ltout(\b2v_inst11.dutycycle_eena_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI6O567_2_LC_8_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI6O567_2_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI6O567_2_LC_8_13_4 .LUT_INIT=16'b0111111100100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI6O567_2_LC_8_13_4  (
            .in0(N__27549),
            .in1(N__24579),
            .in2(N__24556),
            .in3(N__24552),
            .lcout(\b2v_inst11.dutycycleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIEFS24_1_LC_8_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIEFS24_1_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIEFS24_1_LC_8_13_7 .LUT_INIT=16'b0000111111101111;
    LogicCell40 \b2v_inst11.dutycycle_RNIEFS24_1_LC_8_13_7  (
            .in0(N__25308),
            .in1(N__29633),
            .in2(N__27741),
            .in3(N__24831),
            .lcout(\b2v_inst11.dutycycle_eena_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIOJI01_1_LC_8_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIOJI01_1_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIOJI01_1_LC_8_14_0 .LUT_INIT=16'b0000010100110101;
    LogicCell40 \b2v_inst11.func_state_RNIOJI01_1_LC_8_14_0  (
            .in0(N__28582),
            .in1(N__28798),
            .in2(N__29671),
            .in3(N__24525),
            .lcout(\b2v_inst11.un1_clk_100khz_26_and_i_o2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIE5T11_1_LC_8_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIE5T11_1_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIE5T11_1_LC_8_14_1 .LUT_INIT=16'b0100111100000000;
    LogicCell40 \b2v_inst11.func_state_RNIE5T11_1_LC_8_14_1  (
            .in0(N__28581),
            .in1(N__28731),
            .in2(N__28346),
            .in3(N__28412),
            .lcout(\b2v_inst11.N_375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_sx_LC_8_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_sx_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_sx_LC_8_14_2 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_sx_LC_8_14_2  (
            .in0(N__28732),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28336),
            .lcout(),
            .ltout(\b2v_inst11.un1_clk_100khz_52_and_i_a2_1_sxZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_LC_8_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_LC_8_14_3 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_LC_8_14_3  (
            .in0(N__27026),
            .in1(N__27108),
            .in2(N__24487),
            .in3(N__24469),
            .lcout(\b2v_inst11.un1_clk_100khz_52_and_i_a2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNINJ641_0_2_LC_8_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNINJ641_0_2_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNINJ641_0_2_LC_8_14_4 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \b2v_inst11.dutycycle_RNINJ641_0_2_LC_8_14_4  (
            .in0(N__27107),
            .in1(N__27027),
            .in2(N__24481),
            .in3(N__24427),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIVFCT3_1_LC_8_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIVFCT3_1_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIVFCT3_1_LC_8_14_5 .LUT_INIT=16'b0100111010101010;
    LogicCell40 \b2v_inst11.func_state_RNIVFCT3_1_LC_8_14_5  (
            .in0(N__24892),
            .in1(N__24886),
            .in2(N__24877),
            .in3(N__29653),
            .lcout(\b2v_inst11.N_183 ),
            .ltout(\b2v_inst11.N_183_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIG8JO1_1_LC_8_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIG8JO1_1_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIG8JO1_1_LC_8_14_6 .LUT_INIT=16'b1111111101001111;
    LogicCell40 \b2v_inst11.func_state_RNIG8JO1_1_LC_8_14_6  (
            .in0(N__29654),
            .in1(N__24867),
            .in2(N__24838),
            .in3(N__24675),
            .lcout(\b2v_inst11.N_114_f0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_3_LC_8_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_3_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_3_LC_8_14_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_3_LC_8_14_7  (
            .in0(N__29268),
            .in1(N__25552),
            .in2(N__25337),
            .in3(N__24820),
            .lcout(\b2v_inst11.g1_4_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_1_ss0_i_0_a2_3_LC_8_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_1_ss0_i_0_a2_3_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_1_ss0_i_0_a2_3_LC_8_15_0 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \b2v_inst11.func_state_1_ss0_i_0_a2_3_LC_8_15_0  (
            .in0(N__28707),
            .in1(N__28252),
            .in2(_gnd_net_),
            .in3(N__29095),
            .lcout(\b2v_inst11.N_379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst31.un8_output_0_LC_8_15_1 .C_ON=1'b0;
    defparam \b2v_inst31.un8_output_0_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst31.un8_output_0_LC_8_15_1 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \b2v_inst31.un8_output_0_LC_8_15_1  (
            .in0(N__29659),
            .in1(N__34743),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst31.un8_outputZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNI8OKQ2_0_LC_8_15_2 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNI8OKQ2_0_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNI8OKQ2_0_LC_8_15_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \b2v_inst6.curr_state_RNI8OKQ2_0_LC_8_15_2  (
            .in0(N__29510),
            .in1(N__27843),
            .in2(_gnd_net_),
            .in3(N__33713),
            .lcout(\b2v_inst6.curr_state_RNI8OKQ2Z0Z_0 ),
            .ltout(\b2v_inst6.curr_state_RNI8OKQ2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNITH2G3_LC_8_15_3 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNITH2G3_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNITH2G3_LC_8_15_3 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_RNITH2G3_LC_8_15_3  (
            .in0(N__24600),
            .in1(N__29511),
            .in2(N__24697),
            .in3(N__29475),
            .lcout(\b2v_inst6.delayed_vccin_vccinaux_okZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_1_LC_8_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_1_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.func_state_1_LC_8_15_4 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \b2v_inst11.func_state_1_LC_8_15_4  (
            .in0(N__24624),
            .in1(N__27624),
            .in2(N__24689),
            .in3(N__24652),
            .lcout(\b2v_inst11.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34670),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_LC_8_15_5 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_LC_8_15_5 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_LC_8_15_5  (
            .in0(N__24610),
            .in1(N__29513),
            .in2(N__24604),
            .in3(N__29476),
            .lcout(\b2v_inst6.delayed_vccin_vccinaux_ok_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34670),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_LC_8_15_6 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_LC_8_15_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.tmp_1_LC_8_15_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst20.tmp_1_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__33929),
            .in2(_gnd_net_),
            .in3(N__26877),
            .lcout(SYNTHESIZED_WIRE_47keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34670),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNI7OBF3_0_LC_8_15_7 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNI7OBF3_0_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNI7OBF3_0_LC_8_15_7 .LUT_INIT=16'b1010101000100000;
    LogicCell40 \b2v_inst6.curr_state_RNI7OBF3_0_LC_8_15_7  (
            .in0(N__33712),
            .in1(N__29512),
            .in2(N__27844),
            .in3(N__35178),
            .lcout(\b2v_inst6.count_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un1_vddq_en_LC_8_16_4 .C_ON=1'b0;
    defparam \b2v_inst16.un1_vddq_en_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un1_vddq_en_LC_8_16_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst16.un1_vddq_en_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(N__25055),
            .in2(_gnd_net_),
            .in3(N__25006),
            .lcout(VDDQ_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst31.un8_output_LC_8_16_5 .C_ON=1'b0;
    defparam \b2v_inst31.un8_output_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst31.un8_output_LC_8_16_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst31.un8_output_LC_8_16_5  (
            .in0(N__24982),
            .in1(N__24976),
            .in2(N__24970),
            .in3(N__24961),
            .lcout(VCCIN_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_1_c_LC_9_1_0 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_1_c_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_1_c_LC_9_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_1_c_LC_9_1_0  (
            .in0(_gnd_net_),
            .in1(N__32245),
            .in2(N__29818),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_1_0_),
            .carryout(\b2v_inst36.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_9_1_1 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_9_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_9_1_1  (
            .in0(_gnd_net_),
            .in1(N__29967),
            .in2(_gnd_net_),
            .in3(N__24931),
            .lcout(\b2v_inst36.un2_count_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_1 ),
            .carryout(\b2v_inst36.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_9_1_2 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_9_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_9_1_2  (
            .in0(_gnd_net_),
            .in1(N__29905),
            .in2(_gnd_net_),
            .in3(N__24928),
            .lcout(\b2v_inst36.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_2 ),
            .carryout(\b2v_inst36.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_3_c_RNICUC8_LC_9_1_3 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_3_c_RNICUC8_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_3_c_RNICUC8_LC_9_1_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_3_c_RNICUC8_LC_9_1_3  (
            .in0(N__32214),
            .in1(N__30442),
            .in2(_gnd_net_),
            .in3(N__24925),
            .lcout(\b2v_inst36.count_rst_10 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_3 ),
            .carryout(\b2v_inst36.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_9_1_4 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_9_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_9_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_9_1_4  (
            .in0(_gnd_net_),
            .in1(N__24917),
            .in2(_gnd_net_),
            .in3(N__24895),
            .lcout(\b2v_inst36.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_4 ),
            .carryout(\b2v_inst36.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_5_c_RNINEG01_LC_9_1_5 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_5_c_RNINEG01_LC_9_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_5_c_RNINEG01_LC_9_1_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_5_c_RNINEG01_LC_9_1_5  (
            .in0(N__32215),
            .in1(N__29770),
            .in2(_gnd_net_),
            .in3(N__25183),
            .lcout(\b2v_inst36.count_rst_8 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_5 ),
            .carryout(\b2v_inst36.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_9_1_6 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_9_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_9_1_6  (
            .in0(_gnd_net_),
            .in1(N__25172),
            .in2(_gnd_net_),
            .in3(N__25141),
            .lcout(\b2v_inst36.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_6 ),
            .carryout(\b2v_inst36.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_9_1_7 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_9_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_9_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_9_1_7  (
            .in0(_gnd_net_),
            .in1(N__29858),
            .in2(_gnd_net_),
            .in3(N__25123),
            .lcout(\b2v_inst36.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_7 ),
            .carryout(\b2v_inst36.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_8_c_RNIH8I8_LC_9_2_0 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_8_c_RNIH8I8_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_8_c_RNIH8I8_LC_9_2_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst36.un2_count_1_cry_8_c_RNIH8I8_LC_9_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31552),
            .in3(N__25120),
            .lcout(\b2v_inst36.un2_count_1_cry_8_c_RNIH8IZ0Z8 ),
            .ltout(),
            .carryin(bfn_9_2_0_),
            .carryout(\b2v_inst36.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_9_2_1 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_9_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_9_2_1  (
            .in0(_gnd_net_),
            .in1(N__29834),
            .in2(_gnd_net_),
            .in3(N__25108),
            .lcout(\b2v_inst36.un2_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_9 ),
            .carryout(\b2v_inst36.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_9_2_2 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_9_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_9_2_2  (
            .in0(_gnd_net_),
            .in1(N__29745),
            .in2(_gnd_net_),
            .in3(N__25105),
            .lcout(\b2v_inst36.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_10 ),
            .carryout(\b2v_inst36.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_11_c_RNIR5K1_LC_9_2_3 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_11_c_RNIR5K1_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_11_c_RNIR5K1_LC_9_2_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_11_c_RNIR5K1_LC_9_2_3  (
            .in0(N__32199),
            .in1(N__30027),
            .in2(_gnd_net_),
            .in3(N__25102),
            .lcout(\b2v_inst36.count_rst_2 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_11 ),
            .carryout(\b2v_inst36.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_12_c_RNIS7L1_LC_9_2_4 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_12_c_RNIS7L1_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_12_c_RNIS7L1_LC_9_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst36.un2_count_1_cry_12_c_RNIS7L1_LC_9_2_4  (
            .in0(_gnd_net_),
            .in1(N__31569),
            .in2(_gnd_net_),
            .in3(N__25099),
            .lcout(\b2v_inst36.un2_count_1_cry_12_c_RNIS7LZ0Z1 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_12 ),
            .carryout(\b2v_inst36.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_13_c_RNIT9M1_LC_9_2_5 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_13_c_RNIT9M1_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_13_c_RNIT9M1_LC_9_2_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_13_c_RNIT9M1_LC_9_2_5  (
            .in0(N__32200),
            .in1(N__29430),
            .in2(_gnd_net_),
            .in3(N__25246),
            .lcout(\b2v_inst36.count_rst_0 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_13 ),
            .carryout(\b2v_inst36.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_14_c_RNIUBN1_LC_9_2_6 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_14_c_RNIUBN1_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_14_c_RNIUBN1_LC_9_2_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_14_c_RNIUBN1_LC_9_2_6  (
            .in0(N__29415),
            .in1(N__32201),
            .in2(_gnd_net_),
            .in3(N__25243),
            .lcout(\b2v_inst36.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNILPEV_14_LC_9_2_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNILPEV_14_LC_9_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNILPEV_14_LC_9_2_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNILPEV_14_LC_9_2_7  (
            .in0(N__25210),
            .in1(N__31915),
            .in2(_gnd_net_),
            .in3(N__25221),
            .lcout(\b2v_inst36.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_12_LC_9_3_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_12_LC_9_3_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_12_LC_9_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_12_LC_9_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25231),
            .lcout(\b2v_inst36.count_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34677),
            .ce(N__31958),
            .sr(N__31835));
    defparam \b2v_inst36.curr_state_RNIKEBL_1_LC_9_3_1 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNIKEBL_1_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNIKEBL_1_LC_9_3_1 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \b2v_inst36.curr_state_RNIKEBL_1_LC_9_3_1  (
            .in0(N__31800),
            .in1(N__30259),
            .in2(N__30357),
            .in3(N__33716),
            .lcout(\b2v_inst36.count_en ),
            .ltout(\b2v_inst36.count_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIHJCV_12_LC_9_3_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIHJCV_12_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIHJCV_12_LC_9_3_2 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \b2v_inst36.count_RNIHJCV_12_LC_9_3_2  (
            .in0(_gnd_net_),
            .in1(N__25240),
            .in2(N__25234),
            .in3(N__25230),
            .lcout(\b2v_inst36.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_14_LC_9_3_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_14_LC_9_3_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_14_LC_9_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_14_LC_9_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25222),
            .lcout(\b2v_inst36.count_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34677),
            .ce(N__31958),
            .sr(N__31835));
    defparam \b2v_inst36.count_15_LC_9_3_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_15_LC_9_3_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_15_LC_9_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_15_LC_9_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25197),
            .lcout(\b2v_inst36.count_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34677),
            .ce(N__31958),
            .sr(N__31835));
    defparam \b2v_inst36.count_RNINSFV_15_LC_9_3_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNINSFV_15_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNINSFV_15_LC_9_3_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst36.count_RNINSFV_15_LC_9_3_6  (
            .in0(N__31959),
            .in1(_gnd_net_),
            .in2(N__25201),
            .in3(N__25189),
            .lcout(\b2v_inst36.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_4_LC_9_3_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_4_LC_9_3_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_4_LC_9_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_4_LC_9_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30462),
            .lcout(\b2v_inst36.count_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34677),
            .ce(N__31958),
            .sr(N__31835));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_9_4_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_9_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(N__25590),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_4_0_),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_9_4_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_9_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_9_4_1  (
            .in0(_gnd_net_),
            .in1(N__25439),
            .in2(N__25255),
            .in3(N__25466),
            .lcout(G_2890),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_0 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_9_4_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_9_4_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_9_4_2  (
            .in0(_gnd_net_),
            .in1(N__25492),
            .in2(N__25444),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_1 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_9_4_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_9_4_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_9_4_3  (
            .in0(_gnd_net_),
            .in1(N__25467),
            .in2(N__25486),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_9_4_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_9_4_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_9_4_4  (
            .in0(_gnd_net_),
            .in1(N__25477),
            .in2(N__25471),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_9_4_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_9_4_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_9_4_5  (
            .in0(_gnd_net_),
            .in1(N__25443),
            .in2(N__25429),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_9_4_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_9_4_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_9_4_6  (
            .in0(N__25417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25411),
            .lcout(\b2v_inst11.un85_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_9_4_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_9_4_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_9_4_7  (
            .in0(N__25396),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.pwm_out_RNO_0_LC_9_5_0 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_RNO_0_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.pwm_out_RNO_0_LC_9_5_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \b2v_inst11.pwm_out_RNO_0_LC_9_5_0  (
            .in0(N__25663),
            .in1(N__34092),
            .in2(_gnd_net_),
            .in3(N__25679),
            .lcout(\b2v_inst11.pwm_out_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_2_LC_9_5_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_2_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_2_LC_9_5_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst11.count_RNI_2_LC_9_5_1  (
            .in0(N__25919),
            .in1(N__25616),
            .in2(_gnd_net_),
            .in3(N__26021),
            .lcout(\b2v_inst11.un79_clk_100khzlt6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_15_LC_9_5_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_15_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_15_LC_9_5_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst11.count_RNI_15_LC_9_5_2  (
            .in0(N__25889),
            .in1(N__26403),
            .in2(_gnd_net_),
            .in3(N__25862),
            .lcout(\b2v_inst11.un79_clk_100khzlto15_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_9_LC_9_5_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_9_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_9_LC_9_5_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.count_RNI_9_LC_9_5_3  (
            .in0(N__25842),
            .in1(N__25815),
            .in2(N__26365),
            .in3(N__25789),
            .lcout(),
            .ltout(\b2v_inst11.un79_clk_100khzlto15_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_5_LC_9_5_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_5_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_5_LC_9_5_4 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \b2v_inst11.count_RNI_5_LC_9_5_4  (
            .in0(N__25765),
            .in1(N__25757),
            .in2(N__25738),
            .in3(N__25979),
            .lcout(),
            .ltout(\b2v_inst11.un79_clk_100khzlto15_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_13_LC_9_5_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_13_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_13_LC_9_5_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst11.count_RNI_13_LC_9_5_5  (
            .in0(N__25730),
            .in1(N__26066),
            .in2(N__25711),
            .in3(N__25708),
            .lcout(\b2v_inst11.count_RNIZ0Z_13 ),
            .ltout(\b2v_inst11.count_RNIZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.pwm_out_RNO_1_LC_9_5_6 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_RNO_1_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.pwm_out_RNO_1_LC_9_5_6 .LUT_INIT=16'b0101000100010001;
    LogicCell40 \b2v_inst11.pwm_out_RNO_1_LC_9_5_6  (
            .in0(N__25662),
            .in1(N__26610),
            .in2(N__25627),
            .in3(N__34093),
            .lcout(\b2v_inst11.g0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIMQBN_3_LC_9_6_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIMQBN_3_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIMQBN_3_LC_9_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIMQBN_3_LC_9_6_0  (
            .in0(N__34076),
            .in1(N__26077),
            .in2(_gnd_net_),
            .in3(N__26085),
            .lcout(\b2v_inst11.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_3_LC_9_6_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_3_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_3_LC_9_6_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_3_LC_9_6_1  (
            .in0(N__26086),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34662),
            .ce(N__33688),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIOC3M_13_LC_9_6_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIOC3M_13_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIOC3M_13_LC_9_6_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIOC3M_13_LC_9_6_2  (
            .in0(N__34079),
            .in1(N__26035),
            .in2(_gnd_net_),
            .in3(N__26043),
            .lcout(\b2v_inst11.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_13_LC_9_6_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_13_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_13_LC_9_6_3 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_13_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26047),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34662),
            .ce(N__33688),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIOTCN_4_LC_9_6_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIOTCN_4_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIOTCN_4_LC_9_6_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIOTCN_4_LC_9_6_4  (
            .in0(N__34077),
            .in1(N__25993),
            .in2(_gnd_net_),
            .in3(N__26001),
            .lcout(\b2v_inst11.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_4_LC_9_6_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_4_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_4_LC_9_6_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_4_LC_9_6_5  (
            .in0(N__26002),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34662),
            .ce(N__33688),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIQ0EN_5_LC_9_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIQ0EN_5_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIQ0EN_5_LC_9_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIQ0EN_5_LC_9_6_6  (
            .in0(N__34078),
            .in1(N__25951),
            .in2(_gnd_net_),
            .in3(N__25959),
            .lcout(\b2v_inst11.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_5_LC_9_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_5_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_5_LC_9_6_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_5_LC_9_6_7  (
            .in0(N__25960),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34662),
            .ce(N__33688),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI03G9_0_LC_9_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI03G9_0_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI03G9_0_LC_9_7_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNI03G9_0_LC_9_7_0  (
            .in0(N__25945),
            .in1(N__34086),
            .in2(_gnd_net_),
            .in3(N__25933),
            .lcout(\b2v_inst11.countZ0Z_0 ),
            .ltout(\b2v_inst11.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_1_LC_9_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_1_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_1_LC_9_7_1 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \b2v_inst11.count_RNI_1_LC_9_7_1  (
            .in0(N__26555),
            .in1(_gnd_net_),
            .in2(N__25924),
            .in3(N__26486),
            .lcout(),
            .ltout(\b2v_inst11.count_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI14G9_1_LC_9_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI14G9_1_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI14G9_1_LC_9_7_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_RNI14G9_1_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__26413),
            .in2(N__26566),
            .in3(N__34087),
            .lcout(\b2v_inst11.countZ0Z_1 ),
            .ltout(\b2v_inst11.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_1_LC_9_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_1_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_1_LC_9_7_3 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \b2v_inst11.count_1_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(N__26518),
            .in2(N__26494),
            .in3(N__26487),
            .lcout(\b2v_inst11.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34655),
            .ce(N__33685),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI0AHN_8_LC_9_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI0AHN_8_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI0AHN_8_LC_9_7_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNI0AHN_8_LC_9_7_4  (
            .in0(N__26371),
            .in1(N__34088),
            .in2(_gnd_net_),
            .in3(N__26379),
            .lcout(\b2v_inst11.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_8_LC_9_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_8_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_8_LC_9_7_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_8_LC_9_7_5  (
            .in0(N__26380),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34655),
            .ce(N__33685),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI2DIN_9_LC_9_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI2DIN_9_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI2DIN_9_LC_9_7_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNI2DIN_9_LC_9_7_6  (
            .in0(N__26320),
            .in1(N__34089),
            .in2(_gnd_net_),
            .in3(N__26328),
            .lcout(\b2v_inst11.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_9_LC_9_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_9_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_9_LC_9_7_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_9_LC_9_7_7  (
            .in0(N__26329),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34655),
            .ce(N__33685),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNI65HI_0_LC_9_8_0 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNI65HI_0_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNI65HI_0_LC_9_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst5.curr_state_RNI65HI_0_LC_9_8_0  (
            .in0(N__26266),
            .in1(N__26314),
            .in2(_gnd_net_),
            .in3(N__34090),
            .lcout(\b2v_inst5.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst5.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_LC_9_8_1 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_LC_9_8_1 .LUT_INIT=16'b1111111100001010;
    LogicCell40 \b2v_inst5.curr_state_7_1_0__m4_0_LC_9_8_1  (
            .in0(N__26284),
            .in1(_gnd_net_),
            .in2(N__26269),
            .in3(N__27089),
            .lcout(\b2v_inst5.m4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNITBKN1_7_LC_9_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNITBKN1_7_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNITBKN1_7_LC_9_8_2 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNITBKN1_7_LC_9_8_2  (
            .in0(N__27088),
            .in1(N__26260),
            .in2(_gnd_net_),
            .in3(N__26233),
            .lcout(\b2v_inst11.dutycycle_RNITBKN1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_en_LC_9_8_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_en_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_en_LC_9_8_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst5.count_en_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__26667),
            .in2(_gnd_net_),
            .in3(N__27593),
            .lcout(\b2v_inst5.count_enZ0 ),
            .ltout(\b2v_inst5.count_enZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNICVEB2_6_LC_9_8_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNICVEB2_6_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNICVEB2_6_LC_9_8_4 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \b2v_inst5.count_RNICVEB2_6_LC_9_8_4  (
            .in0(N__30676),
            .in1(N__30745),
            .in2(N__26656),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.un2_count_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.pwm_out_LC_9_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_LC_9_8_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.pwm_out_LC_9_8_5 .LUT_INIT=16'b0010001011101010;
    LogicCell40 \b2v_inst11.pwm_out_LC_9_8_5  (
            .in0(N__26606),
            .in1(N__27594),
            .in2(N__26653),
            .in3(N__26620),
            .lcout(\b2v_inst11.pwm_outZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34651),
            .ce(),
            .sr(N__26587));
    defparam \b2v_inst5.count_RNIE2GB2_7_LC_9_8_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIE2GB2_7_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIE2GB2_7_LC_9_8_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNIE2GB2_7_LC_9_8_6  (
            .in0(N__30214),
            .in1(N__32546),
            .in2(_gnd_net_),
            .in3(N__30868),
            .lcout(\b2v_inst5.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIA2IH2_14_LC_9_8_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIA2IH2_14_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIA2IH2_14_LC_9_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst5.count_RNIA2IH2_14_LC_9_8_7  (
            .in0(N__32547),
            .in1(N__30229),
            .in2(_gnd_net_),
            .in3(N__30774),
            .lcout(\b2v_inst5.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_0_c_LC_9_9_0 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_0_c_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_0_c_LC_9_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_0_c_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26575),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\b2v_inst20.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_1_c_LC_9_9_1 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_1_c_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_1_c_LC_9_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_1_c_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26689),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_0 ),
            .carryout(\b2v_inst20.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_2_c_LC_9_9_2 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_2_c_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_2_c_LC_9_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_2_c_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33370),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_1 ),
            .carryout(\b2v_inst20.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_3_c_LC_9_9_3 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_3_c_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_3_c_LC_9_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_3_c_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__33304),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_2 ),
            .carryout(\b2v_inst20.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_4_c_LC_9_9_4 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_4_c_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_4_c_LC_9_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_4_c_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33241),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_3 ),
            .carryout(\b2v_inst20.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_5_c_LC_9_9_5 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_5_c_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_5_c_LC_9_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_5_c_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33175),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_4 ),
            .carryout(\b2v_inst20.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_6_c_LC_9_9_6 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_6_c_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_6_c_LC_9_9_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_6_c_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33100),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_5 ),
            .carryout(\b2v_inst20.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_7_c_LC_9_9_7 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_7_c_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_7_c_LC_9_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_7_c_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__33433),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_6 ),
            .carryout(b2v_inst20_un4_counter_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_9_10_0.C_ON=1'b0;
    defparam b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_9_10_0.SEQ_MODE=4'b0000;
    defparam b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_9_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_9_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26692),
            .lcout(b2v_inst20_un4_counter_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_6_LC_9_10_1 .C_ON=1'b0;
    defparam \b2v_inst20.counter_6_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_6_LC_9_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst20.counter_6_LC_9_10_1  (
            .in0(N__26848),
            .in1(N__30929),
            .in2(_gnd_net_),
            .in3(N__30913),
            .lcout(\b2v_inst20.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34650),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_2_LC_9_10_2 .C_ON=1'b0;
    defparam \b2v_inst20.counter_2_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_2_LC_9_10_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \b2v_inst20.counter_2_LC_9_10_2  (
            .in0(N__31063),
            .in1(N__31083),
            .in2(_gnd_net_),
            .in3(N__26849),
            .lcout(\b2v_inst20.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34650),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_5_LC_9_10_3 .C_ON=1'b0;
    defparam \b2v_inst20.counter_5_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_5_LC_9_10_3 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \b2v_inst20.counter_5_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__30966),
            .in2(N__26867),
            .in3(N__30952),
            .lcout(\b2v_inst20.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34650),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_1_c_RNO_LC_9_10_4 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_1_c_RNO_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_1_c_RNO_LC_9_10_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst20.un4_counter_1_c_RNO_LC_9_10_4  (
            .in0(N__30965),
            .in1(N__31136),
            .in2(N__30933),
            .in3(N__31231),
            .lcout(\b2v_inst20.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.SYNTHESIZED_WIRE_48_i_0_o3_2_LC_9_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.SYNTHESIZED_WIRE_48_i_0_o3_2_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.SYNTHESIZED_WIRE_48_i_0_o3_2_LC_9_10_5 .LUT_INIT=16'b0111011101011111;
    LogicCell40 \b2v_inst11.SYNTHESIZED_WIRE_48_i_0_o3_2_LC_9_10_5  (
            .in0(N__28348),
            .in1(N__27087),
            .in2(N__27025),
            .in3(N__26923),
            .lcout(SYNTHESIZED_WIRE_48_i_0_o3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_LC_9_10_6 .C_ON=1'b0;
    defparam \b2v_inst20.counter_1_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_1_LC_9_10_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \b2v_inst20.counter_1_LC_9_10_6  (
            .in0(N__31140),
            .in1(N__26844),
            .in2(_gnd_net_),
            .in3(N__31112),
            .lcout(\b2v_inst20.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34650),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_3_LC_9_10_7 .C_ON=1'b0;
    defparam \b2v_inst20.counter_3_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_3_LC_9_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst20.counter_3_LC_9_10_7  (
            .in0(N__26843),
            .in1(N__31021),
            .in2(_gnd_net_),
            .in3(N__31043),
            .lcout(\b2v_inst20.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34650),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_5_LC_9_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_5_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_5_LC_9_11_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_5_LC_9_11_0  (
            .in0(N__28434),
            .in1(N__26742),
            .in2(_gnd_net_),
            .in3(N__29285),
            .lcout(),
            .ltout(\b2v_inst11.N_234_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIG8JO1_5_LC_9_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIG8JO1_5_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIG8JO1_5_LC_9_11_1 .LUT_INIT=16'b1000100010001111;
    LogicCell40 \b2v_inst11.dutycycle_RNIG8JO1_5_LC_9_11_1  (
            .in0(N__29072),
            .in1(N__27442),
            .in2(N__26971),
            .in3(N__29639),
            .lcout(),
            .ltout(\b2v_inst11.un1_clk_100khz_52_and_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI8S5P2_5_LC_9_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI8S5P2_5_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI8S5P2_5_LC_9_11_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \b2v_inst11.dutycycle_RNI8S5P2_5_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__29615),
            .in2(N__26968),
            .in3(N__28575),
            .lcout(\b2v_inst11.g2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_rep1_LC_9_11_5 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_rep1_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.tmp_1_rep1_LC_9_11_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst20.tmp_1_rep1_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__26851),
            .in2(_gnd_net_),
            .in3(N__26942),
            .lcout(SYNTHESIZED_WIRE_47keep_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34654),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_0_LC_9_11_7 .C_ON=1'b0;
    defparam \b2v_inst20.counter_0_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_0_LC_9_11_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \b2v_inst20.counter_0_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__26850),
            .in2(_gnd_net_),
            .in3(N__31113),
            .lcout(\b2v_inst20.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34654),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_S4n_ibuf_RNINJ641_LC_9_12_0.C_ON=1'b0;
    defparam SLP_S4n_ibuf_RNINJ641_LC_9_12_0.SEQ_MODE=4'b0000;
    defparam SLP_S4n_ibuf_RNINJ641_LC_9_12_0.LUT_INIT=16'b1000100011111000;
    LogicCell40 SLP_S4n_ibuf_RNINJ641_LC_9_12_0 (
            .in0(N__27118),
            .in1(N__29093),
            .in2(N__26764),
            .in3(N__28830),
            .lcout(G_26_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_9_4_LC_9_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_9_4_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_9_4_LC_9_12_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_9_4_LC_9_12_1  (
            .in0(N__28831),
            .in1(N__28762),
            .in2(_gnd_net_),
            .in3(N__27331),
            .lcout(),
            .ltout(G_26_0_a5_2_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_S4n_ibuf_RNIE7D82_LC_9_12_2.C_ON=1'b0;
    defparam SLP_S4n_ibuf_RNIE7D82_LC_9_12_2.SEQ_MODE=4'b0000;
    defparam SLP_S4n_ibuf_RNIE7D82_LC_9_12_2.LUT_INIT=16'b1111111111100100;
    LogicCell40 SLP_S4n_ibuf_RNIE7D82_LC_9_12_2 (
            .in0(N__27832),
            .in1(N__27826),
            .in2(N__27820),
            .in3(N__27817),
            .lcout(),
            .ltout(b2v_inst11_un1_dutycycle_172_m3_0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIL3755_0_LC_9_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIL3755_0_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIL3755_0_LC_9_12_3 .LUT_INIT=16'b0001101111111111;
    LogicCell40 \b2v_inst11.dutycycle_RNIL3755_0_LC_9_12_3  (
            .in0(N__27811),
            .in1(N__27799),
            .in2(N__27793),
            .in3(N__29619),
            .lcout(),
            .ltout(\b2v_inst11.g4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIM0L9A_0_LC_9_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIM0L9A_0_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIM0L9A_0_LC_9_12_4 .LUT_INIT=16'b0100000011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNIM0L9A_0_LC_9_12_4  (
            .in0(N__27790),
            .in1(N__27695),
            .in2(N__27628),
            .in3(N__27545),
            .lcout(\b2v_inst11.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_x_LC_9_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_x_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_x_LC_9_12_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.un1_clk_100khz_52_and_i_a2_1_x_LC_9_12_5  (
            .in0(N__28745),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28332),
            .lcout(\b2v_inst11.un1_clk_100khz_52_and_i_a2_1_xZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_2_LC_9_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_2_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_2_LC_9_12_7 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_2_LC_9_12_7  (
            .in0(N__27390),
            .in1(N__28761),
            .in2(_gnd_net_),
            .in3(N__27330),
            .lcout(N_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNINJ641_6_LC_9_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNINJ641_6_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNINJ641_6_LC_9_13_0 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \b2v_inst11.dutycycle_RNINJ641_6_LC_9_13_0  (
            .in0(N__28031),
            .in1(N__27311),
            .in2(_gnd_net_),
            .in3(N__28165),
            .lcout(\b2v_inst11.g3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_S4n_ibuf_RNIF6NL_LC_9_13_1.C_ON=1'b0;
    defparam SLP_S4n_ibuf_RNIF6NL_LC_9_13_1.SEQ_MODE=4'b0000;
    defparam SLP_S4n_ibuf_RNIF6NL_LC_9_13_1.LUT_INIT=16'b0000010000000000;
    LogicCell40 SLP_S4n_ibuf_RNIF6NL_LC_9_13_1 (
            .in0(N__28309),
            .in1(N__28705),
            .in2(N__28837),
            .in3(N__27124),
            .lcout(G_26_0_a5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIE5T11_6_LC_9_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIE5T11_6_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIE5T11_6_LC_9_13_2 .LUT_INIT=16'b0101010101000101;
    LogicCell40 \b2v_inst11.dutycycle_RNIE5T11_6_LC_9_13_2  (
            .in0(N__28029),
            .in1(N__29354),
            .in2(N__29293),
            .in3(N__28592),
            .lcout(),
            .ltout(\b2v_inst11.g2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI2C4V3_6_LC_9_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI2C4V3_6_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI2C4V3_6_LC_9_13_3 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI2C4V3_6_LC_9_13_3  (
            .in0(N__29128),
            .in1(N__27862),
            .in2(N__29122),
            .in3(N__29094),
            .lcout(\b2v_inst11.N_228_N_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIM6F44_LC_9_13_4 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIM6F44_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIM6F44_LC_9_13_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_RNIM6F44_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__29011),
            .in2(_gnd_net_),
            .in3(N__29638),
            .lcout(N_219),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_4_LC_9_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_4_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_4_LC_9_13_5 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_4_LC_9_13_5  (
            .in0(N__28166),
            .in1(N__29002),
            .in2(N__28995),
            .in3(N__28836),
            .lcout(\b2v_inst11.g0_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIE5T11_0_1_LC_9_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIE5T11_0_1_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIE5T11_0_1_LC_9_13_6 .LUT_INIT=16'b0010000000001010;
    LogicCell40 \b2v_inst11.func_state_RNIE5T11_0_1_LC_9_13_6  (
            .in0(N__28706),
            .in1(N__28593),
            .in2(N__28433),
            .in3(N__28311),
            .lcout(),
            .ltout(\b2v_inst11.g1_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIL5HA1_6_LC_9_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIL5HA1_6_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIL5HA1_6_LC_9_13_7 .LUT_INIT=16'b1011010111111111;
    LogicCell40 \b2v_inst11.dutycycle_RNIL5HA1_6_LC_9_13_7  (
            .in0(N__28310),
            .in1(N__28167),
            .in2(N__28039),
            .in3(N__28030),
            .lcout(\b2v_inst11.g1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIRLUM4_11_LC_9_14_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIRLUM4_11_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIRLUM4_11_LC_9_14_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst6.count_RNIRLUM4_11_LC_9_14_0  (
            .in0(N__34346),
            .in1(N__27850),
            .in2(_gnd_net_),
            .in3(N__29395),
            .lcout(\b2v_inst6.countZ0Z_11 ),
            .ltout(\b2v_inst6.countZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_11_LC_9_14_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_11_LC_9_14_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_11_LC_9_14_1 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst6.count_11_LC_9_14_1  (
            .in0(N__35203),
            .in1(N__34939),
            .in2(N__27853),
            .in3(N__31297),
            .lcout(\b2v_inst6.count_3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34671),
            .ce(N__34429),
            .sr(N__35270));
    defparam \b2v_inst6.curr_state_RNIDMSJ1_1_LC_9_14_2 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIDMSJ1_1_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIDMSJ1_1_LC_9_14_2 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \b2v_inst6.curr_state_RNIDMSJ1_1_LC_9_14_2  (
            .in0(N__29706),
            .in1(N__29536),
            .in2(N__29670),
            .in3(N__29722),
            .lcout(\b2v_inst6.curr_state_RNIDMSJ1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_10_c_RNI6P001_LC_9_14_3 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_10_c_RNI6P001_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_10_c_RNI6P001_LC_9_14_3 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_10_c_RNI6P001_LC_9_14_3  (
            .in0(N__35202),
            .in1(N__34937),
            .in2(N__31488),
            .in3(N__31296),
            .lcout(\b2v_inst6.count_rst_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_3_c_RNIO6IO_LC_9_14_4 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_3_c_RNIO6IO_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_3_c_RNIO6IO_LC_9_14_4 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_3_c_RNIO6IO_LC_9_14_4  (
            .in0(N__34936),
            .in1(N__31332),
            .in2(N__35054),
            .in3(N__35201),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIVJVD4_4_LC_9_14_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIVJVD4_4_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIVJVD4_4_LC_9_14_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNIVJVD4_4_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__29383),
            .in2(N__29389),
            .in3(N__34345),
            .lcout(\b2v_inst6.countZ0Z_4 ),
            .ltout(\b2v_inst6.countZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_4_LC_9_14_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_4_LC_9_14_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_4_LC_9_14_6 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \b2v_inst6.count_4_LC_9_14_6  (
            .in0(N__34938),
            .in1(N__31333),
            .in2(N__29386),
            .in3(N__35205),
            .lcout(\b2v_inst6.count_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34671),
            .ce(N__34429),
            .sr(N__35270));
    defparam \b2v_inst6.count_5_LC_9_14_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_5_LC_9_14_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_5_LC_9_14_7 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst6.count_5_LC_9_14_7  (
            .in0(N__35204),
            .in1(N__34940),
            .in2(N__31378),
            .in3(N__35131),
            .lcout(\b2v_inst6.count_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34671),
            .ce(N__34429),
            .sr(N__35270));
    defparam \b2v_inst6.curr_state_RNIVVMK_0_LC_9_15_0 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIVVMK_0_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIVVMK_0_LC_9_15_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst6.curr_state_RNIVVMK_0_LC_9_15_0  (
            .in0(N__29472),
            .in1(N__29505),
            .in2(_gnd_net_),
            .in3(N__33906),
            .lcout(\b2v_inst6.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_7_1_0__m4_0_LC_9_15_1 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_7_1_0__m4_0_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_7_1_0__m4_0_LC_9_15_1 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \b2v_inst6.curr_state_7_1_0__m4_0_LC_9_15_1  (
            .in0(N__29533),
            .in1(N__34960),
            .in2(N__29515),
            .in3(N__29471),
            .lcout(),
            .ltout(G_2746_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNI7JCH_0_LC_9_15_2 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNI7JCH_0_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNI7JCH_0_LC_9_15_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.curr_state_RNI7JCH_0_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__29371),
            .in2(N__29377),
            .in3(N__33905),
            .lcout(\b2v_inst6.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst6.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_0_LC_9_15_3 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_0_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst6.curr_state_0_LC_9_15_3 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \b2v_inst6.curr_state_0_LC_9_15_3  (
            .in0(N__29534),
            .in1(N__34959),
            .in2(N__29374),
            .in3(N__29473),
            .lcout(\b2v_inst6.curr_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34676),
            .ce(N__33678),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIDMSJ1_0_1_LC_9_15_4 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIDMSJ1_0_1_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIDMSJ1_0_1_LC_9_15_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst6.curr_state_RNIDMSJ1_0_1_LC_9_15_4  (
            .in0(N__29721),
            .in1(N__29532),
            .in2(N__29707),
            .in3(N__29658),
            .lcout(\b2v_inst6.N_413 ),
            .ltout(\b2v_inst6.N_413_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_7_1_0__m6_0_LC_9_15_5 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_7_1_0__m6_0_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_7_1_0__m6_0_LC_9_15_5 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \b2v_inst6.curr_state_7_1_0__m6_0_LC_9_15_5  (
            .in0(N__29535),
            .in1(N__34942),
            .in2(N__29542),
            .in3(N__29514),
            .lcout(),
            .ltout(\b2v_inst6.curr_state_7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIF7P21_1_LC_9_15_6 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIF7P21_1_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIF7P21_1_LC_9_15_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.curr_state_RNIF7P21_1_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__29452),
            .in2(N__29539),
            .in3(N__33904),
            .lcout(\b2v_inst6.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst6.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_1_LC_9_15_7 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_1_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst6.curr_state_1_LC_9_15_7 .LUT_INIT=16'b0101010101000000;
    LogicCell40 \b2v_inst6.curr_state_1_LC_9_15_7  (
            .in0(N__29506),
            .in1(N__34941),
            .in2(N__29479),
            .in3(N__29474),
            .lcout(\b2v_inst6.curr_state_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34676),
            .ce(N__33678),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI471O_1_LC_11_1_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI471O_1_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI471O_1_LC_11_1_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNI471O_1_LC_11_1_0  (
            .in0(N__29401),
            .in1(N__31960),
            .in2(_gnd_net_),
            .in3(N__29443),
            .lcout(\b2v_inst36.countZ0Z_1 ),
            .ltout(\b2v_inst36.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI_1_LC_11_1_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI_1_LC_11_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI_1_LC_11_1_1 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \b2v_inst36.count_RNI_1_LC_11_1_1  (
            .in0(N__32236),
            .in1(_gnd_net_),
            .in2(N__29446),
            .in3(N__32143),
            .lcout(\b2v_inst36.count_rst_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI_15_LC_11_1_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI_15_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI_15_LC_11_1_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst36.count_RNI_15_LC_11_1_2  (
            .in0(N__29437),
            .in1(N__32235),
            .in2(N__31570),
            .in3(N__29419),
            .lcout(\b2v_inst36.un12_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_1_LC_11_1_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_1_LC_11_1_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_1_LC_11_1_3 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \b2v_inst36.count_1_LC_11_1_3  (
            .in0(N__32237),
            .in1(N__29810),
            .in2(_gnd_net_),
            .in3(N__32146),
            .lcout(\b2v_inst36.count_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34689),
            .ce(N__31962),
            .sr(N__31828));
    defparam \b2v_inst36.un2_count_1_cry_1_c_RNIAQA8_LC_11_1_4 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_1_c_RNIAQA8_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_1_c_RNIAQA8_LC_11_1_4 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_1_c_RNIAQA8_LC_11_1_4  (
            .in0(N__32144),
            .in1(N__32038),
            .in2(N__29941),
            .in3(N__29963),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIF2C01_2_LC_11_1_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIF2C01_2_LC_11_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIF2C01_2_LC_11_1_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst36.count_RNIF2C01_2_LC_11_1_5  (
            .in0(N__31961),
            .in1(_gnd_net_),
            .in2(N__29971),
            .in3(N__29920),
            .lcout(\b2v_inst36.countZ0Z_2 ),
            .ltout(\b2v_inst36.countZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_2_LC_11_1_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_2_LC_11_1_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_2_LC_11_1_6 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \b2v_inst36.count_2_LC_11_1_6  (
            .in0(N__32145),
            .in1(N__32042),
            .in2(N__29944),
            .in3(N__29940),
            .lcout(\b2v_inst36.count_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34689),
            .ce(N__31962),
            .sr(N__31828));
    defparam \b2v_inst36.count_3_LC_11_1_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_3_LC_11_1_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_3_LC_11_1_7 .LUT_INIT=16'b0000011000000000;
    LogicCell40 \b2v_inst36.count_3_LC_11_1_7  (
            .in0(N__29913),
            .in1(N__29887),
            .in2(N__32056),
            .in3(N__32147),
            .lcout(\b2v_inst36.count_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34689),
            .ce(N__31962),
            .sr(N__31828));
    defparam \b2v_inst36.count_RNI_0_1_LC_11_2_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI_0_1_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI_0_1_LC_11_2_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst36.count_RNI_0_1_LC_11_2_0  (
            .in0(N__29863),
            .in1(N__29842),
            .in2(N__29817),
            .in3(N__29741),
            .lcout(),
            .ltout(\b2v_inst36.un12_clk_100khz_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI9C1O_2_6_LC_11_2_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI9C1O_2_6_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI9C1O_2_6_LC_11_2_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst36.count_RNI9C1O_2_6_LC_11_2_1  (
            .in0(N__29791),
            .in1(N__30013),
            .in2(N__29779),
            .in3(N__29776),
            .lcout(\b2v_inst36.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_6_LC_11_2_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_6_LC_11_2_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_6_LC_11_2_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst36.count_6_LC_11_2_2  (
            .in0(N__30060),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.count_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34687),
            .ce(N__31977),
            .sr(N__31815));
    defparam \b2v_inst36.count_RNI9C1O_6_LC_11_2_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI9C1O_6_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI9C1O_6_LC_11_2_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNI9C1O_6_LC_11_2_3  (
            .in0(N__30042),
            .in1(N__31964),
            .in2(_gnd_net_),
            .in3(N__30059),
            .lcout(\b2v_inst36.un2_count_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIFGBV_11_LC_11_2_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIFGBV_11_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIFGBV_11_LC_11_2_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst36.count_RNIFGBV_11_LC_11_2_4  (
            .in0(N__31965),
            .in1(N__30070),
            .in2(_gnd_net_),
            .in3(N__29758),
            .lcout(\b2v_inst36.countZ0Z_11 ),
            .ltout(\b2v_inst36.countZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_11_LC_11_2_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_11_LC_11_2_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_11_LC_11_2_5 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst36.count_11_LC_11_2_5  (
            .in0(N__30091),
            .in1(N__32182),
            .in2(N__30073),
            .in3(N__32054),
            .lcout(\b2v_inst36.count_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34687),
            .ce(N__31977),
            .sr(N__31815));
    defparam \b2v_inst36.count_RNI9C1O_0_6_LC_11_2_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI9C1O_0_6_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI9C1O_0_6_LC_11_2_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst36.count_RNI9C1O_0_6_LC_11_2_6  (
            .in0(N__31966),
            .in1(_gnd_net_),
            .in2(N__30064),
            .in3(N__30043),
            .lcout(),
            .ltout(\b2v_inst36.countZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI9C1O_1_6_LC_11_2_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI9C1O_1_6_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI9C1O_1_6_LC_11_2_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst36.count_RNI9C1O_1_6_LC_11_2_7  (
            .in0(N__30034),
            .in1(N__31548),
            .in2(N__30016),
            .in3(N__30441),
            .lcout(\b2v_inst36.un12_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNI3NTL_1_LC_11_3_0 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI3NTL_1_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI3NTL_1_LC_11_3_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst36.curr_state_RNI3NTL_1_LC_11_3_0  (
            .in0(N__29983),
            .in1(N__29977),
            .in2(_gnd_net_),
            .in3(N__34073),
            .lcout(\b2v_inst36.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst36.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_7_1_0__m4_LC_11_3_1 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_7_1_0__m4_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_7_1_0__m4_LC_11_3_1 .LUT_INIT=16'b0011100000001000;
    LogicCell40 \b2v_inst36.curr_state_7_1_0__m4_LC_11_3_1  (
            .in0(N__30301),
            .in1(N__30389),
            .in2(N__30007),
            .in3(N__32034),
            .lcout(),
            .ltout(\b2v_inst36.curr_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNI2MTL_0_LC_11_3_2 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI2MTL_0_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI2MTL_0_LC_11_3_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.curr_state_RNI2MTL_0_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__30364),
            .in2(N__30004),
            .in3(N__34074),
            .lcout(\b2v_inst36.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst36.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.DSW_PWROK_LC_11_3_3 .C_ON=1'b0;
    defparam \b2v_inst36.DSW_PWROK_LC_11_3_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst36.DSW_PWROK_LC_11_3_3 .LUT_INIT=16'b0010000000100000;
    LogicCell40 \b2v_inst36.DSW_PWROK_LC_11_3_3  (
            .in0(N__30298),
            .in1(N__30336),
            .in2(N__30001),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.DSW_PWROK_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34684),
            .ce(N__33689),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_1_LC_11_3_4 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_1_LC_11_3_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst36.curr_state_1_LC_11_3_4 .LUT_INIT=16'b0010101000100000;
    LogicCell40 \b2v_inst36.curr_state_1_LC_11_3_4  (
            .in0(N__30257),
            .in1(N__32052),
            .in2(N__30349),
            .in3(N__30300),
            .lcout(\b2v_inst36.curr_state_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34684),
            .ce(N__33689),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_7_1_0__m6_LC_11_3_5 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_7_1_0__m6_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_7_1_0__m6_LC_11_3_5 .LUT_INIT=16'b0000100011001000;
    LogicCell40 \b2v_inst36.curr_state_7_1_0__m6_LC_11_3_5  (
            .in0(N__30302),
            .in1(N__30258),
            .in2(N__30353),
            .in3(N__32033),
            .lcout(\b2v_inst36.curr_state_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_0_LC_11_3_6 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_0_LC_11_3_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst36.curr_state_0_LC_11_3_6 .LUT_INIT=16'b0100010010100000;
    LogicCell40 \b2v_inst36.curr_state_0_LC_11_3_6  (
            .in0(N__30335),
            .in1(N__30299),
            .in2(N__32055),
            .in3(N__30388),
            .lcout(\b2v_inst36.curr_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34684),
            .ce(N__33689),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNI0A86_1_LC_11_3_7 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI0A86_1_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI0A86_1_LC_11_3_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst36.curr_state_RNI0A86_1_LC_11_3_7  (
            .in0(N__34075),
            .in1(N__30334),
            .in2(N__30307),
            .in3(N__30256),
            .lcout(\b2v_inst36.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_14_LC_11_4_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_14_LC_11_4_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_14_LC_11_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.count_14_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30775),
            .lcout(\b2v_inst5.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34679),
            .ce(N__32686),
            .sr(N__32867));
    defparam \b2v_inst5.count_6_LC_11_4_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_6_LC_11_4_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_6_LC_11_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.count_6_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30669),
            .lcout(\b2v_inst5.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34679),
            .ce(N__32686),
            .sr(N__32867));
    defparam \b2v_inst5.count_7_LC_11_4_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_7_LC_11_4_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_7_LC_11_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.count_7_LC_11_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30867),
            .lcout(\b2v_inst5.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34679),
            .ce(N__32686),
            .sr(N__32867));
    defparam \b2v_inst16.count_RNIPM3K1_8_LC_11_5_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIPM3K1_8_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIPM3K1_8_LC_11_5_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst16.count_RNIPM3K1_8_LC_11_5_0  (
            .in0(N__30174),
            .in1(N__30157),
            .in2(_gnd_net_),
            .in3(N__30603),
            .lcout(\b2v_inst16.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_8_LC_11_5_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_8_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_8_LC_11_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_8_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30175),
            .lcout(\b2v_inst16.count_4_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34672),
            .ce(N__30604),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIRP4K1_9_LC_11_5_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIRP4K1_9_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIRP4K1_9_LC_11_5_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst16.count_RNIRP4K1_9_LC_11_5_2  (
            .in0(N__30118),
            .in1(N__30097),
            .in2(_gnd_net_),
            .in3(N__30602),
            .lcout(\b2v_inst16.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_9_LC_11_5_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_9_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.count_9_LC_11_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_9_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30117),
            .lcout(\b2v_inst16.count_4_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34672),
            .ce(N__30604),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIJ8E01_4_LC_11_5_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIJ8E01_4_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIJ8E01_4_LC_11_5_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIJ8E01_4_LC_11_5_4  (
            .in0(N__30475),
            .in1(N__31963),
            .in2(_gnd_net_),
            .in3(N__30463),
            .lcout(\b2v_inst36.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI_0_0_LC_11_5_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI_0_0_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI_0_0_LC_11_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst5.count_RNI_0_0_LC_11_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32332),
            .lcout(\b2v_inst5.N_2906_i ),
            .ltout(\b2v_inst5.N_2906_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIU55SG_2_LC_11_5_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIU55SG_2_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIU55SG_2_LC_11_5_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \b2v_inst5.count_RNIU55SG_2_LC_11_5_6  (
            .in0(N__32443),
            .in1(_gnd_net_),
            .in2(N__30424),
            .in3(N__32302),
            .lcout(\b2v_inst5.N_390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIC5JH2_15_LC_11_5_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIC5JH2_15_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIC5JH2_15_LC_11_5_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst5.count_RNIC5JH2_15_LC_11_5_7  (
            .in0(N__32642),
            .in1(N__31153),
            .in2(_gnd_net_),
            .in3(N__31168),
            .lcout(\b2v_inst5.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_12_LC_11_6_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_12_LC_11_6_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_12_LC_11_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst5.count_12_LC_11_6_0  (
            .in0(N__30820),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34666),
            .ce(N__32680),
            .sr(N__32893));
    defparam \b2v_inst5.count_RNI6SFH2_12_LC_11_6_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI6SFH2_12_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI6SFH2_12_LC_11_6_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNI6SFH2_12_LC_11_6_1  (
            .in0(N__30417),
            .in1(N__32637),
            .in2(_gnd_net_),
            .in3(N__30818),
            .lcout(\b2v_inst5.un2_count_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIASDB2_0_5_LC_11_6_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIASDB2_0_5_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIASDB2_0_5_LC_11_6_2 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \b2v_inst5.count_RNIASDB2_0_5_LC_11_6_2  (
            .in0(N__32681),
            .in1(N__30754),
            .in2(N__30799),
            .in3(N__30703),
            .lcout(),
            .ltout(\b2v_inst5.count_1_i_a2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNISNC87_5_LC_11_6_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNISNC87_5_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNISNC87_5_LC_11_6_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst5.count_RNISNC87_5_LC_11_6_3  (
            .in0(N__30724),
            .in1(N__32509),
            .in2(N__30421),
            .in3(N__30409),
            .lcout(\b2v_inst5.count_1_i_a2_11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI6SFH2_0_12_LC_11_6_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI6SFH2_0_12_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI6SFH2_0_12_LC_11_6_4 .LUT_INIT=16'b0000000001010011;
    LogicCell40 \b2v_inst5.count_RNI6SFH2_0_12_LC_11_6_4  (
            .in0(N__30819),
            .in1(N__30418),
            .in2(N__32664),
            .in3(N__31182),
            .lcout(\b2v_inst5.count_1_i_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_5_LC_11_6_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_5_LC_11_6_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_5_LC_11_6_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst5.count_5_LC_11_6_5  (
            .in0(N__30702),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34666),
            .ce(N__32680),
            .sr(N__32893));
    defparam \b2v_inst5.count_RNIASDB2_5_LC_11_6_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIASDB2_5_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIASDB2_5_LC_11_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst5.count_RNIASDB2_5_LC_11_6_6  (
            .in0(N__32641),
            .in1(N__30753),
            .in2(_gnd_net_),
            .in3(N__30701),
            .lcout(\b2v_inst5.un2_count_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNICVEB2_0_6_LC_11_6_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNICVEB2_0_6_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNICVEB2_0_6_LC_11_6_7 .LUT_INIT=16'b0000000100001101;
    LogicCell40 \b2v_inst5.count_RNICVEB2_0_6_LC_11_6_7  (
            .in0(N__30744),
            .in1(N__32682),
            .in2(N__30895),
            .in3(N__30665),
            .lcout(\b2v_inst5.count_1_i_a2_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_1_c_LC_11_7_0 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_1_c_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_1_c_LC_11_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_1_c_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__32331),
            .in2(N__32398),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\b2v_inst5.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_1_c_RNIJQ1L1_LC_11_7_1 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_1_c_RNIJQ1L1_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_1_c_RNIJQ1L1_LC_11_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_1_c_RNIJQ1L1_LC_11_7_1  (
            .in0(N__32808),
            .in1(N__32404),
            .in2(_gnd_net_),
            .in3(N__30718),
            .lcout(\b2v_inst5.count_rst_12 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_1 ),
            .carryout(\b2v_inst5.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_11_7_2 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_11_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__32469),
            .in2(_gnd_net_),
            .in3(N__30715),
            .lcout(\b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_2 ),
            .carryout(\b2v_inst5.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_11_7_3 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_11_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__32997),
            .in2(_gnd_net_),
            .in3(N__30712),
            .lcout(\b2v_inst5.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_3 ),
            .carryout(\b2v_inst5.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_4_c_RNIM05L1_LC_11_7_4 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_4_c_RNIM05L1_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_4_c_RNIM05L1_LC_11_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_4_c_RNIM05L1_LC_11_7_4  (
            .in0(N__32803),
            .in1(N__30709),
            .in2(_gnd_net_),
            .in3(N__30691),
            .lcout(\b2v_inst5.count_rst_9 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_4 ),
            .carryout(\b2v_inst5.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_5_c_RNIN26L1_LC_11_7_5 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_5_c_RNIN26L1_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_5_c_RNIN26L1_LC_11_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_5_c_RNIN26L1_LC_11_7_5  (
            .in0(N__32809),
            .in1(N__30688),
            .in2(_gnd_net_),
            .in3(N__30646),
            .lcout(\b2v_inst5.count_rst_8 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_5 ),
            .carryout(\b2v_inst5.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_6_c_RNIO47L1_LC_11_7_6 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_6_c_RNIO47L1_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_6_c_RNIO47L1_LC_11_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_6_c_RNIO47L1_LC_11_7_6  (
            .in0(N__32802),
            .in1(N__30891),
            .in2(_gnd_net_),
            .in3(N__30847),
            .lcout(\b2v_inst5.count_rst_7 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_6 ),
            .carryout(\b2v_inst5.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_11_7_7 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_11_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__33046),
            .in2(_gnd_net_),
            .in3(N__30844),
            .lcout(\b2v_inst5.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_7 ),
            .carryout(\b2v_inst5.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_11_8_0 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_11_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__31750),
            .in2(_gnd_net_),
            .in3(N__30841),
            .lcout(\b2v_inst5.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\b2v_inst5.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_11_8_1 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_11_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__31705),
            .in2(_gnd_net_),
            .in3(N__30838),
            .lcout(\b2v_inst5.un2_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_9 ),
            .carryout(\b2v_inst5.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_10_c_RNI3GUD1_LC_11_8_2 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_10_c_RNI3GUD1_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_10_c_RNI3GUD1_LC_11_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_10_c_RNI3GUD1_LC_11_8_2  (
            .in0(N__32804),
            .in1(N__32347),
            .in2(_gnd_net_),
            .in3(N__30835),
            .lcout(\b2v_inst5.count_rst_3 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_10 ),
            .carryout(\b2v_inst5.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_11_c_RNI4IVD1_LC_11_8_3 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_11_c_RNI4IVD1_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_11_c_RNI4IVD1_LC_11_8_3 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_11_c_RNI4IVD1_LC_11_8_3  (
            .in0(N__32806),
            .in1(_gnd_net_),
            .in2(N__30832),
            .in3(N__30805),
            .lcout(\b2v_inst5.count_rst_2 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_11 ),
            .carryout(\b2v_inst5.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_11_8_4 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_11_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__32500),
            .in2(_gnd_net_),
            .in3(N__30802),
            .lcout(\b2v_inst5.un2_count_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_12 ),
            .carryout(\b2v_inst5.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_13_c_RNI6M1E1_LC_11_8_5 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_13_c_RNI6M1E1_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_13_c_RNI6M1E1_LC_11_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_13_c_RNI6M1E1_LC_11_8_5  (
            .in0(N__32807),
            .in1(N__30792),
            .in2(_gnd_net_),
            .in3(N__30757),
            .lcout(\b2v_inst5.count_rst_0 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_13 ),
            .carryout(\b2v_inst5.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_14_c_RNI7O2E1_LC_11_8_6 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_14_c_RNI7O2E1_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_14_c_RNI7O2E1_LC_11_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_14_c_RNI7O2E1_LC_11_8_6  (
            .in0(N__32805),
            .in1(N__31186),
            .in2(_gnd_net_),
            .in3(N__31171),
            .lcout(\b2v_inst5.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_15_LC_11_8_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_15_LC_11_8_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_15_LC_11_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.count_15_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31167),
            .lcout(\b2v_inst5.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34658),
            .ce(N__32679),
            .sr(N__32880));
    defparam \b2v_inst20.counter_1_cry_1_c_LC_11_9_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_1_c_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_1_c_LC_11_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.counter_1_cry_1_c_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__31144),
            .in2(N__31120),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\b2v_inst20.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_11_9_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_11_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__31087),
            .in2(_gnd_net_),
            .in3(N__31051),
            .lcout(\b2v_inst20.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_1 ),
            .carryout(\b2v_inst20.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_11_9_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_11_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__31048),
            .in2(_gnd_net_),
            .in3(N__31009),
            .lcout(\b2v_inst20.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_2 ),
            .carryout(\b2v_inst20.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_11_9_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_11_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__31006),
            .in2(_gnd_net_),
            .in3(N__30976),
            .lcout(\b2v_inst20.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_3 ),
            .carryout(\b2v_inst20.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_11_9_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_11_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__30973),
            .in2(_gnd_net_),
            .in3(N__30940),
            .lcout(\b2v_inst20.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_4 ),
            .carryout(\b2v_inst20.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_11_9_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_11_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__30937),
            .in2(_gnd_net_),
            .in3(N__30898),
            .lcout(\b2v_inst20.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_5 ),
            .carryout(\b2v_inst20.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_7_LC_11_9_6 .C_ON=1'b1;
    defparam \b2v_inst20.counter_7_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_7_LC_11_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_7_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__31227),
            .in2(_gnd_net_),
            .in3(N__31213),
            .lcout(\b2v_inst20.counterZ0Z_7 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_6 ),
            .carryout(\b2v_inst20.counter_1_cry_7 ),
            .clk(N__34652),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_8_LC_11_9_7 .C_ON=1'b1;
    defparam \b2v_inst20.counter_8_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_8_LC_11_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_8_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__33409),
            .in2(_gnd_net_),
            .in3(N__31210),
            .lcout(\b2v_inst20.counterZ0Z_8 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_7 ),
            .carryout(\b2v_inst20.counter_1_cry_8 ),
            .clk(N__34652),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_9_LC_11_10_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_9_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_9_LC_11_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_9_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__33382),
            .in2(_gnd_net_),
            .in3(N__31207),
            .lcout(\b2v_inst20.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\b2v_inst20.counter_1_cry_9 ),
            .clk(N__34657),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_10_LC_11_10_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_10_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_10_LC_11_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_10_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__33396),
            .in2(_gnd_net_),
            .in3(N__31204),
            .lcout(\b2v_inst20.counterZ0Z_10 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_9 ),
            .carryout(\b2v_inst20.counter_1_cry_10 ),
            .clk(N__34657),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_11_LC_11_10_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_11_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_11_LC_11_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_11_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__33421),
            .in2(_gnd_net_),
            .in3(N__31201),
            .lcout(\b2v_inst20.counterZ0Z_11 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_10 ),
            .carryout(\b2v_inst20.counter_1_cry_11 ),
            .clk(N__34657),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_12_LC_11_10_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_12_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_12_LC_11_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_12_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__33355),
            .in2(_gnd_net_),
            .in3(N__31198),
            .lcout(\b2v_inst20.counterZ0Z_12 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_11 ),
            .carryout(\b2v_inst20.counter_1_cry_12 ),
            .clk(N__34657),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_13_LC_11_10_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_13_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_13_LC_11_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_13_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__33316),
            .in2(_gnd_net_),
            .in3(N__31195),
            .lcout(\b2v_inst20.counterZ0Z_13 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_12 ),
            .carryout(\b2v_inst20.counter_1_cry_13 ),
            .clk(N__34657),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_14_LC_11_10_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_14_LC_11_10_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_14_LC_11_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_14_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__33343),
            .in2(_gnd_net_),
            .in3(N__31192),
            .lcout(\b2v_inst20.counterZ0Z_14 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_13 ),
            .carryout(\b2v_inst20.counter_1_cry_14 ),
            .clk(N__34657),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_15_LC_11_10_6 .C_ON=1'b1;
    defparam \b2v_inst20.counter_15_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_15_LC_11_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_15_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__33330),
            .in2(_gnd_net_),
            .in3(N__31189),
            .lcout(\b2v_inst20.counterZ0Z_15 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_14 ),
            .carryout(\b2v_inst20.counter_1_cry_15 ),
            .clk(N__34657),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_16_LC_11_10_7 .C_ON=1'b1;
    defparam \b2v_inst20.counter_16_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_16_LC_11_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_16_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__33280),
            .in2(_gnd_net_),
            .in3(N__31258),
            .lcout(\b2v_inst20.counterZ0Z_16 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_15 ),
            .carryout(\b2v_inst20.counter_1_cry_16 ),
            .clk(N__34657),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_17_LC_11_11_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_17_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_17_LC_11_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_17_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__33267),
            .in2(_gnd_net_),
            .in3(N__31255),
            .lcout(\b2v_inst20.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\b2v_inst20.counter_1_cry_17 ),
            .clk(N__34663),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_18_LC_11_11_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_18_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_18_LC_11_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_18_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__33253),
            .in2(_gnd_net_),
            .in3(N__31252),
            .lcout(\b2v_inst20.counterZ0Z_18 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_17 ),
            .carryout(\b2v_inst20.counter_1_cry_18 ),
            .clk(N__34663),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_19_LC_11_11_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_19_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_19_LC_11_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_19_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__33292),
            .in2(_gnd_net_),
            .in3(N__31249),
            .lcout(\b2v_inst20.counterZ0Z_19 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_18 ),
            .carryout(\b2v_inst20.counter_1_cry_19 ),
            .clk(N__34663),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_20_LC_11_11_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_20_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_20_LC_11_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_20_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__33187),
            .in2(_gnd_net_),
            .in3(N__31246),
            .lcout(\b2v_inst20.counterZ0Z_20 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_19 ),
            .carryout(\b2v_inst20.counter_1_cry_20 ),
            .clk(N__34663),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_21_LC_11_11_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_21_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_21_LC_11_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_21_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__33201),
            .in2(_gnd_net_),
            .in3(N__31243),
            .lcout(\b2v_inst20.counterZ0Z_21 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_20 ),
            .carryout(\b2v_inst20.counter_1_cry_21 ),
            .clk(N__34663),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_22_LC_11_11_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_22_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_22_LC_11_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_22_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__33214),
            .in2(_gnd_net_),
            .in3(N__31240),
            .lcout(\b2v_inst20.counterZ0Z_22 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_21 ),
            .carryout(\b2v_inst20.counter_1_cry_22 ),
            .clk(N__34663),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_23_LC_11_11_6 .C_ON=1'b1;
    defparam \b2v_inst20.counter_23_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_23_LC_11_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_23_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__33226),
            .in2(_gnd_net_),
            .in3(N__31237),
            .lcout(\b2v_inst20.counterZ0Z_23 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_22 ),
            .carryout(\b2v_inst20.counter_1_cry_23 ),
            .clk(N__34663),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_24_LC_11_11_7 .C_ON=1'b1;
    defparam \b2v_inst20.counter_24_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_24_LC_11_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_24_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(N__33160),
            .in2(_gnd_net_),
            .in3(N__31234),
            .lcout(\b2v_inst20.counterZ0Z_24 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_23 ),
            .carryout(\b2v_inst20.counter_1_cry_24 ),
            .clk(N__34663),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_25_LC_11_12_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_25_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_25_LC_11_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_25_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__33129),
            .in2(_gnd_net_),
            .in3(N__31282),
            .lcout(\b2v_inst20.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\b2v_inst20.counter_1_cry_25 ),
            .clk(N__34665),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_26_LC_11_12_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_26_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_26_LC_11_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_26_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__33114),
            .in2(_gnd_net_),
            .in3(N__31279),
            .lcout(\b2v_inst20.counterZ0Z_26 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_25 ),
            .carryout(\b2v_inst20.counter_1_cry_26 ),
            .clk(N__34665),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_27_LC_11_12_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_27_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_27_LC_11_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_27_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__33147),
            .in2(_gnd_net_),
            .in3(N__31276),
            .lcout(\b2v_inst20.counterZ0Z_27 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_26 ),
            .carryout(\b2v_inst20.counter_1_cry_27 ),
            .clk(N__34665),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_28_LC_11_12_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_28_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_28_LC_11_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_28_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__33472),
            .in2(_gnd_net_),
            .in3(N__31273),
            .lcout(\b2v_inst20.counterZ0Z_28 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_27 ),
            .carryout(\b2v_inst20.counter_1_cry_28 ),
            .clk(N__34665),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_29_LC_11_12_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_29_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_29_LC_11_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_29_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(N__33484),
            .in2(_gnd_net_),
            .in3(N__31270),
            .lcout(\b2v_inst20.counterZ0Z_29 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_28 ),
            .carryout(\b2v_inst20.counter_1_cry_29 ),
            .clk(N__34665),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_30_LC_11_12_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_30_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_30_LC_11_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_30_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(N__33445),
            .in2(_gnd_net_),
            .in3(N__31267),
            .lcout(\b2v_inst20.counterZ0Z_30 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_29 ),
            .carryout(\b2v_inst20.counter_1_cry_30 ),
            .clk(N__34665),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_31_LC_11_12_6 .C_ON=1'b0;
    defparam \b2v_inst20.counter_31_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_31_LC_11_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst20.counter_31_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__33459),
            .in2(_gnd_net_),
            .in3(N__31264),
            .lcout(\b2v_inst20.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34665),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_1_c_LC_11_13_0 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_1_c_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_1_c_LC_11_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_1_c_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__34214),
            .in2(N__35026),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\b2v_inst6.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNIM2GO_LC_11_13_1 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNIM2GO_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNIM2GO_LC_11_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_1_c_RNIM2GO_LC_11_13_1  (
            .in0(N__35273),
            .in1(N__34230),
            .in2(_gnd_net_),
            .in3(N__31261),
            .lcout(\b2v_inst6.count_rst_1 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_1 ),
            .carryout(\b2v_inst6.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_13_2 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__35093),
            .in2(_gnd_net_),
            .in3(N__31336),
            .lcout(\b2v_inst6.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_2 ),
            .carryout(\b2v_inst6.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_13_3 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__35058),
            .in2(_gnd_net_),
            .in3(N__31318),
            .lcout(\b2v_inst6.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_3 ),
            .carryout(\b2v_inst6.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_13_4 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__35126),
            .in2(_gnd_net_),
            .in3(N__31315),
            .lcout(\b2v_inst6.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_4 ),
            .carryout(\b2v_inst6.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_5_c_RNIQAKO_LC_11_13_5 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_5_c_RNIQAKO_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_5_c_RNIQAKO_LC_11_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_5_c_RNIQAKO_LC_11_13_5  (
            .in0(N__35274),
            .in1(N__34255),
            .in2(_gnd_net_),
            .in3(N__31312),
            .lcout(\b2v_inst6.count_rst_5 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_5 ),
            .carryout(\b2v_inst6.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_13_6 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__31455),
            .in2(_gnd_net_),
            .in3(N__31309),
            .lcout(\b2v_inst6.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_6 ),
            .carryout(\b2v_inst6.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_13_7 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__31410),
            .in2(_gnd_net_),
            .in3(N__31306),
            .lcout(\b2v_inst6.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_7 ),
            .carryout(\b2v_inst6.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_14_0 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__31633),
            .in2(_gnd_net_),
            .in3(N__31303),
            .lcout(\b2v_inst6.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\b2v_inst6.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNIUIOO_LC_11_14_1 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNIUIOO_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNIUIOO_LC_11_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_9_c_RNIUIOO_LC_11_14_1  (
            .in0(N__35290),
            .in1(N__34242),
            .in2(_gnd_net_),
            .in3(N__31300),
            .lcout(\b2v_inst6.count_rst_9 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_9 ),
            .carryout(\b2v_inst6.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_14_2 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__31484),
            .in2(_gnd_net_),
            .in3(N__31285),
            .lcout(\b2v_inst6.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_10 ),
            .carryout(\b2v_inst6.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNI7R101_LC_11_14_3 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNI7R101_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNI7R101_LC_11_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_11_c_RNI7R101_LC_11_14_3  (
            .in0(N__35291),
            .in1(N__34200),
            .in2(_gnd_net_),
            .in3(N__31390),
            .lcout(\b2v_inst6.count_rst_11 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_11 ),
            .carryout(\b2v_inst6.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNI8T201_LC_11_14_4 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNI8T201_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNI8T201_LC_11_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_12_c_RNI8T201_LC_11_14_4  (
            .in0(N__35296),
            .in1(N__34173),
            .in2(_gnd_net_),
            .in3(N__31387),
            .lcout(\b2v_inst6.count_rst_12 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_12 ),
            .carryout(\b2v_inst6.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_13_c_RNI9V301_LC_11_14_5 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_13_c_RNI9V301_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_13_c_RNI9V301_LC_11_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_13_c_RNI9V301_LC_11_14_5  (
            .in0(N__35292),
            .in1(N__34848),
            .in2(_gnd_net_),
            .in3(N__31384),
            .lcout(\b2v_inst6.count_rst_13 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_13 ),
            .carryout(\b2v_inst6.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_14_c_RNIA1501_LC_11_14_6 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_14_c_RNIA1501_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_14_c_RNIA1501_LC_11_14_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_14_c_RNIA1501_LC_11_14_6  (
            .in0(N__34803),
            .in1(N__35293),
            .in2(_gnd_net_),
            .in3(N__31381),
            .lcout(\b2v_inst6.count_rst_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_15_LC_11_14_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_15_LC_11_14_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_15_LC_11_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.count_15_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34816),
            .lcout(\b2v_inst6.count_3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34678),
            .ce(N__34430),
            .sr(N__35297));
    defparam \b2v_inst6.un2_count_1_cry_4_c_RNIP8JO_LC_11_15_0 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_4_c_RNIP8JO_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_4_c_RNIP8JO_LC_11_15_0 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_4_c_RNIP8JO_LC_11_15_0  (
            .in0(N__34895),
            .in1(N__31371),
            .in2(N__35130),
            .in3(N__35226),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI1N0E4_5_LC_11_15_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI1N0E4_5_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI1N0E4_5_LC_11_15_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst6.count_RNI1N0E4_5_LC_11_15_1  (
            .in0(N__34370),
            .in1(_gnd_net_),
            .in2(N__31354),
            .in3(N__31351),
            .lcout(\b2v_inst6.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_2_c_RNIN4HO_LC_11_15_2 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_2_c_RNIN4HO_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_2_c_RNIN4HO_LC_11_15_2 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_2_c_RNIN4HO_LC_11_15_2  (
            .in0(N__34894),
            .in1(N__34716),
            .in2(N__35095),
            .in3(N__35225),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNITGUD4_3_LC_11_15_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNITGUD4_3_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNITGUD4_3_LC_11_15_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst6.count_RNITGUD4_3_LC_11_15_3  (
            .in0(N__34369),
            .in1(_gnd_net_),
            .in2(N__31339),
            .in3(N__34699),
            .lcout(\b2v_inst6.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_8_c_RNITGNO_LC_11_15_4 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_8_c_RNITGNO_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_8_c_RNITGNO_LC_11_15_4 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_8_c_RNITGNO_LC_11_15_4  (
            .in0(N__34896),
            .in1(N__31611),
            .in2(N__31639),
            .in3(N__35227),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI935E4_9_LC_11_15_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI935E4_9_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI935E4_9_LC_11_15_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst6.count_RNI935E4_9_LC_11_15_5  (
            .in0(N__34371),
            .in1(_gnd_net_),
            .in2(N__31510),
            .in3(N__31600),
            .lcout(\b2v_inst6.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIIEMF4_10_LC_11_15_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIIEMF4_10_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIIEMF4_10_LC_11_15_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNIIEMF4_10_LC_11_15_6  (
            .in0(N__31498),
            .in1(N__31506),
            .in2(_gnd_net_),
            .in3(N__34372),
            .lcout(\b2v_inst6.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_10_LC_11_15_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_10_LC_11_15_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_10_LC_11_15_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst6.count_10_LC_11_15_7  (
            .in0(N__31507),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.count_3_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34683),
            .ce(N__34420),
            .sr(N__35294));
    defparam \b2v_inst6.count_RNI_7_LC_11_16_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_7_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_7_LC_11_16_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst6.count_RNI_7_LC_11_16_0  (
            .in0(N__31406),
            .in1(N__31634),
            .in2(N__31456),
            .in3(N__31489),
            .lcout(\b2v_inst6.un12_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_6_c_RNIRCLO_LC_11_16_1 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_6_c_RNIRCLO_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_6_c_RNIRCLO_LC_11_16_1 .LUT_INIT=16'b0000000001100000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_6_c_RNIRCLO_LC_11_16_1  (
            .in0(N__31434),
            .in1(N__31454),
            .in2(N__34928),
            .in3(N__35275),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI5T2E4_7_LC_11_16_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI5T2E4_7_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI5T2E4_7_LC_11_16_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNI5T2E4_7_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__31420),
            .in2(N__31459),
            .in3(N__34418),
            .lcout(\b2v_inst6.countZ0Z_7 ),
            .ltout(\b2v_inst6.countZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_7_LC_11_16_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_7_LC_11_16_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_7_LC_11_16_3 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst6.count_7_LC_11_16_3  (
            .in0(N__31435),
            .in1(N__34935),
            .in2(N__31423),
            .in3(N__35278),
            .lcout(\b2v_inst6.count_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34686),
            .ce(N__34434),
            .sr(N__35307));
    defparam \b2v_inst6.un2_count_1_cry_7_c_RNISEMO_LC_11_16_4 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_7_c_RNISEMO_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_7_c_RNISEMO_LC_11_16_4 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_7_c_RNISEMO_LC_11_16_4  (
            .in0(N__35276),
            .in1(N__31656),
            .in2(N__31411),
            .in3(N__34903),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI704E4_8_LC_11_16_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI704E4_8_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI704E4_8_LC_11_16_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst6.count_RNI704E4_8_LC_11_16_5  (
            .in0(N__34419),
            .in1(_gnd_net_),
            .in2(N__31414),
            .in3(N__31645),
            .lcout(\b2v_inst6.countZ0Z_8 ),
            .ltout(\b2v_inst6.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_8_LC_11_16_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_8_LC_11_16_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_8_LC_11_16_6 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst6.count_8_LC_11_16_6  (
            .in0(N__35277),
            .in1(N__34904),
            .in2(N__31660),
            .in3(N__31657),
            .lcout(\b2v_inst6.count_3_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34686),
            .ce(N__34434),
            .sr(N__35307));
    defparam \b2v_inst6.count_9_LC_11_16_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_9_LC_11_16_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_9_LC_11_16_7 .LUT_INIT=16'b0000000001100000;
    LogicCell40 \b2v_inst6.count_9_LC_11_16_7  (
            .in0(N__31635),
            .in1(N__31615),
            .in2(N__34929),
            .in3(N__35279),
            .lcout(\b2v_inst6.count_3_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34686),
            .ce(N__34434),
            .sr(N__35307));
    defparam \b2v_inst36.count_RNI_0_LC_12_1_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI_0_LC_12_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI_0_LC_12_1_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst36.count_RNI_0_LC_12_1_0  (
            .in0(N__32241),
            .in1(N__32181),
            .in2(_gnd_net_),
            .in3(N__32051),
            .lcout(\b2v_inst36.count_rst_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNI_1_LC_12_2_0 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI_1_LC_12_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI_1_LC_12_2_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst36.curr_state_RNI_1_LC_12_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31785),
            .lcout(\b2v_inst36.N_2928_i ),
            .ltout(\b2v_inst36.N_2928_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_13_LC_12_2_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_13_LC_12_2_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_13_LC_12_2_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \b2v_inst36.count_13_LC_12_2_1  (
            .in0(N__31582),
            .in1(_gnd_net_),
            .in2(N__31591),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.count_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34690),
            .ce(N__31975),
            .sr(N__31836));
    defparam \b2v_inst36.count_RNIJMDV_13_LC_12_2_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIJMDV_13_LC_12_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIJMDV_13_LC_12_2_2 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \b2v_inst36.count_RNIJMDV_13_LC_12_2_2  (
            .in0(N__32178),
            .in1(N__31588),
            .in2(N__31978),
            .in3(N__31581),
            .lcout(\b2v_inst36.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNITNJ01_9_LC_12_2_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNITNJ01_9_LC_12_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNITNJ01_9_LC_12_2_3 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \b2v_inst36.count_RNITNJ01_9_LC_12_2_3  (
            .in0(N__31516),
            .in1(N__31970),
            .in2(N__31534),
            .in3(N__32177),
            .lcout(\b2v_inst36.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_9_LC_12_2_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_9_LC_12_2_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_9_LC_12_2_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst36.count_9_LC_12_2_4  (
            .in0(N__32179),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31530),
            .lcout(\b2v_inst36.count_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34690),
            .ce(N__31975),
            .sr(N__31836));
    defparam \b2v_inst36.count_RNI361O_0_LC_12_2_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI361O_0_LC_12_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI361O_0_LC_12_2_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst36.count_RNI361O_0_LC_12_2_6  (
            .in0(N__31974),
            .in1(N__32251),
            .in2(_gnd_net_),
            .in3(N__31984),
            .lcout(\b2v_inst36.countZ0Z_0 ),
            .ltout(\b2v_inst36.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_0_LC_12_2_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_0_LC_12_2_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_0_LC_12_2_7 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \b2v_inst36.count_0_LC_12_2_7  (
            .in0(_gnd_net_),
            .in1(N__32180),
            .in2(N__32092),
            .in3(N__32053),
            .lcout(\b2v_inst36.count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34690),
            .ce(N__31975),
            .sr(N__31836));
    defparam \b2v_inst5.count_RNII8IB2_0_9_LC_12_5_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNII8IB2_0_9_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNII8IB2_0_9_LC_12_5_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \b2v_inst5.count_RNII8IB2_0_9_LC_12_5_0  (
            .in0(N__31697),
            .in1(N__31759),
            .in2(N__32678),
            .in3(N__31717),
            .lcout(\b2v_inst5.count_1_i_a2_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_8_c_RNIQ89L1_LC_12_5_1 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_8_c_RNIQ89L1_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_8_c_RNIQ89L1_LC_12_5_1 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_8_c_RNIQ89L1_LC_12_5_1  (
            .in0(N__31731),
            .in1(N__31743),
            .in2(N__32883),
            .in3(N__32946),
            .lcout(\b2v_inst5.count_rst_5 ),
            .ltout(\b2v_inst5.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNII8IB2_9_LC_12_5_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNII8IB2_9_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNII8IB2_9_LC_12_5_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \b2v_inst5.count_RNII8IB2_9_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(N__32650),
            .in2(N__31753),
            .in3(N__31716),
            .lcout(\b2v_inst5.un2_count_1_axb_9 ),
            .ltout(\b2v_inst5.un2_count_1_axb_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_9_LC_12_5_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_9_LC_12_5_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_9_LC_12_5_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.count_9_LC_12_5_3  (
            .in0(N__31732),
            .in1(N__32866),
            .in2(N__31720),
            .in3(N__32950),
            .lcout(\b2v_inst5.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34681),
            .ce(N__32660),
            .sr(N__32892));
    defparam \b2v_inst5.un2_count_1_cry_9_c_RNIRAAL1_LC_12_5_4 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_9_c_RNIRAAL1_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_9_c_RNIRAAL1_LC_12_5_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_9_c_RNIRAAL1_LC_12_5_4  (
            .in0(N__32947),
            .in1(N__32861),
            .in2(N__31704),
            .in3(N__31680),
            .lcout(),
            .ltout(\b2v_inst5.count_rst_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIRIQO2_10_LC_12_5_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIRIQO2_10_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIRIQO2_10_LC_12_5_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst5.count_RNIRIQO2_10_LC_12_5_5  (
            .in0(N__32651),
            .in1(_gnd_net_),
            .in2(N__31708),
            .in3(N__31666),
            .lcout(\b2v_inst5.countZ0Z_10 ),
            .ltout(\b2v_inst5.countZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_10_LC_12_5_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_10_LC_12_5_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_10_LC_12_5_6 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst5.count_10_LC_12_5_6  (
            .in0(N__32948),
            .in1(N__32865),
            .in2(N__31684),
            .in3(N__31681),
            .lcout(\b2v_inst5.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34681),
            .ce(N__32660),
            .sr(N__32892));
    defparam \b2v_inst5.count_13_LC_12_5_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_13_LC_12_5_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_13_LC_12_5_7 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \b2v_inst5.count_13_LC_12_5_7  (
            .in0(N__32504),
            .in1(N__32908),
            .in2(N__32884),
            .in3(N__32949),
            .lcout(\b2v_inst5.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34681),
            .ce(N__32660),
            .sr(N__32892));
    defparam \b2v_inst5.count_RNIRHC7I_2_LC_12_6_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIRHC7I_2_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIRHC7I_2_LC_12_6_0 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \b2v_inst5.count_RNIRHC7I_2_LC_12_6_0  (
            .in0(N__32297),
            .in1(N__32442),
            .in2(N__32868),
            .in3(N__32284),
            .lcout(),
            .ltout(\b2v_inst5.count_RNIRHC7IZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIA8LTI_0_LC_12_6_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIA8LTI_0_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIA8LTI_0_LC_12_6_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst5.count_RNIA8LTI_0_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__32275),
            .in2(N__32335),
            .in3(N__32643),
            .lcout(\b2v_inst5.countZ0Z_0 ),
            .ltout(\b2v_inst5.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI_0_LC_12_6_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI_0_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI_0_LC_12_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst5.count_RNI_0_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32320),
            .in3(N__32397),
            .lcout(\b2v_inst5.count_RNIZ0Z_0 ),
            .ltout(\b2v_inst5.count_RNIZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNID3G12_1_LC_12_6_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNID3G12_1_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNID3G12_1_LC_12_6_3 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst5.count_RNID3G12_1_LC_12_6_3  (
            .in0(N__32832),
            .in1(N__32308),
            .in2(N__32317),
            .in3(N__32644),
            .lcout(\b2v_inst5.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_1_LC_12_6_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_1_LC_12_6_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_1_LC_12_6_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst5.count_1_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__32314),
            .in2(_gnd_net_),
            .in3(N__32834),
            .lcout(\b2v_inst5.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34674),
            .ce(N__32646),
            .sr(N__32882));
    defparam \b2v_inst5.count_3_LC_12_6_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_3_LC_12_6_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_3_LC_12_6_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst5.count_3_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__32828),
            .in2(_gnd_net_),
            .in3(N__32260),
            .lcout(\b2v_inst5.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34674),
            .ce(N__32646),
            .sr(N__32882));
    defparam \b2v_inst5.count_0_LC_12_6_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_0_LC_12_6_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_0_LC_12_6_6 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \b2v_inst5.count_0_LC_12_6_6  (
            .in0(N__32298),
            .in1(N__32283),
            .in2(N__32869),
            .in3(N__32441),
            .lcout(\b2v_inst5.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34674),
            .ce(N__32646),
            .sr(N__32882));
    defparam \b2v_inst5.count_RNI6MBB2_3_LC_12_6_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI6MBB2_3_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI6MBB2_3_LC_12_6_7 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \b2v_inst5.count_RNI6MBB2_3_LC_12_6_7  (
            .in0(N__32833),
            .in1(N__32645),
            .in2(N__32269),
            .in3(N__32259),
            .lcout(\b2v_inst5.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_2_LC_12_7_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_2_LC_12_7_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_2_LC_12_7_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst5.count_2_LC_12_7_0  (
            .in0(N__32416),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34668),
            .ce(N__32635),
            .sr(N__32885));
    defparam \b2v_inst5.count_RNI4JAB2_0_2_LC_12_7_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI4JAB2_0_2_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI4JAB2_0_2_LC_12_7_1 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \b2v_inst5.count_RNI4JAB2_0_2_LC_12_7_1  (
            .in0(N__32633),
            .in1(N__32425),
            .in2(N__32473),
            .in3(N__32415),
            .lcout(),
            .ltout(\b2v_inst5.count_1_i_a2_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI2EOJ9_2_LC_12_7_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI2EOJ9_2_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI2EOJ9_2_LC_12_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst5.count_RNI2EOJ9_2_LC_12_7_2  (
            .in0(N__32455),
            .in1(N__32341),
            .in2(N__32446),
            .in3(N__32377),
            .lcout(\b2v_inst5.count_1_i_a2_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI4JAB2_2_LC_12_7_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI4JAB2_2_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI4JAB2_2_LC_12_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst5.count_RNI4JAB2_2_LC_12_7_3  (
            .in0(N__32632),
            .in1(N__32424),
            .in2(_gnd_net_),
            .in3(N__32414),
            .lcout(\b2v_inst5.un2_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI4PEH2_0_11_LC_12_7_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI4PEH2_0_11_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI4PEH2_0_11_LC_12_7_4 .LUT_INIT=16'b0000000000100111;
    LogicCell40 \b2v_inst5.count_RNI4PEH2_0_11_LC_12_7_4  (
            .in0(N__32634),
            .in1(N__32358),
            .in2(N__32371),
            .in3(N__32396),
            .lcout(\b2v_inst5.count_1_i_a2_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_11_LC_12_7_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_11_LC_12_7_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_11_LC_12_7_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst5.count_11_LC_12_7_5  (
            .in0(N__32359),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34668),
            .ce(N__32635),
            .sr(N__32885));
    defparam \b2v_inst5.count_RNI4PEH2_11_LC_12_7_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI4PEH2_11_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI4PEH2_11_LC_12_7_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNI4PEH2_11_LC_12_7_6  (
            .in0(N__32367),
            .in1(N__32631),
            .in2(_gnd_net_),
            .in3(N__32357),
            .lcout(\b2v_inst5.un2_count_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI8PCB2_0_4_LC_12_7_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI8PCB2_0_4_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI8PCB2_0_4_LC_12_7_7 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \b2v_inst5.count_RNI8PCB2_0_4_LC_12_7_7  (
            .in0(N__33045),
            .in1(N__33010),
            .in2(N__32974),
            .in3(N__32636),
            .lcout(\b2v_inst5.count_1_i_a2_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_7_c_RNIP68L1_LC_12_8_0 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_7_c_RNIP68L1_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_7_c_RNIP68L1_LC_12_8_0 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_7_c_RNIP68L1_LC_12_8_0  (
            .in0(N__32953),
            .in1(N__33027),
            .in2(N__32870),
            .in3(N__33044),
            .lcout(),
            .ltout(\b2v_inst5.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIG5HB2_8_LC_12_8_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIG5HB2_8_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIG5HB2_8_LC_12_8_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst5.count_RNIG5HB2_8_LC_12_8_1  (
            .in0(N__32649),
            .in1(_gnd_net_),
            .in2(N__33049),
            .in3(N__33016),
            .lcout(\b2v_inst5.countZ0Z_8 ),
            .ltout(\b2v_inst5.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_8_LC_12_8_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_8_LC_12_8_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_8_LC_12_8_2 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst5.count_8_LC_12_8_2  (
            .in0(N__32955),
            .in1(N__33028),
            .in2(N__33019),
            .in3(N__32841),
            .lcout(\b2v_inst5.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34664),
            .ce(N__32659),
            .sr(N__32881));
    defparam \b2v_inst5.un2_count_1_cry_3_c_RNILU3L1_LC_12_8_3 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_3_c_RNILU3L1_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_3_c_RNILU3L1_LC_12_8_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.un2_count_1_cry_3_c_RNILU3L1_LC_12_8_3  (
            .in0(N__32985),
            .in1(N__32951),
            .in2(N__33001),
            .in3(N__32835),
            .lcout(\b2v_inst5.count_rst_10 ),
            .ltout(\b2v_inst5.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI8PCB2_4_LC_12_8_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI8PCB2_4_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI8PCB2_4_LC_12_8_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst5.count_RNI8PCB2_4_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(N__32970),
            .in2(N__33004),
            .in3(N__32647),
            .lcout(\b2v_inst5.un2_count_1_axb_4 ),
            .ltout(\b2v_inst5.un2_count_1_axb_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_4_LC_12_8_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_4_LC_12_8_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_4_LC_12_8_5 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.count_4_LC_12_8_5  (
            .in0(N__32986),
            .in1(N__32954),
            .in2(N__32977),
            .in3(N__32839),
            .lcout(\b2v_inst5.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34664),
            .ce(N__32659),
            .sr(N__32881));
    defparam \b2v_inst5.un2_count_1_cry_12_c_RNI5K0E1_LC_12_8_6 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_12_c_RNI5K0E1_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_12_c_RNI5K0E1_LC_12_8_6 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_12_c_RNI5K0E1_LC_12_8_6  (
            .in0(N__32952),
            .in1(N__32904),
            .in2(N__32505),
            .in3(N__32840),
            .lcout(),
            .ltout(\b2v_inst5.count_rst_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI8VGH2_13_LC_12_8_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI8VGH2_13_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI8VGH2_13_LC_12_8_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst5.count_RNI8VGH2_13_LC_12_8_7  (
            .in0(N__32648),
            .in1(_gnd_net_),
            .in2(N__32521),
            .in3(N__32518),
            .lcout(\b2v_inst5.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_2_LC_12_9_3 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_2_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.curr_state_2_LC_12_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst200.curr_state_2_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34114),
            .lcout(\b2v_inst200.curr_state_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34656),
            .ce(N__33686),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_2_c_RNO_LC_12_10_0 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_2_c_RNO_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_2_c_RNO_LC_12_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_2_c_RNO_LC_12_10_0  (
            .in0(N__33420),
            .in1(N__33408),
            .in2(N__33397),
            .in3(N__33381),
            .lcout(\b2v_inst20.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_3_c_RNO_LC_12_10_1 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_3_c_RNO_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_3_c_RNO_LC_12_10_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_3_c_RNO_LC_12_10_1  (
            .in0(N__33354),
            .in1(N__33342),
            .in2(N__33331),
            .in3(N__33315),
            .lcout(\b2v_inst20.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_4_c_RNO_LC_12_10_2 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_4_c_RNO_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_4_c_RNO_LC_12_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_4_c_RNO_LC_12_10_2  (
            .in0(N__33291),
            .in1(N__33279),
            .in2(N__33268),
            .in3(N__33252),
            .lcout(\b2v_inst20.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_5_c_RNO_LC_12_10_3 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_5_c_RNO_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_5_c_RNO_LC_12_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_5_c_RNO_LC_12_10_3  (
            .in0(N__33225),
            .in1(N__33213),
            .in2(N__33202),
            .in3(N__33186),
            .lcout(\b2v_inst20.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_6_c_RNO_LC_12_10_4 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_6_c_RNO_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_6_c_RNO_LC_12_10_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_6_c_RNO_LC_12_10_4  (
            .in0(N__33159),
            .in1(N__33148),
            .in2(N__33133),
            .in3(N__33115),
            .lcout(\b2v_inst20.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNIQ7EG4_1_LC_12_11_0 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNIQ7EG4_1_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNIQ7EG4_1_LC_12_11_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.curr_state_RNIQ7EG4_1_LC_12_11_0  (
            .in0(N__33514),
            .in1(N__33532),
            .in2(_gnd_net_),
            .in3(N__34069),
            .lcout(\b2v_inst200.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst200.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_12_11_1 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_12_11_1 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33085),
            .in3(N__33821),
            .lcout(N_405),
            .ltout(N_405_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_12_11_2 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_12_11_2 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_12_11_2  (
            .in0(N__33622),
            .in1(N__33616),
            .in2(N__33547),
            .in3(N__33522),
            .lcout(\b2v_inst200.m6_i_0 ),
            .ltout(\b2v_inst200.m6_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_LC_12_11_3 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_LC_12_11_3 .LUT_INIT=16'b1111010011110001;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m6_i_LC_12_11_3  (
            .in0(N__33768),
            .in1(N__33802),
            .in2(N__33544),
            .in3(N__33822),
            .lcout(),
            .ltout(\b2v_inst200.N_57_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNIKHBJ4_0_LC_12_11_4 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNIKHBJ4_0_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNIKHBJ4_0_LC_12_11_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst200.curr_state_RNIKHBJ4_0_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__33724),
            .in2(N__33541),
            .in3(N__34070),
            .lcout(\b2v_inst200.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst200.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_a2_LC_12_11_5 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_a2_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_a2_LC_12_11_5 .LUT_INIT=16'b0000110000001100;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m8_i_a2_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__33803),
            .in2(N__33538),
            .in3(_gnd_net_),
            .lcout(N_406),
            .ltout(N_406_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_LC_12_11_6 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_LC_12_11_6 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m8_i_LC_12_11_6  (
            .in0(N__33805),
            .in1(N__34147),
            .in2(N__33535),
            .in3(N__33767),
            .lcout(\b2v_inst200.N_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_1_LC_12_11_7 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_1_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.curr_state_1_LC_12_11_7 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \b2v_inst200.curr_state_1_LC_12_11_7  (
            .in0(N__33769),
            .in1(N__33804),
            .in2(N__33526),
            .in3(N__34146),
            .lcout(\b2v_inst200.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34667),
            .ce(N__33683),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNI_0_LC_12_12_0 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNI_0_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNI_0_LC_12_12_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \b2v_inst200.curr_state_RNI_0_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__33806),
            .in2(_gnd_net_),
            .in3(N__33830),
            .lcout(\b2v_inst200.N_202 ),
            .ltout(\b2v_inst200.N_202_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.HDA_SDO_FPGA_RNIJCSM_LC_12_12_1 .C_ON=1'b0;
    defparam \b2v_inst200.HDA_SDO_FPGA_RNIJCSM_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.HDA_SDO_FPGA_RNIJCSM_LC_12_12_1 .LUT_INIT=16'b1110111001001110;
    LogicCell40 \b2v_inst200.HDA_SDO_FPGA_RNIJCSM_LC_12_12_1  (
            .in0(N__34072),
            .in1(N__33838),
            .in2(N__33508),
            .in3(N__33850),
            .lcout(HDA_SDO_FPGA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_7_c_RNO_LC_12_12_2 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_7_c_RNO_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_7_c_RNO_LC_12_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_7_c_RNO_LC_12_12_2  (
            .in0(N__33483),
            .in1(N__33471),
            .in2(N__33460),
            .in3(N__33444),
            .lcout(\b2v_inst20.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_LC_12_12_3 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_LC_12_12_3 .LUT_INIT=16'b1100110011111101;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m11_0_LC_12_12_3  (
            .in0(N__33770),
            .in1(N__34145),
            .in2(N__34123),
            .in3(N__33849),
            .lcout(G_2788),
            .ltout(G_2788_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNI52VB_2_LC_12_12_4 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNI52VB_2_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNI52VB_2_LC_12_12_4 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \b2v_inst200.curr_state_RNI52VB_2_LC_12_12_4  (
            .in0(N__34105),
            .in1(_gnd_net_),
            .in2(N__34096),
            .in3(N__34071),
            .lcout(\b2v_inst200.curr_stateZ0Z_2 ),
            .ltout(\b2v_inst200.curr_stateZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.HDA_SDO_FPGA_LC_12_12_5 .C_ON=1'b0;
    defparam \b2v_inst200.HDA_SDO_FPGA_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.HDA_SDO_FPGA_LC_12_12_5 .LUT_INIT=16'b1111100011111000;
    LogicCell40 \b2v_inst200.HDA_SDO_FPGA_LC_12_12_5  (
            .in0(N__33831),
            .in1(N__33808),
            .in2(N__33841),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.HDA_SDO_FPGA_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34673),
            .ce(N__33681),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_0_LC_12_12_7 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_0_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.curr_state_0_LC_12_12_7 .LUT_INIT=16'b1111111100001001;
    LogicCell40 \b2v_inst200.curr_state_0_LC_12_12_7  (
            .in0(N__33832),
            .in1(N__33807),
            .in2(N__33777),
            .in3(N__33730),
            .lcout(\b2v_inst200.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34673),
            .ce(N__33681),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_6_LC_12_13_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_6_LC_12_13_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_6_LC_12_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.count_6_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34264),
            .lcout(\b2v_inst6.count_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34680),
            .ce(N__34417),
            .sr(N__35295));
    defparam \b2v_inst6.count_RNIRDTD4_2_LC_12_13_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIRDTD4_2_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIRDTD4_2_LC_12_13_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNIRDTD4_2_LC_12_13_1  (
            .in0(N__34276),
            .in1(N__34284),
            .in2(_gnd_net_),
            .in3(N__34415),
            .lcout(\b2v_inst6.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIVVMK_1_LC_12_13_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIVVMK_1_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIVVMK_1_LC_12_13_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \b2v_inst6.count_RNIVVMK_1_LC_12_13_2  (
            .in0(N__34216),
            .in1(N__35020),
            .in2(_gnd_net_),
            .in3(N__35271),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI3A4A4_1_LC_12_13_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI3A4A4_1_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI3A4A4_1_LC_12_13_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNI3A4A4_1_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__34291),
            .in2(N__33625),
            .in3(N__34414),
            .lcout(\b2v_inst6.countZ0Z_1 ),
            .ltout(\b2v_inst6.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_1_LC_12_13_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_1_LC_12_13_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_1_LC_12_13_4 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \b2v_inst6.count_1_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__35021),
            .in2(N__34294),
            .in3(N__35272),
            .lcout(\b2v_inst6.count_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34680),
            .ce(N__34417),
            .sr(N__35295));
    defparam \b2v_inst6.count_2_LC_12_13_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_2_LC_12_13_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_2_LC_12_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.count_2_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34285),
            .lcout(\b2v_inst6.count_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34680),
            .ce(N__34417),
            .sr(N__35295));
    defparam \b2v_inst6.count_RNI3Q1E4_6_LC_12_13_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI3Q1E4_6_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI3Q1E4_6_LC_12_13_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst6.count_RNI3Q1E4_6_LC_12_13_6  (
            .in0(N__34416),
            .in1(N__34270),
            .in2(_gnd_net_),
            .in3(N__34263),
            .lcout(\b2v_inst6.countZ0Z_6 ),
            .ltout(\b2v_inst6.countZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI_1_LC_12_13_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_1_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_1_LC_12_13_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst6.count_RNI_1_LC_12_13_7  (
            .in0(N__34249),
            .in1(N__34231),
            .in2(N__34219),
            .in3(N__34215),
            .lcout(\b2v_inst6.un12_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI_15_LC_12_14_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_15_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_15_LC_12_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst6.count_RNI_15_LC_12_14_0  (
            .in0(N__34174),
            .in1(N__34201),
            .in2(N__34804),
            .in3(N__34849),
            .lcout(\b2v_inst6.un12_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNITOVM4_12_LC_12_14_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNITOVM4_12_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNITOVM4_12_LC_12_14_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNITOVM4_12_LC_12_14_1  (
            .in0(N__34180),
            .in1(N__34188),
            .in2(_gnd_net_),
            .in3(N__34425),
            .lcout(\b2v_inst6.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_12_LC_12_14_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_12_LC_12_14_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_12_LC_12_14_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst6.count_12_LC_12_14_2  (
            .in0(N__34189),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.count_3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34685),
            .ce(N__34435),
            .sr(N__35308));
    defparam \b2v_inst6.count_RNIVR0N4_13_LC_12_14_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIVR0N4_13_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIVR0N4_13_LC_12_14_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst6.count_RNIVR0N4_13_LC_12_14_3  (
            .in0(N__34153),
            .in1(N__34426),
            .in2(_gnd_net_),
            .in3(N__34161),
            .lcout(\b2v_inst6.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_13_LC_12_14_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_13_LC_12_14_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_13_LC_12_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst6.count_13_LC_12_14_4  (
            .in0(N__34162),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.count_3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34685),
            .ce(N__34435),
            .sr(N__35308));
    defparam \b2v_inst6.count_RNI1V1N4_14_LC_12_14_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI1V1N4_14_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI1V1N4_14_LC_12_14_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNI1V1N4_14_LC_12_14_5  (
            .in0(N__34828),
            .in1(N__34836),
            .in2(_gnd_net_),
            .in3(N__34427),
            .lcout(\b2v_inst6.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_14_LC_12_14_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_14_LC_12_14_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_14_LC_12_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst6.count_14_LC_12_14_6  (
            .in0(N__34837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.count_3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34685),
            .ce(N__34435),
            .sr(N__35308));
    defparam \b2v_inst6.count_RNI323N4_15_LC_12_14_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI323N4_15_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI323N4_15_LC_12_14_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNI323N4_15_LC_12_14_7  (
            .in0(N__34822),
            .in1(N__34815),
            .in2(_gnd_net_),
            .in3(N__34428),
            .lcout(\b2v_inst6.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un8_rsmrst_pwrgd_4_LC_12_15_0 .C_ON=1'b0;
    defparam \b2v_inst5.un8_rsmrst_pwrgd_4_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un8_rsmrst_pwrgd_4_LC_12_15_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst5.un8_rsmrst_pwrgd_4_LC_12_15_0  (
            .in0(N__34789),
            .in1(N__34783),
            .in2(N__34777),
            .in3(N__34768),
            .lcout(SYNTHESIZED_WIRE_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIVVMK_0_LC_12_15_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIVVMK_0_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIVVMK_0_LC_12_15_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst6.count_RNIVVMK_0_LC_12_15_4  (
            .in0(N__35025),
            .in1(N__34915),
            .in2(_gnd_net_),
            .in3(N__35222),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI294A4_0_LC_12_15_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI294A4_0_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI294A4_0_LC_12_15_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNI294A4_0_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(N__34723),
            .in2(N__34729),
            .in3(N__34368),
            .lcout(\b2v_inst6.countZ0Z_0 ),
            .ltout(\b2v_inst6.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_0_LC_12_15_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_0_LC_12_15_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_0_LC_12_15_6 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \b2v_inst6.count_0_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__34914),
            .in2(N__34726),
            .in3(N__35224),
            .lcout(\b2v_inst6.count_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34688),
            .ce(N__34421),
            .sr(N__35228));
    defparam \b2v_inst6.count_3_LC_12_15_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_3_LC_12_15_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_3_LC_12_15_7 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst6.count_3_LC_12_15_7  (
            .in0(N__35223),
            .in1(N__34916),
            .in2(N__35094),
            .in3(N__34717),
            .lcout(\b2v_inst6.count_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34688),
            .ce(N__34421),
            .sr(N__35228));
    defparam \b2v_inst6.count_RNI_3_LC_12_16_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_3_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_3_LC_12_16_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst6.count_RNI_3_LC_12_16_5  (
            .in0(N__35125),
            .in1(N__35092),
            .in2(N__35062),
            .in3(N__35016),
            .lcout(),
            .ltout(\b2v_inst6.un12_clk_100khz_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI_0_1_LC_12_16_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_0_1_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_0_1_LC_12_16_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst6.count_RNI_0_1_LC_12_16_6  (
            .in0(N__34987),
            .in1(N__34981),
            .in2(N__34972),
            .in3(N__34969),
            .lcout(\b2v_inst6.N_1_i ),
            .ltout(\b2v_inst6.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI_1_1_LC_12_16_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_1_1_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_1_1_LC_12_16_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst6.count_RNI_1_1_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34945),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.N_1_i_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TOP
