-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Aug 28 2022 11:53:56

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : in std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : out std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : out std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : out std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__21309\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \VCCG0\ : std_logic;
signal \PCH_PWRGD.un4_count_11\ : std_logic;
signal \PCH_PWRGD.un4_count_9\ : std_logic;
signal \PCH_PWRGD.un4_count_10_cascade_\ : std_logic;
signal \PCH_PWRGD.N_1_i_cascade_\ : std_logic;
signal \PCH_PWRGD.un1_curr_state_0_sqmuxa_0_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_RNI7N705Z0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.un4_count_8\ : std_logic;
signal \PCH_PWRGD.N_3_i_cascade_\ : std_logic;
signal vr_ready_vccin : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \PCH_PWRGD.N_1_i\ : std_logic;
signal \PCH_PWRGD.N_3_i\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \bfn_1_5_0_\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8_cascade_\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un96_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8_cascade_\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un103_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8_cascade_\ : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un110_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un110_sum_s_8_cascade_\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un124_sum_s_8_cascade_\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un131_sum_s_8_cascade_\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un138_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8_cascade_\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7_cascade_\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_0\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5_s\ : std_logic;
signal \G_407\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un166_sum_axb_6\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum_i\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8\ : std_logic;
signal pwrbtn_led : std_logic;
signal \PCH_PWRGD.un1_curr_state10_0\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0\ : std_logic;
signal \bfn_2_2_0_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_1\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \PCH_PWRGD.countZ0Z_2\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \PCH_PWRGD.countZ0Z_3\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \PCH_PWRGD.countZ0Z_5\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \PCH_PWRGD.countZ0Z_7\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \PCH_PWRGD.countZ0Z_8\ : std_logic;
signal \bfn_2_3_0_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \PCH_PWRGD.countZ0Z_10\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \PCH_PWRGD.countZ0Z_11\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \PCH_PWRGD.countZ0Z_12\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \PCH_PWRGD.countZ0Z_13\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \PCH_PWRGD.countZ0Z_14\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_2_4_0_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15\ : std_logic;
signal \PCH_PWRGD.N_65_3\ : std_logic;
signal \PCH_PWRGD.curr_state_RNI7N705Z0Z_0\ : std_logic;
signal \bfn_2_5_0_\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un89_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un82_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_0_8\ : std_logic;
signal \bfn_2_6_0_\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un82_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_0_8\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un75_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_i\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_i\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un110_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un117_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un117_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_i\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_4_l_fx\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8_cascade_\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \POWERLED.mult1_un145_sum_i\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un159_sum_axb_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un152_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un152_sum_i_0_8\ : std_logic;
signal \POWERLED.un1_count_2_0\ : std_logic;
signal \POWERLED.count_i_0_0\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \POWERLED.un1_count_2_1\ : std_logic;
signal \POWERLED.count_i_1\ : std_logic;
signal \POWERLED.un1_count_2_cry_0\ : std_logic;
signal \POWERLED.un1_count_2_2\ : std_logic;
signal \POWERLED.count_i_2\ : std_logic;
signal \POWERLED.un1_count_2_cry_1\ : std_logic;
signal \POWERLED.un1_count_2_3\ : std_logic;
signal \POWERLED.count_i_3\ : std_logic;
signal \POWERLED.un1_count_2_cry_2\ : std_logic;
signal \POWERLED.count_i_4\ : std_logic;
signal \POWERLED.un1_count_2_cry_3\ : std_logic;
signal \POWERLED.un1_count_2_5\ : std_logic;
signal \POWERLED.count_i_5\ : std_logic;
signal \POWERLED.un1_count_2_cry_4\ : std_logic;
signal \POWERLED.un1_count_2_6\ : std_logic;
signal \POWERLED.count_i_6\ : std_logic;
signal \POWERLED.un1_count_2_cry_5\ : std_logic;
signal \POWERLED.un1_count_2_7\ : std_logic;
signal \POWERLED.count_i_7\ : std_logic;
signal \POWERLED.un1_count_2_cry_6\ : std_logic;
signal \POWERLED.un1_count_2_cry_7\ : std_logic;
signal \POWERLED.un1_count_2_8\ : std_logic;
signal \POWERLED.count_i_8\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \POWERLED.un1_count_2_9\ : std_logic;
signal \POWERLED.count_i_9\ : std_logic;
signal \POWERLED.un1_count_2_cry_8\ : std_logic;
signal \POWERLED.un1_count_2_10\ : std_logic;
signal \POWERLED.count_i_10\ : std_logic;
signal \POWERLED.un1_count_2_cry_9\ : std_logic;
signal \POWERLED.un1_count_2_11\ : std_logic;
signal \POWERLED.count_i_11\ : std_logic;
signal \POWERLED.un1_count_2_cry_10\ : std_logic;
signal \POWERLED.un1_count_2_12\ : std_logic;
signal \POWERLED.count_i_12\ : std_logic;
signal \POWERLED.un1_count_2_cry_11\ : std_logic;
signal \POWERLED.un1_count_2_13\ : std_logic;
signal \POWERLED.count_i_13\ : std_logic;
signal \POWERLED.un1_count_2_cry_12\ : std_logic;
signal \POWERLED.un1_count_2_14\ : std_logic;
signal \POWERLED.count_i_14\ : std_logic;
signal \POWERLED.un1_count_2_cry_13\ : std_logic;
signal \POWERLED.un1_count_2_15\ : std_logic;
signal \POWERLED.count_i_15\ : std_logic;
signal \POWERLED.un1_count_2_cry_14\ : std_logic;
signal \POWERLED.un1_count_2_cry_15\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \POWERLED.un1_count_2_cry_15_THRU_CO\ : std_logic;
signal \POWERLED.un1_count_2_cry_15_THRU_CO_cascade_\ : std_logic;
signal \POWERLED.pwm_out_RNOZ0\ : std_logic;
signal vpp_ok : std_logic;
signal vddq_en : std_logic;
signal gpio_fpga_soc_1 : std_logic;
signal \HDA_STRAP.N_5_0_cascade_\ : std_logic;
signal pch_pwrok : std_logic;
signal \HDA_STRAP.m14_ns_1\ : std_logic;
signal \bfn_4_5_0_\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7\ : std_logic;
signal \bfn_4_6_0_\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7_THRU_CO\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un68_sum_i\ : std_logic;
signal \bfn_4_7_0_\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6_THRU_CO\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_i\ : std_logic;
signal \POWERLED.mult1_un138_sum_i\ : std_logic;
signal \POWERLED.mult1_un124_sum_i\ : std_logic;
signal \POWERLED.mult1_un117_sum_i\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_7_l_fx\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8\ : std_logic;
signal \POWERLED.un1_count_2_4\ : std_logic;
signal v5s_enn : std_logic;
signal \POWERLED.mult1_un159_sum_i\ : std_logic;
signal \POWERLED.mult1_un152_sum_i\ : std_logic;
signal \POWERLED.un1_countlt6_0_cascade_\ : std_logic;
signal \POWERLED.g0_0_7_cascade_\ : std_logic;
signal \POWERLED.un1_count_0\ : std_logic;
signal \POWERLED.un1_countlto15_5_cascade_\ : std_logic;
signal \POWERLED.g0_0_4\ : std_logic;
signal \POWERLED.un1_countlt6\ : std_logic;
signal \POWERLED.g0_0_5\ : std_logic;
signal \POWERLED.un1_countlto15_4_cascade_\ : std_logic;
signal \POWERLED.un1_countlto15_7\ : std_logic;
signal \POWERLED.count_RNIOVT24Z0Z_11\ : std_logic;
signal \POWERLED.curr_stateZ0Z_0\ : std_logic;
signal \POWERLED.count_RNIOVT24Z0Z_11_cascade_\ : std_logic;
signal \HDA_STRAP.N_5_0\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_2\ : std_logic;
signal hda_sdo_atp : std_logic;
signal \POWERLED.mult1_un82_sum_i\ : std_logic;
signal \POWERLED.un1_dutycycle_1_i_28\ : std_logic;
signal \POWERLED.un1_dutycycle_1_19_0_cascade_\ : std_logic;
signal \POWERLED.mult1_un75_sum_i\ : std_logic;
signal \POWERLED.N_53\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_4\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_5\ : std_logic;
signal \POWERLED.mult1_un47_sum_axb_4\ : std_logic;
signal \POWERLED.un1_dutycycle_1_i_29\ : std_logic;
signal \POWERLED.mult1_un61_sum_i\ : std_logic;
signal \POWERLED.mult1_un54_sum_i\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_0\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_1\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_2\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_3\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_4\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_5\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_6\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_7\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_8\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_9\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_10\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_11\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_12\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_13\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_14\ : std_logic;
signal \POWERLED.count_offZ0Z_12\ : std_logic;
signal \POWERLED.count_offZ0Z_13\ : std_logic;
signal \POWERLED.count_offZ0Z_15\ : std_logic;
signal \POWERLED.count_offZ0Z_1\ : std_logic;
signal \POWERLED.count_offZ0Z_11\ : std_logic;
signal \POWERLED.count_offZ0Z_0\ : std_logic;
signal \POWERLED.count_offZ0Z_14\ : std_logic;
signal \POWERLED.count_offZ0Z_10\ : std_logic;
signal \POWERLED.count_offZ0Z_8\ : std_logic;
signal \POWERLED.count_offZ0Z_6\ : std_logic;
signal \POWERLED.count_offZ0Z_9\ : std_logic;
signal \POWERLED.count_offZ0Z_5\ : std_logic;
signal \POWERLED.func_state_ns_0_a2_11_0\ : std_logic;
signal \POWERLED.func_state_ns_0_a2_10_0\ : std_logic;
signal \POWERLED.func_state_ns_0_a2_9_0_cascade_\ : std_logic;
signal \POWERLED.count_off_0_sqmuxa\ : std_logic;
signal \POWERLED.count_off_0_sqmuxa_cascade_\ : std_logic;
signal \POWERLED.N_85_1\ : std_logic;
signal \POWERLED.countZ0Z_0\ : std_logic;
signal \POWERLED.countZ0Z_1\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \POWERLED.countZ0Z_2\ : std_logic;
signal \POWERLED.un1_count_1_cry_1\ : std_logic;
signal \POWERLED.countZ0Z_3\ : std_logic;
signal \POWERLED.un1_count_1_cry_2\ : std_logic;
signal \POWERLED.countZ0Z_4\ : std_logic;
signal \POWERLED.un1_count_1_cry_3\ : std_logic;
signal \POWERLED.countZ0Z_5\ : std_logic;
signal \POWERLED.un1_count_1_cry_4\ : std_logic;
signal \POWERLED.countZ0Z_6\ : std_logic;
signal \POWERLED.un1_count_1_cry_5\ : std_logic;
signal \POWERLED.countZ0Z_7\ : std_logic;
signal \POWERLED.un1_count_1_cry_6\ : std_logic;
signal \POWERLED.countZ0Z_8\ : std_logic;
signal \POWERLED.un1_count_1_cry_7\ : std_logic;
signal \POWERLED.un1_count_1_cry_8\ : std_logic;
signal \POWERLED.countZ0Z_9\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \POWERLED.countZ0Z_10\ : std_logic;
signal \POWERLED.un1_count_1_cry_9\ : std_logic;
signal \POWERLED.countZ0Z_11\ : std_logic;
signal \POWERLED.un1_count_1_cry_10\ : std_logic;
signal \POWERLED.countZ0Z_12\ : std_logic;
signal \POWERLED.un1_count_1_cry_11\ : std_logic;
signal \POWERLED.countZ0Z_13\ : std_logic;
signal \POWERLED.un1_count_1_cry_12\ : std_logic;
signal \POWERLED.countZ0Z_14\ : std_logic;
signal \POWERLED.un1_count_1_cry_13\ : std_logic;
signal \POWERLED.un1_count_1_cry_14\ : std_logic;
signal \POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO\ : std_logic;
signal \bfn_5_16_0_\ : std_logic;
signal \POWERLED.countZ0Z_15\ : std_logic;
signal \POWERLED.N_65_5\ : std_logic;
signal \POWERLED.curr_state_RNI75RB5Z0Z_0\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_0\ : std_logic;
signal \bfn_6_1_0_\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_0\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_1\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_2\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_3\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_4\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_5\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_6\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_7\ : std_logic;
signal \bfn_6_2_0_\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_8\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_9\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_11\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_10\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_11\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_12\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_13\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_14\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_15\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_16\ : std_logic;
signal \POWERLED.un1_dutycycle_1_axb_0\ : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_1_axb_1\ : std_logic;
signal \POWERLED.mult1_un138_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_0\ : std_logic;
signal \POWERLED.dutycycle_RNI16B71Z0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNIFHLJZ0Z_0\ : std_logic;
signal \POWERLED.mult1_un131_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_1\ : std_logic;
signal \POWERLED.mult1_un124_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_3\ : std_logic;
signal \POWERLED.dutycycle_RNIEJ021Z0Z_4\ : std_logic;
signal \POWERLED.mult1_un110_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_4\ : std_logic;
signal \POWERLED.dutycycle_RNI6NI81Z0Z_5\ : std_logic;
signal \POWERLED.mult1_un103_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_5\ : std_logic;
signal \POWERLED.dutycycle_RNIJNBA1Z0Z_6\ : std_logic;
signal \POWERLED.mult1_un96_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_6\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_7\ : std_logic;
signal \POWERLED.mult1_un89_sum\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \POWERLED.mult1_un82_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_8\ : std_logic;
signal \POWERLED.mult1_un75_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_9\ : std_logic;
signal \POWERLED.mult1_un68_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_10\ : std_logic;
signal \POWERLED.mult1_un61_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_11\ : std_logic;
signal \POWERLED.mult1_un54_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_12\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_15\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71\ : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal \POWERLED.CO2\ : std_logic;
signal \POWERLED.CO2_THRU_CO\ : std_logic;
signal \POWERLED.dutycycle_fastZ0Z_5\ : std_logic;
signal \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNIE4FLZ0Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNI53MGZ0Z_14\ : std_logic;
signal \POWERLED.dutycycle_RNI84C11Z0Z_14\ : std_logic;
signal \POWERLED.dutycycle_RNIB1FLZ0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNI75MGZ0Z_15\ : std_logic;
signal \POWERLED.un1_dutycycle_1_34_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_1_axb_8_cascade_\ : std_logic;
signal \POWERLED.dutycycle_fast_RNILMLMZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNIJL1R1Z0Z_6\ : std_logic;
signal \POWERLED.dutycycle_fastZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNI2V0PZ0Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNI2V0PZ0Z_10_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI712I1Z0Z_15\ : std_logic;
signal \POWERLED.dutycycle_RNIQ09G1Z0Z_10\ : std_logic;
signal \POWERLED.count_offZ0Z_3\ : std_logic;
signal \POWERLED.count_offZ0Z_7\ : std_logic;
signal \POWERLED.count_offZ0Z_4\ : std_logic;
signal \POWERLED.count_offZ0Z_2\ : std_logic;
signal \POWERLED.func_state_ns_0_a2_8_0\ : std_logic;
signal \POWERLED.un1_dutycycle_1_44_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIF3561Z0Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNIC8C11Z0Z_15\ : std_logic;
signal \POWERLED.dutycycle_RNI73C11Z0Z_15\ : std_logic;
signal \POWERLED.N_368_0_i_i_a6_0\ : std_logic;
signal \POWERLED.N_207_cascade_\ : std_logic;
signal \POWERLED.N_48\ : std_logic;
signal \POWERLED.N_149\ : std_logic;
signal \POWERLED.N_149_cascade_\ : std_logic;
signal \POWERLED.N_214\ : std_logic;
signal \POWERLED.N_213\ : std_logic;
signal \POWERLED.N_234\ : std_logic;
signal \POWERLED.N_218_cascade_\ : std_logic;
signal \POWERLED.N_248\ : std_logic;
signal \POWERLED.N_88_cascade_\ : std_logic;
signal \POWERLED.N_208_cascade_\ : std_logic;
signal \POWERLED.func_state_ns_i_0_1_1\ : std_logic;
signal \POWERLED.N_222\ : std_logic;
signal \POWERLED.N_222_cascade_\ : std_logic;
signal \POWERLED.N_228\ : std_logic;
signal \POWERLED.N_211_cascade_\ : std_logic;
signal \POWERLED.func_state_ns_i_0_0_1\ : std_logic;
signal \POWERLED.N_179\ : std_logic;
signal \POWERLED.N_178\ : std_logic;
signal \POWERLED.N_180\ : std_logic;
signal \POWERLED.N_250\ : std_logic;
signal \HDA_STRAP.curr_state_RNIH91AZ0Z_0\ : std_logic;
signal \HDA_STRAP.countZ0Z_2\ : std_logic;
signal \HDA_STRAP.countZ0Z_1\ : std_logic;
signal \HDA_STRAP.countZ0Z_3\ : std_logic;
signal \HDA_STRAP.countZ0Z_0\ : std_logic;
signal \HDA_STRAP.countZ0Z_14\ : std_logic;
signal \HDA_STRAP.countZ0Z_15\ : std_logic;
signal \HDA_STRAP.countZ0Z_12\ : std_logic;
signal \HDA_STRAP.un4_count_9_cascade_\ : std_logic;
signal \HDA_STRAP.countZ0Z_13\ : std_logic;
signal \HDA_STRAP.countZ0Z_7\ : std_logic;
signal \HDA_STRAP.countZ0Z_5\ : std_logic;
signal \HDA_STRAP.countZ0Z_9\ : std_logic;
signal \HDA_STRAP.countZ0Z_4\ : std_logic;
signal \HDA_STRAP.countZ0Z_11\ : std_logic;
signal \HDA_STRAP.un4_count_12\ : std_logic;
signal \HDA_STRAP.un4_count_11\ : std_logic;
signal \HDA_STRAP.un4_count_10_cascade_\ : std_logic;
signal \HDA_STRAP.un4_count_13\ : std_logic;
signal \HDA_STRAP.count_RNIB5IA5Z0Z_0_cascade_\ : std_logic;
signal \HDA_STRAP.curr_state_RNO_0Z0Z_2\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_10\ : std_logic;
signal \HDA_STRAP.countZ0Z_10\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_16\ : std_logic;
signal \HDA_STRAP.countZ0Z_16\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_17\ : std_logic;
signal \HDA_STRAP.countZ0Z_17\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_8\ : std_logic;
signal \HDA_STRAP.countZ0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNI31MG_0Z0Z_12\ : std_logic;
signal \POWERLED.dutycycle_RNI31MGZ0Z_12\ : std_logic;
signal \POWERLED.un1_dutycycle_1_39_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI34C41Z0Z_8\ : std_logic;
signal \POWERLED.N_117\ : std_logic;
signal \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNIK4I81Z0Z_6\ : std_logic;
signal \POWERLED.dutycycle_lm_0_1_2\ : std_logic;
signal \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNIQAI81Z0Z_4\ : std_logic;
signal \POWERLED.dutycycle_RNIOQLJZ0Z_4\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_0\ : std_logic;
signal \POWERLED.dutycycle_s_0\ : std_logic;
signal \POWERLED.dutycycle_cry_c_0_THRU_CO\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1\ : std_logic;
signal \POWERLED.dutycycle_s_1\ : std_logic;
signal \POWERLED.dutycycle_cry_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2\ : std_logic;
signal \POWERLED.dutycycle_s_2\ : std_logic;
signal \POWERLED.dutycycle_cry_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_3\ : std_logic;
signal \POWERLED.dutycycle_cry_2\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4\ : std_logic;
signal \POWERLED.dutycycle_cry_3\ : std_logic;
signal \POWERLED.dutycycleZ0Z_5\ : std_logic;
signal \POWERLED.dutycycle_s_5\ : std_logic;
signal \POWERLED.dutycycle_cry_4\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_s_6\ : std_logic;
signal \POWERLED.dutycycle_cry_5\ : std_logic;
signal \POWERLED.dutycycle_cry_6\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7\ : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal \POWERLED.dutycycle_cry_7\ : std_logic;
signal \POWERLED.dutycycle_cry_8\ : std_logic;
signal \POWERLED.dutycycle_cry_9\ : std_logic;
signal \POWERLED.dutycycle_cry_10\ : std_logic;
signal \POWERLED.dutycycle_cry_11\ : std_logic;
signal \POWERLED.dutycycle_cry_12\ : std_logic;
signal \POWERLED.dutycycle_cry_13\ : std_logic;
signal \POWERLED.dutycycle_cry_14\ : std_logic;
signal \POWERLED.N_177\ : std_logic;
signal \bfn_7_9_0_\ : std_logic;
signal \POWERLED.N_246_cascade_\ : std_logic;
signal \POWERLED.N_203_4\ : std_logic;
signal \POWERLED.N_203_4_cascade_\ : std_logic;
signal \POWERLED.N_203_cascade_\ : std_logic;
signal \POWERLED.N_251_cascade_\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_1_0\ : std_logic;
signal \POWERLED.count_clk_139_tz_0\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_cascade_\ : std_logic;
signal \POWERLED.N_246\ : std_logic;
signal \POWERLED.N_205\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_a6_3_0_cascade_\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_1\ : std_logic;
signal \POWERLED.N_127\ : std_logic;
signal \POWERLED.count_clk_1_sqmuxa_5_0_1\ : std_logic;
signal \POWERLED.N_127_cascade_\ : std_logic;
signal \POWERLED.count_clk_1_sqmuxa_5_0_0\ : std_logic;
signal \POWERLED.N_88\ : std_logic;
signal \POWERLED.dutycycle_3_sqmuxa_1_i_0_1_1_cascade_\ : std_logic;
signal \POWERLED.N_200_2\ : std_logic;
signal \POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_1\ : std_logic;
signal \POWERLED.N_366_1_cascade_\ : std_logic;
signal \POWERLED.N_251\ : std_logic;
signal \POWERLED.dutycycle\ : std_logic;
signal \POWERLED.N_243\ : std_logic;
signal slp_s4n : std_logic;
signal \POWERLED.func_stateZ0Z_1\ : std_logic;
signal \POWERLED.func_stateZ0Z_0\ : std_logic;
signal \POWERLED.count_off_RNIIKVR3Z0Z_10\ : std_logic;
signal \POWERLED.N_148\ : std_logic;
signal slp_s3n : std_logic;
signal vccst_en : std_logic;
signal vpp_en : std_logic;
signal \N_55\ : std_logic;
signal \VPP_VDDQ.N_238\ : std_logic;
signal \VPP_VDDQ.N_238_cascade_\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\ : std_logic;
signal \VPP_VDDQ.G_127_0\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgdZ0\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_1\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_0\ : std_logic;
signal \VPP_VDDQ.N_128\ : std_logic;
signal \VPP_VDDQ.N_154_cascade_\ : std_logic;
signal \HDA_STRAP.count_RNO_0Z0Z_6\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_1\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_0\ : std_logic;
signal \HDA_STRAP.count_RNIB5IA5Z0Z_0\ : std_logic;
signal \HDA_STRAP.countZ0Z_6\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \POWERLED.dutycycle_RNIO18NZ0Z_9\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13\ : std_logic;
signal \POWERLED.dutycycleZ0Z_12\ : std_logic;
signal \POWERLED.dutycycleZ0Z_14\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11\ : std_logic;
signal \POWERLED.dutycycleZ0Z_15\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_o2_3_7\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_o2_3_8_cascade_\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_o2_3_6\ : std_logic;
signal \POWERLED.N_112\ : std_logic;
signal \POWERLED.N_366_1\ : std_logic;
signal \POWERLED.un1_dutycycle_4_sqmuxa_0\ : std_logic;
signal \POWERLED.N_177_5\ : std_logic;
signal \POWERLED.count_clk_0_sqmuxa_5_0_o2_0_0_cascade_\ : std_logic;
signal \POWERLED.N_141\ : std_logic;
signal \POWERLED.N_136_cascade_\ : std_logic;
signal \POWERLED.N_146\ : std_logic;
signal \POWERLED.count_clk_0_sqmuxa_5_0_a6_1\ : std_logic;
signal \POWERLED.count_clk_0_sqmuxa_5_0_o2_4\ : std_logic;
signal gpio_fpga_soc_4 : std_logic;
signal \POWERLED.count_off_1_sqmuxa_i_a6_0_1_cascade_\ : std_logic;
signal \POWERLED.N_136\ : std_logic;
signal \POWERLED.count_off_1_sqmuxa_i_a6_0_3\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \VPP_VDDQ.N_108_i\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_0\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_1\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_2\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_3\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_4\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_5\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_7\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_8\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_9\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_10\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_11\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_12\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_13\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \VPP_VDDQ.N_65_1\ : std_logic;
signal \VPP_VDDQ.curr_state_RNIGR9S7Z0Z_0\ : std_logic;
signal \COUNTER.counterZ0Z_1\ : std_logic;
signal \bfn_9_1_0_\ : std_logic;
signal \COUNTER.counter_1_cry_1\ : std_logic;
signal \COUNTER.counter_1_cry_2\ : std_logic;
signal \COUNTER.counter_1_cry_3\ : std_logic;
signal \COUNTER.counterZ0Z_5\ : std_logic;
signal \COUNTER.counter_1_cry_4_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_4\ : std_logic;
signal \COUNTER.counterZ0Z_6\ : std_logic;
signal \COUNTER.counter_1_cry_5_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_5\ : std_logic;
signal \COUNTER.counterZ0Z_7\ : std_logic;
signal \COUNTER.counter_1_cry_6\ : std_logic;
signal \COUNTER.counter_1_cry_7\ : std_logic;
signal \COUNTER.counter_1_cry_8\ : std_logic;
signal \bfn_9_2_0_\ : std_logic;
signal \COUNTER.counter_1_cry_9\ : std_logic;
signal \COUNTER.counter_1_cry_10\ : std_logic;
signal \COUNTER.counter_1_cry_11\ : std_logic;
signal \COUNTER.counter_1_cry_12\ : std_logic;
signal \COUNTER.counter_1_cry_13\ : std_logic;
signal \COUNTER.counter_1_cry_14\ : std_logic;
signal \COUNTER.counter_1_cry_15\ : std_logic;
signal \COUNTER.counter_1_cry_16\ : std_logic;
signal \bfn_9_3_0_\ : std_logic;
signal \COUNTER.counter_1_cry_17\ : std_logic;
signal \COUNTER.counter_1_cry_18\ : std_logic;
signal \COUNTER.counter_1_cry_19\ : std_logic;
signal \COUNTER.counter_1_cry_20\ : std_logic;
signal \COUNTER.counter_1_cry_21\ : std_logic;
signal \COUNTER.counter_1_cry_22\ : std_logic;
signal \COUNTER.counter_1_cry_23\ : std_logic;
signal \COUNTER.counter_1_cry_24\ : std_logic;
signal \bfn_9_4_0_\ : std_logic;
signal \COUNTER.counter_1_cry_25\ : std_logic;
signal \COUNTER.counter_1_cry_26\ : std_logic;
signal \COUNTER.counter_1_cry_27\ : std_logic;
signal \COUNTER.counter_1_cry_28\ : std_logic;
signal \COUNTER.counter_1_cry_29\ : std_logic;
signal \COUNTER.counter_1_cry_30\ : std_logic;
signal \COUNTER.counterZ0Z_22\ : std_logic;
signal \COUNTER.counterZ0Z_21\ : std_logic;
signal \COUNTER.counterZ0Z_23\ : std_logic;
signal \COUNTER.counterZ0Z_20\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_5\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_3\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_11\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_2\ : std_logic;
signal \COUNTER.counterZ0Z_26\ : std_logic;
signal \COUNTER.counterZ0Z_25\ : std_logic;
signal \COUNTER.counterZ0Z_27\ : std_logic;
signal \COUNTER.counterZ0Z_24\ : std_logic;
signal \COUNTER.counterZ0Z_30\ : std_logic;
signal \COUNTER.counterZ0Z_28\ : std_logic;
signal \COUNTER.counterZ0Z_29\ : std_logic;
signal \COUNTER.counterZ0Z_31\ : std_logic;
signal \COUNTER.counter_1_cry_3_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_4\ : std_logic;
signal \COUNTER.counterZ0Z_0\ : std_logic;
signal \COUNTER.counter_1_cry_1_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_2\ : std_logic;
signal \COUNTER.counter_1_cry_2_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_3\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_7\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_8\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_6\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_4\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_14\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_15\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_13\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_12\ : std_logic;
signal \ALL_SYS_PWRGD.un4_count_10\ : std_logic;
signal \ALL_SYS_PWRGD.un4_count_11_cascade_\ : std_logic;
signal \ALL_SYS_PWRGD.un4_count_8\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_1\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_9\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_10\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_0\ : std_logic;
signal \ALL_SYS_PWRGD.un4_count_9\ : std_logic;
signal \ALL_SYS_PWRGD.curr_state_RNIKNST6Z0Z_0\ : std_logic;
signal \ALL_SYS_PWRGD.curr_state_RNIKNST6Z0Z_0_cascade_\ : std_logic;
signal \ALL_SYS_PWRGD.N_65_4\ : std_logic;
signal slp_susn : std_logic;
signal v5a_ok : std_logic;
signal v33a_ok : std_logic;
signal v1p8a_ok : std_logic;
signal \COUNTER.tmp_i\ : std_logic;
signal \tmp_RNIRH3P\ : std_logic;
signal \POWERLED.count_clk_1_sqmuxa_5_i\ : std_logic;
signal \POWERLED.count_clkZ0Z_0\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \POWERLED.count_clkZ0Z_1\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_0\ : std_logic;
signal \POWERLED.count_clkZ0Z_2\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_1\ : std_logic;
signal \POWERLED.count_clkZ0Z_3\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_2\ : std_logic;
signal \POWERLED.count_clkZ0Z_4\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_3\ : std_logic;
signal \POWERLED.count_clkZ0Z_5\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_4\ : std_logic;
signal \POWERLED.count_clkZ0Z_6\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_5\ : std_logic;
signal \POWERLED.count_clkZ0Z_7\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_6\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_7\ : std_logic;
signal \POWERLED.count_clkZ0Z_8\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \POWERLED.count_clkZ0Z_9\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_8\ : std_logic;
signal \POWERLED.count_clkZ0Z_10\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_9\ : std_logic;
signal \POWERLED.count_clkZ0Z_11\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_10\ : std_logic;
signal \POWERLED.count_clkZ0Z_12\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_11\ : std_logic;
signal \POWERLED.count_clkZ0Z_13\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_12\ : std_logic;
signal \POWERLED.count_clkZ0Z_14\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_13\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_14\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \POWERLED.count_clkZ0Z_15\ : std_logic;
signal \POWERLED.N_65_0\ : std_logic;
signal \POWERLED.count_clk_RNIOH1J11Z0Z_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_11\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_13\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_6\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_9\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_12\ : std_logic;
signal \RSMRST_PWRGD.m4_i_i_a2_0_11\ : std_logic;
signal \RSMRST_PWRGD.m4_i_i_a2_0_9_cascade_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_15\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_7\ : std_logic;
signal \RSMRST_PWRGD.m4_i_i_a2_0_7_cascade_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_3\ : std_logic;
signal \RSMRST_PWRGD.m4_i_i_a2_0_12\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_4\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_2\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_5\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.m4_i_i_a2_0_10\ : std_logic;
signal \RSMRST_PWRGD.N_240_cascade_\ : std_logic;
signal \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0\ : std_logic;
signal \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_65_2\ : std_logic;
signal \RSMRST_PWRGD.N_37\ : std_logic;
signal \VPP_VDDQ.countZ0Z_5\ : std_logic;
signal \VPP_VDDQ.countZ0Z_4\ : std_logic;
signal \VPP_VDDQ.countZ0Z_7\ : std_logic;
signal \VPP_VDDQ.countZ0Z_3\ : std_logic;
signal \VPP_VDDQ.countZ0Z_14\ : std_logic;
signal \VPP_VDDQ.countZ0Z_15\ : std_logic;
signal \VPP_VDDQ.countZ0Z_13\ : std_logic;
signal \VPP_VDDQ.countZ0Z_12\ : std_logic;
signal \VPP_VDDQ.countZ0Z_6\ : std_logic;
signal \VPP_VDDQ.countZ0Z_2\ : std_logic;
signal \VPP_VDDQ.countZ0Z_10\ : std_logic;
signal \VPP_VDDQ.countZ0Z_1\ : std_logic;
signal \VPP_VDDQ.countZ0Z_9\ : std_logic;
signal \VPP_VDDQ.countZ0Z_8\ : std_logic;
signal \VPP_VDDQ.countZ0Z_11\ : std_logic;
signal \VPP_VDDQ.countZ0Z_0\ : std_logic;
signal \VPP_VDDQ.un6_count_11\ : std_logic;
signal \VPP_VDDQ.un6_count_10\ : std_logic;
signal \VPP_VDDQ.un6_count_9_cascade_\ : std_logic;
signal \VPP_VDDQ.un6_count_8\ : std_logic;
signal \VPP_VDDQ.count_esr_RNIRFM64Z0Z_15\ : std_logic;
signal \COUNTER.counterZ0Z_14\ : std_logic;
signal \COUNTER.counterZ0Z_13\ : std_logic;
signal \COUNTER.counterZ0Z_15\ : std_logic;
signal \COUNTER.counterZ0Z_12\ : std_logic;
signal \COUNTER.counterZ0Z_18\ : std_logic;
signal \COUNTER.counterZ0Z_17\ : std_logic;
signal \COUNTER.counterZ0Z_19\ : std_logic;
signal \COUNTER.counterZ0Z_16\ : std_logic;
signal \COUNTER.counterZ0Z_10\ : std_logic;
signal \COUNTER.counterZ0Z_9\ : std_logic;
signal \COUNTER.counterZ0Z_11\ : std_logic;
signal \COUNTER.counterZ0Z_8\ : std_logic;
signal \COUNTER.un4_counter_0_and\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \COUNTER.un4_counter_1_and\ : std_logic;
signal \COUNTER.un4_counter_0\ : std_logic;
signal \COUNTER.un4_counter_2_and\ : std_logic;
signal \COUNTER.un4_counter_1\ : std_logic;
signal \COUNTER.un4_counter_3_and\ : std_logic;
signal \COUNTER.un4_counter_2\ : std_logic;
signal \COUNTER.un4_counter_4_and\ : std_logic;
signal \COUNTER.un4_counter_3\ : std_logic;
signal \COUNTER.un4_counter_5_and\ : std_logic;
signal \COUNTER.un4_counter_4\ : std_logic;
signal \COUNTER.un4_counter_6_and\ : std_logic;
signal \COUNTER.un4_counter_5\ : std_logic;
signal \COUNTER.un4_counter_7_and\ : std_logic;
signal \COUNTER.un4_counter_6\ : std_logic;
signal \COUNTER.un4_counter_7\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \COUNTER.un4_counter_7_THRU_CO\ : std_logic;
signal \ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa_cascade_\ : std_logic;
signal \ALL_SYS_PWRGD.un1_curr_state10_0\ : std_logic;
signal \ALL_SYS_PWRGD.N_1_i\ : std_logic;
signal \ALL_SYS_PWRGD.N_36\ : std_logic;
signal \ALL_SYS_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \ALL_SYS_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal vccst_pwrgd : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.N_241\ : std_logic;
signal \RSMRST_PWRGD.N_240\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal rsmrstn : std_logic;
signal fpga_osc : std_logic;
signal \N_65_g\ : std_logic;
signal vddq_ok : std_logic;
signal v5s_ok : std_logic;
signal rsmrst_pwrgd_signal : std_logic;
signal vccst_cpu_ok : std_logic;
signal \ALL_SYS_PWRGD.m4_0_0_a2_1_cascade_\ : std_logic;
signal v33s_ok : std_logic;
signal \ALL_SYS_PWRGD.N_245\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \VCCST_OVERRIDE_3V3_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \SLP_S0n_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \PWRBTNn_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \GPIO_FPGA_SoC_2_wire\ : std_logic;
signal \VCCIN_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \CPU_C10_GATE_N_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \TPM_GPIO_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \PLTRSTn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \FPGA_OSC_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \SPI_FP_IO2_wire\ : std_logic;
signal \SATAXPCIE1_FPGA_wire\ : std_logic;
signal \GPIO_FPGA_EXP_1_wire\ : std_logic;
signal \VCCINAUX_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \GPIO_FPGA_EXP_2_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSACK_N_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \GPIO_FPGA_SoC_3_wire\ : std_logic;
signal \VR_PROCHOT_FPGA_OUT_N_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \SOC_SPKR_wire\ : std_logic;
signal \SLP_S5n_wire\ : std_logic;
signal \V12_MAIN_MON_wire\ : std_logic;
signal \SPI_FP_IO3_wire\ : std_logic;
signal \SATAXPCIE0_FPGA_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \FPGA_SLP_WLAN_N_wire\ : std_logic;

begin
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    V33A_ENn <= \V33A_ENn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \VCCST_OVERRIDE_3V3_wire\ <= VCCST_OVERRIDE_3V3;
    \V5S_OK_wire\ <= V5S_OK;
    \SLP_S3n_wire\ <= SLP_S3n;
    \SLP_S0n_wire\ <= SLP_S0n;
    V5S_ENn <= \V5S_ENn_wire\;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \PWRBTNn_wire\ <= PWRBTNn;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \GPIO_FPGA_SoC_2_wire\ <= GPIO_FPGA_SoC_2;
    \VCCIN_VR_PROCHOT_FPGA_wire\ <= VCCIN_VR_PROCHOT_FPGA;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    \CPU_C10_GATE_N_wire\ <= CPU_C10_GATE_N;
    VCCST_EN <= \VCCST_EN_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \TPM_GPIO_wire\ <= TPM_GPIO;
    SUSWARN_N <= \SUSWARN_N_wire\;
    \PLTRSTn_wire\ <= PLTRSTn;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    \V5A_OK_wire\ <= V5A_OK;
    RSMRSTn <= \RSMRSTn_wire\;
    \FPGA_OSC_wire\ <= FPGA_OSC;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \SPI_FP_IO2_wire\ <= SPI_FP_IO2;
    \SATAXPCIE1_FPGA_wire\ <= SATAXPCIE1_FPGA;
    \GPIO_FPGA_EXP_1_wire\ <= GPIO_FPGA_EXP_1;
    \VCCINAUX_VR_PROCHOT_FPGA_wire\ <= VCCINAUX_VR_PROCHOT_FPGA;
    VCCINAUX_VR_PE <= \VCCINAUX_VR_PE_wire\;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    \GPIO_FPGA_EXP_2_wire\ <= GPIO_FPGA_EXP_2;
    VPP_EN <= \VPP_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    \SUSACK_N_wire\ <= SUSACK_N;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    DSW_PWROK <= \DSW_PWROK_wire\;
    V5A_EN <= \V5A_EN_wire\;
    \GPIO_FPGA_SoC_3_wire\ <= GPIO_FPGA_SoC_3;
    \VR_PROCHOT_FPGA_OUT_N_wire\ <= VR_PROCHOT_FPGA_OUT_N;
    \VPP_OK_wire\ <= VPP_OK;
    VCCIN_VR_PE <= \VCCIN_VR_PE_wire\;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \SOC_SPKR_wire\ <= SOC_SPKR;
    \SLP_S5n_wire\ <= SLP_S5n;
    \V12_MAIN_MON_wire\ <= V12_MAIN_MON;
    \SPI_FP_IO3_wire\ <= SPI_FP_IO3;
    \SATAXPCIE0_FPGA_wire\ <= SATAXPCIE0_FPGA;
    \V33A_OK_wire\ <= V33A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    \FPGA_SLP_WLAN_N_wire\ <= FPGA_SLP_WLAN_N;

    \ipInertedIOPad_VR_READY_VCCINAUX_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__21309\,
            DIN => \N__21308\,
            DOUT => \N__21307\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \ipInertedIOPad_VR_READY_VCCINAUX_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21309\,
            PADOUT => \N__21308\,
            PADIN => \N__21307\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21300\,
            DIN => \N__21299\,
            DOUT => \N__21298\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \ipInertedIOPad_V33A_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21300\,
            PADOUT => \N__21299\,
            PADIN => \N__21298\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21291\,
            DIN => \N__21290\,
            DOUT => \N__21289\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \ipInertedIOPad_V1P8A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21291\,
            PADOUT => \N__21290\,
            PADIN => \N__21289\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17852\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21282\,
            DIN => \N__21281\,
            DOUT => \N__21280\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \ipInertedIOPad_VDDQ_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21282\,
            PADOUT => \N__21281\,
            PADIN => \N__21280\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__11063\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21273\,
            DIN => \N__21272\,
            DOUT => \N__21271\,
            PACKAGEPIN => \VCCST_OVERRIDE_3V3_wire\
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21273\,
            PADOUT => \N__21272\,
            PADIN => \N__21271\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21264\,
            DIN => \N__21263\,
            DOUT => \N__21262\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \ipInertedIOPad_V5S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21264\,
            PADOUT => \N__21263\,
            PADIN => \N__21262\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S3n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21255\,
            DIN => \N__21254\,
            DOUT => \N__21253\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \ipInertedIOPad_SLP_S3n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21255\,
            PADOUT => \N__21254\,
            PADIN => \N__21253\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s3n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S0n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21246\,
            DIN => \N__21245\,
            DOUT => \N__21244\,
            PACKAGEPIN => \SLP_S0n_wire\
        );

    \ipInertedIOPad_SLP_S0n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21246\,
            PADOUT => \N__21245\,
            PADIN => \N__21244\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21237\,
            DIN => \N__21236\,
            DOUT => \N__21235\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \ipInertedIOPad_V5S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21237\,
            PADOUT => \N__21236\,
            PADIN => \N__21235\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__11573\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__21228\,
            DIN => \N__21227\,
            DOUT => \N__21226\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \ipInertedIOPad_V1P8A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21228\,
            PADOUT => \N__21227\,
            PADIN => \N__21226\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v1p8a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTNn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21219\,
            DIN => \N__21218\,
            DOUT => \N__21217\,
            PACKAGEPIN => \PWRBTNn_wire\
        );

    \ipInertedIOPad_PWRBTNn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21219\,
            PADOUT => \N__21218\,
            PADIN => \N__21217\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTN_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21210\,
            DIN => \N__21209\,
            DOUT => \N__21208\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \ipInertedIOPad_PWRBTN_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21210\,
            PADOUT => \N__21209\,
            PADIN => \N__21208\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__9542\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21201\,
            DIN => \N__21200\,
            DOUT => \N__21199\,
            PACKAGEPIN => \GPIO_FPGA_SoC_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21201\,
            PADOUT => \N__21200\,
            PADIN => \N__21199\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21192\,
            DIN => \N__21191\,
            DOUT => \N__21190\,
            PACKAGEPIN => \VCCIN_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21192\,
            PADOUT => \N__21191\,
            PADIN => \N__21190\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_SUSn_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__21183\,
            DIN => \N__21182\,
            DOUT => \N__21181\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \ipInertedIOPad_SLP_SUSn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21183\,
            PADOUT => \N__21182\,
            PADIN => \N__21181\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_susn,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CPU_C10_GATE_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21174\,
            DIN => \N__21173\,
            DOUT => \N__21172\,
            PACKAGEPIN => \CPU_C10_GATE_N_wire\
        );

    \ipInertedIOPad_CPU_C10_GATE_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21174\,
            PADOUT => \N__21173\,
            PADIN => \N__21172\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21165\,
            DIN => \N__21164\,
            DOUT => \N__21163\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \ipInertedIOPad_VCCST_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21165\,
            PADOUT => \N__21164\,
            PADIN => \N__21163\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__15023\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33DSW_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__21156\,
            DIN => \N__21155\,
            DOUT => \N__21154\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \ipInertedIOPad_V33DSW_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21156\,
            PADOUT => \N__21155\,
            PADIN => \N__21154\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TPM_GPIO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21147\,
            DIN => \N__21146\,
            DOUT => \N__21145\,
            PACKAGEPIN => \TPM_GPIO_wire\
        );

    \ipInertedIOPad_TPM_GPIO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21147\,
            PADOUT => \N__21146\,
            PADIN => \N__21145\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSWARN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21138\,
            DIN => \N__21137\,
            DOUT => \N__21136\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \ipInertedIOPad_SUSWARN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21138\,
            PADOUT => \N__21137\,
            PADIN => \N__21136\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16592\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PLTRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21129\,
            DIN => \N__21128\,
            DOUT => \N__21127\,
            PACKAGEPIN => \PLTRSTn_wire\
        );

    \ipInertedIOPad_PLTRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21129\,
            PADOUT => \N__21128\,
            PADIN => \N__21127\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21120\,
            DIN => \N__21119\,
            DOUT => \N__21118\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21120\,
            PADOUT => \N__21119\,
            PADIN => \N__21118\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_4,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_READY_VCCIN_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__21111\,
            DIN => \N__21110\,
            DOUT => \N__21109\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \ipInertedIOPad_VR_READY_VCCIN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21111\,
            PADOUT => \N__21110\,
            PADIN => \N__21109\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccin,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__21102\,
            DIN => \N__21101\,
            DOUT => \N__21100\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \ipInertedIOPad_V5A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21102\,
            PADOUT => \N__21101\,
            PADIN => \N__21100\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RSMRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21093\,
            DIN => \N__21092\,
            DOUT => \N__21091\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \ipInertedIOPad_RSMRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21093\,
            PADOUT => \N__21092\,
            PADIN => \N__21091\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20717\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_OSC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21084\,
            DIN => \N__21083\,
            DOUT => \N__21082\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \ipInertedIOPad_FPGA_OSC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21084\,
            PADOUT => \N__21083\,
            PADIN => \N__21082\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => fpga_osc,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_PWRGD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21075\,
            DIN => \N__21074\,
            DOUT => \N__21073\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \ipInertedIOPad_VCCST_PWRGD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21075\,
            PADOUT => \N__21074\,
            PADIN => \N__21073\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19285\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SYS_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21066\,
            DIN => \N__21065\,
            DOUT => \N__21064\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \ipInertedIOPad_SYS_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21066\,
            PADOUT => \N__21065\,
            PADIN => \N__21064\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__11033\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21057\,
            DIN => \N__21056\,
            DOUT => \N__21055\,
            PACKAGEPIN => \SPI_FP_IO2_wire\
        );

    \ipInertedIOPad_SPI_FP_IO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21057\,
            PADOUT => \N__21056\,
            PADIN => \N__21055\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21048\,
            DIN => \N__21047\,
            DOUT => \N__21046\,
            PACKAGEPIN => \SATAXPCIE1_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21048\,
            PADOUT => \N__21047\,
            PADIN => \N__21046\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21039\,
            DIN => \N__21038\,
            DOUT => \N__21037\,
            PACKAGEPIN => \GPIO_FPGA_EXP_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21039\,
            PADOUT => \N__21038\,
            PADIN => \N__21037\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21030\,
            DIN => \N__21029\,
            DOUT => \N__21028\,
            PACKAGEPIN => \VCCINAUX_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21030\,
            PADOUT => \N__21029\,
            PADIN => \N__21028\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21021\,
            DIN => \N__21020\,
            DOUT => \N__21019\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21021\,
            PADOUT => \N__21020\,
            PADIN => \N__21019\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_HDA_SDO_ATP_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21012\,
            DIN => \N__21011\,
            DOUT => \N__21010\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \ipInertedIOPad_HDA_SDO_ATP_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21012\,
            PADOUT => \N__21011\,
            PADIN => \N__21010\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__11681\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__21003\,
            DIN => \N__21002\,
            DOUT => \N__21001\,
            PACKAGEPIN => \GPIO_FPGA_EXP_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__21003\,
            PADOUT => \N__21002\,
            PADIN => \N__21001\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20994\,
            DIN => \N__20993\,
            DOUT => \N__20992\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \ipInertedIOPad_VPP_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20994\,
            PADOUT => \N__20993\,
            PADIN => \N__20992\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__14969\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__20985\,
            DIN => \N__20984\,
            DOUT => \N__20983\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \ipInertedIOPad_VDDQ_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20985\,
            PADOUT => \N__20984\,
            PADIN => \N__20983\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vddq_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSACK_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20976\,
            DIN => \N__20975\,
            DOUT => \N__20974\,
            PACKAGEPIN => \SUSACK_N_wire\
        );

    \ipInertedIOPad_SUSACK_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20976\,
            PADOUT => \N__20975\,
            PADIN => \N__20974\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S4n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20967\,
            DIN => \N__20966\,
            DOUT => \N__20965\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \ipInertedIOPad_SLP_S4n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20967\,
            PADOUT => \N__20966\,
            PADIN => \N__20965\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s4n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_CPU_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20958\,
            DIN => \N__20957\,
            DOUT => \N__20956\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \ipInertedIOPad_VCCST_CPU_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20958\,
            PADOUT => \N__20957\,
            PADIN => \N__20956\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vccst_cpu_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20949\,
            DIN => \N__20948\,
            DOUT => \N__20947\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \ipInertedIOPad_VCCINAUX_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20949\,
            PADOUT => \N__20948\,
            PADIN => \N__20947\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17783\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20940\,
            DIN => \N__20939\,
            DOUT => \N__20938\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \ipInertedIOPad_V33S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20940\,
            PADOUT => \N__20939\,
            PADIN => \N__20938\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20931\,
            DIN => \N__20930\,
            DOUT => \N__20929\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \ipInertedIOPad_V33S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20931\,
            PADOUT => \N__20930\,
            PADIN => \N__20929\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__11569\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20922\,
            DIN => \N__20921\,
            DOUT => \N__20920\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20922\,
            PADOUT => \N__20921\,
            PADIN => \N__20920\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_1,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DSW_PWROK_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__20913\,
            DIN => \N__20912\,
            DOUT => \N__20911\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \ipInertedIOPad_DSW_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20913\,
            PADOUT => \N__20912\,
            PADIN => \N__20911\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__18374\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20904\,
            DIN => \N__20903\,
            DOUT => \N__20902\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \ipInertedIOPad_V5A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20904\,
            PADOUT => \N__20903\,
            PADIN => \N__20902\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17848\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20895\,
            DIN => \N__20894\,
            DOUT => \N__20893\,
            PACKAGEPIN => \GPIO_FPGA_SoC_3_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20895\,
            PADOUT => \N__20894\,
            PADIN => \N__20893\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20886\,
            DIN => \N__20885\,
            DOUT => \N__20884\,
            PACKAGEPIN => \VR_PROCHOT_FPGA_OUT_N_wire\
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20886\,
            PADOUT => \N__20885\,
            PADIN => \N__20884\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__20877\,
            DIN => \N__20876\,
            DOUT => \N__20875\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \ipInertedIOPad_VPP_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20877\,
            PADOUT => \N__20876\,
            PADIN => \N__20875\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vpp_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20868\,
            DIN => \N__20867\,
            DOUT => \N__20866\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20868\,
            PADOUT => \N__20867\,
            PADIN => \N__20866\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20859\,
            DIN => \N__20858\,
            DOUT => \N__20857\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \ipInertedIOPad_VCCIN_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20859\,
            PADOUT => \N__20858\,
            PADIN => \N__20857\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19284\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SOC_SPKR_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20850\,
            DIN => \N__20849\,
            DOUT => \N__20848\,
            PACKAGEPIN => \SOC_SPKR_wire\
        );

    \ipInertedIOPad_SOC_SPKR_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20850\,
            PADOUT => \N__20849\,
            PADIN => \N__20848\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S5n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20841\,
            DIN => \N__20840\,
            DOUT => \N__20839\,
            PACKAGEPIN => \SLP_S5n_wire\
        );

    \ipInertedIOPad_SLP_S5n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20841\,
            PADOUT => \N__20840\,
            PADIN => \N__20839\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V12_MAIN_MON_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20832\,
            DIN => \N__20831\,
            DOUT => \N__20830\,
            PACKAGEPIN => \V12_MAIN_MON_wire\
        );

    \ipInertedIOPad_V12_MAIN_MON_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20832\,
            PADOUT => \N__20831\,
            PADIN => \N__20830\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20823\,
            DIN => \N__20822\,
            DOUT => \N__20821\,
            PACKAGEPIN => \SPI_FP_IO3_wire\
        );

    \ipInertedIOPad_SPI_FP_IO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20823\,
            PADOUT => \N__20822\,
            PADIN => \N__20821\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20814\,
            DIN => \N__20813\,
            DOUT => \N__20812\,
            PACKAGEPIN => \SATAXPCIE0_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20814\,
            PADOUT => \N__20813\,
            PADIN => \N__20812\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20805\,
            DIN => \N__20804\,
            DOUT => \N__20803\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \ipInertedIOPad_V33A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20805\,
            PADOUT => \N__20804\,
            PADIN => \N__20803\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PCH_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20796\,
            DIN => \N__20795\,
            DOUT => \N__20794\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \ipInertedIOPad_PCH_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20796\,
            PADOUT => \N__20795\,
            PADIN => \N__20794\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__11025\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__20787\,
            DIN => \N__20786\,
            DOUT => \N__20785\,
            PACKAGEPIN => \FPGA_SLP_WLAN_N_wire\
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__20787\,
            PADOUT => \N__20786\,
            PADIN => \N__20785\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__4744\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20765\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__20765\,
            I => \N__20761\
        );

    \I__4742\ : InMux
    port map (
            O => \N__20764\,
            I => \N__20758\
        );

    \I__4741\ : Span4Mux_s2_h
    port map (
            O => \N__20761\,
            I => \N__20755\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__20758\,
            I => \N__20752\
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__20755\,
            I => \RSMRST_PWRGD.N_240\
        );

    \I__4738\ : Odrv12
    port map (
            O => \N__20752\,
            I => \RSMRST_PWRGD.N_240\
        );

    \I__4737\ : InMux
    port map (
            O => \N__20747\,
            I => \N__20740\
        );

    \I__4736\ : InMux
    port map (
            O => \N__20746\,
            I => \N__20737\
        );

    \I__4735\ : InMux
    port map (
            O => \N__20745\,
            I => \N__20734\
        );

    \I__4734\ : InMux
    port map (
            O => \N__20744\,
            I => \N__20729\
        );

    \I__4733\ : InMux
    port map (
            O => \N__20743\,
            I => \N__20729\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__20740\,
            I => \N__20724\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__20737\,
            I => \N__20724\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__20734\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__20729\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__4728\ : Odrv4
    port map (
            O => \N__20724\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__4727\ : IoInMux
    port map (
            O => \N__20717\,
            I => \N__20712\
        );

    \I__4726\ : InMux
    port map (
            O => \N__20716\,
            I => \N__20709\
        );

    \I__4725\ : InMux
    port map (
            O => \N__20715\,
            I => \N__20705\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__20712\,
            I => \N__20699\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__20709\,
            I => \N__20696\
        );

    \I__4722\ : InMux
    port map (
            O => \N__20708\,
            I => \N__20693\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__20705\,
            I => \N__20690\
        );

    \I__4720\ : InMux
    port map (
            O => \N__20704\,
            I => \N__20687\
        );

    \I__4719\ : InMux
    port map (
            O => \N__20703\,
            I => \N__20684\
        );

    \I__4718\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20681\
        );

    \I__4717\ : IoSpan4Mux
    port map (
            O => \N__20699\,
            I => \N__20678\
        );

    \I__4716\ : Span4Mux_h
    port map (
            O => \N__20696\,
            I => \N__20675\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__20693\,
            I => \N__20672\
        );

    \I__4714\ : Span4Mux_v
    port map (
            O => \N__20690\,
            I => \N__20663\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__20687\,
            I => \N__20663\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__20684\,
            I => \N__20663\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__20681\,
            I => \N__20663\
        );

    \I__4710\ : IoSpan4Mux
    port map (
            O => \N__20678\,
            I => \N__20660\
        );

    \I__4709\ : Span4Mux_v
    port map (
            O => \N__20675\,
            I => \N__20657\
        );

    \I__4708\ : Span12Mux_s10_h
    port map (
            O => \N__20672\,
            I => \N__20654\
        );

    \I__4707\ : Span4Mux_v
    port map (
            O => \N__20663\,
            I => \N__20651\
        );

    \I__4706\ : Odrv4
    port map (
            O => \N__20660\,
            I => rsmrstn
        );

    \I__4705\ : Odrv4
    port map (
            O => \N__20657\,
            I => rsmrstn
        );

    \I__4704\ : Odrv12
    port map (
            O => \N__20654\,
            I => rsmrstn
        );

    \I__4703\ : Odrv4
    port map (
            O => \N__20651\,
            I => rsmrstn
        );

    \I__4702\ : ClkMux
    port map (
            O => \N__20642\,
            I => \N__20638\
        );

    \I__4701\ : ClkMux
    port map (
            O => \N__20641\,
            I => \N__20632\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__20638\,
            I => \N__20625\
        );

    \I__4699\ : ClkMux
    port map (
            O => \N__20637\,
            I => \N__20622\
        );

    \I__4698\ : ClkMux
    port map (
            O => \N__20636\,
            I => \N__20619\
        );

    \I__4697\ : ClkMux
    port map (
            O => \N__20635\,
            I => \N__20616\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__20632\,
            I => \N__20612\
        );

    \I__4695\ : ClkMux
    port map (
            O => \N__20631\,
            I => \N__20609\
        );

    \I__4694\ : ClkMux
    port map (
            O => \N__20630\,
            I => \N__20606\
        );

    \I__4693\ : ClkMux
    port map (
            O => \N__20629\,
            I => \N__20601\
        );

    \I__4692\ : ClkMux
    port map (
            O => \N__20628\,
            I => \N__20597\
        );

    \I__4691\ : Span4Mux_s3_v
    port map (
            O => \N__20625\,
            I => \N__20586\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__20622\,
            I => \N__20586\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__20619\,
            I => \N__20586\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__20616\,
            I => \N__20582\
        );

    \I__4687\ : ClkMux
    port map (
            O => \N__20615\,
            I => \N__20579\
        );

    \I__4686\ : Span4Mux_s3_v
    port map (
            O => \N__20612\,
            I => \N__20574\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__20609\,
            I => \N__20574\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__20606\,
            I => \N__20571\
        );

    \I__4683\ : ClkMux
    port map (
            O => \N__20605\,
            I => \N__20568\
        );

    \I__4682\ : ClkMux
    port map (
            O => \N__20604\,
            I => \N__20565\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__20601\,
            I => \N__20561\
        );

    \I__4680\ : ClkMux
    port map (
            O => \N__20600\,
            I => \N__20554\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__20597\,
            I => \N__20551\
        );

    \I__4678\ : ClkMux
    port map (
            O => \N__20596\,
            I => \N__20548\
        );

    \I__4677\ : ClkMux
    port map (
            O => \N__20595\,
            I => \N__20544\
        );

    \I__4676\ : ClkMux
    port map (
            O => \N__20594\,
            I => \N__20539\
        );

    \I__4675\ : ClkMux
    port map (
            O => \N__20593\,
            I => \N__20535\
        );

    \I__4674\ : Span4Mux_v
    port map (
            O => \N__20586\,
            I => \N__20529\
        );

    \I__4673\ : ClkMux
    port map (
            O => \N__20585\,
            I => \N__20526\
        );

    \I__4672\ : Span4Mux_s3_v
    port map (
            O => \N__20582\,
            I => \N__20521\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__20579\,
            I => \N__20521\
        );

    \I__4670\ : Span4Mux_v
    port map (
            O => \N__20574\,
            I => \N__20518\
        );

    \I__4669\ : Span4Mux_s3_v
    port map (
            O => \N__20571\,
            I => \N__20511\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__20568\,
            I => \N__20511\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__20565\,
            I => \N__20511\
        );

    \I__4666\ : ClkMux
    port map (
            O => \N__20564\,
            I => \N__20508\
        );

    \I__4665\ : Span4Mux_v
    port map (
            O => \N__20561\,
            I => \N__20505\
        );

    \I__4664\ : ClkMux
    port map (
            O => \N__20560\,
            I => \N__20502\
        );

    \I__4663\ : ClkMux
    port map (
            O => \N__20559\,
            I => \N__20499\
        );

    \I__4662\ : ClkMux
    port map (
            O => \N__20558\,
            I => \N__20496\
        );

    \I__4661\ : ClkMux
    port map (
            O => \N__20557\,
            I => \N__20492\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__20554\,
            I => \N__20488\
        );

    \I__4659\ : Span4Mux_s2_h
    port map (
            O => \N__20551\,
            I => \N__20483\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__20548\,
            I => \N__20483\
        );

    \I__4657\ : ClkMux
    port map (
            O => \N__20547\,
            I => \N__20480\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__20544\,
            I => \N__20477\
        );

    \I__4655\ : ClkMux
    port map (
            O => \N__20543\,
            I => \N__20474\
        );

    \I__4654\ : ClkMux
    port map (
            O => \N__20542\,
            I => \N__20468\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__20539\,
            I => \N__20462\
        );

    \I__4652\ : ClkMux
    port map (
            O => \N__20538\,
            I => \N__20459\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__20535\,
            I => \N__20455\
        );

    \I__4650\ : ClkMux
    port map (
            O => \N__20534\,
            I => \N__20452\
        );

    \I__4649\ : ClkMux
    port map (
            O => \N__20533\,
            I => \N__20447\
        );

    \I__4648\ : ClkMux
    port map (
            O => \N__20532\,
            I => \N__20444\
        );

    \I__4647\ : Span4Mux_h
    port map (
            O => \N__20529\,
            I => \N__20438\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__20526\,
            I => \N__20438\
        );

    \I__4645\ : Span4Mux_v
    port map (
            O => \N__20521\,
            I => \N__20429\
        );

    \I__4644\ : Span4Mux_h
    port map (
            O => \N__20518\,
            I => \N__20429\
        );

    \I__4643\ : Span4Mux_v
    port map (
            O => \N__20511\,
            I => \N__20429\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__20508\,
            I => \N__20429\
        );

    \I__4641\ : Span4Mux_v
    port map (
            O => \N__20505\,
            I => \N__20423\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__20502\,
            I => \N__20423\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__20499\,
            I => \N__20418\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__20496\,
            I => \N__20418\
        );

    \I__4637\ : ClkMux
    port map (
            O => \N__20495\,
            I => \N__20415\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__20492\,
            I => \N__20412\
        );

    \I__4635\ : ClkMux
    port map (
            O => \N__20491\,
            I => \N__20409\
        );

    \I__4634\ : Span4Mux_h
    port map (
            O => \N__20488\,
            I => \N__20404\
        );

    \I__4633\ : Span4Mux_h
    port map (
            O => \N__20483\,
            I => \N__20399\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__20480\,
            I => \N__20399\
        );

    \I__4631\ : Span4Mux_v
    port map (
            O => \N__20477\,
            I => \N__20394\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__20474\,
            I => \N__20394\
        );

    \I__4629\ : ClkMux
    port map (
            O => \N__20473\,
            I => \N__20391\
        );

    \I__4628\ : ClkMux
    port map (
            O => \N__20472\,
            I => \N__20388\
        );

    \I__4627\ : ClkMux
    port map (
            O => \N__20471\,
            I => \N__20385\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__20468\,
            I => \N__20381\
        );

    \I__4625\ : ClkMux
    port map (
            O => \N__20467\,
            I => \N__20378\
        );

    \I__4624\ : ClkMux
    port map (
            O => \N__20466\,
            I => \N__20374\
        );

    \I__4623\ : ClkMux
    port map (
            O => \N__20465\,
            I => \N__20371\
        );

    \I__4622\ : Span4Mux_v
    port map (
            O => \N__20462\,
            I => \N__20365\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__20459\,
            I => \N__20365\
        );

    \I__4620\ : ClkMux
    port map (
            O => \N__20458\,
            I => \N__20362\
        );

    \I__4619\ : Span4Mux_s3_v
    port map (
            O => \N__20455\,
            I => \N__20357\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__20452\,
            I => \N__20357\
        );

    \I__4617\ : ClkMux
    port map (
            O => \N__20451\,
            I => \N__20354\
        );

    \I__4616\ : ClkMux
    port map (
            O => \N__20450\,
            I => \N__20351\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__20447\,
            I => \N__20348\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__20444\,
            I => \N__20345\
        );

    \I__4613\ : ClkMux
    port map (
            O => \N__20443\,
            I => \N__20342\
        );

    \I__4612\ : Span4Mux_v
    port map (
            O => \N__20438\,
            I => \N__20336\
        );

    \I__4611\ : Span4Mux_v
    port map (
            O => \N__20429\,
            I => \N__20336\
        );

    \I__4610\ : ClkMux
    port map (
            O => \N__20428\,
            I => \N__20333\
        );

    \I__4609\ : Span4Mux_v
    port map (
            O => \N__20423\,
            I => \N__20330\
        );

    \I__4608\ : Span4Mux_v
    port map (
            O => \N__20418\,
            I => \N__20325\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__20415\,
            I => \N__20325\
        );

    \I__4606\ : Span4Mux_h
    port map (
            O => \N__20412\,
            I => \N__20320\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__20409\,
            I => \N__20320\
        );

    \I__4604\ : ClkMux
    port map (
            O => \N__20408\,
            I => \N__20317\
        );

    \I__4603\ : ClkMux
    port map (
            O => \N__20407\,
            I => \N__20314\
        );

    \I__4602\ : Span4Mux_v
    port map (
            O => \N__20404\,
            I => \N__20305\
        );

    \I__4601\ : Span4Mux_v
    port map (
            O => \N__20399\,
            I => \N__20305\
        );

    \I__4600\ : Span4Mux_h
    port map (
            O => \N__20394\,
            I => \N__20305\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__20391\,
            I => \N__20305\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__20388\,
            I => \N__20302\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__20385\,
            I => \N__20299\
        );

    \I__4596\ : ClkMux
    port map (
            O => \N__20384\,
            I => \N__20296\
        );

    \I__4595\ : Span4Mux_v
    port map (
            O => \N__20381\,
            I => \N__20291\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__20378\,
            I => \N__20291\
        );

    \I__4593\ : ClkMux
    port map (
            O => \N__20377\,
            I => \N__20288\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__20374\,
            I => \N__20285\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__20371\,
            I => \N__20282\
        );

    \I__4590\ : ClkMux
    port map (
            O => \N__20370\,
            I => \N__20279\
        );

    \I__4589\ : Span4Mux_v
    port map (
            O => \N__20365\,
            I => \N__20274\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__20362\,
            I => \N__20274\
        );

    \I__4587\ : Span4Mux_v
    port map (
            O => \N__20357\,
            I => \N__20265\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__20354\,
            I => \N__20265\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__20351\,
            I => \N__20265\
        );

    \I__4584\ : Span4Mux_h
    port map (
            O => \N__20348\,
            I => \N__20265\
        );

    \I__4583\ : Span4Mux_v
    port map (
            O => \N__20345\,
            I => \N__20260\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__20342\,
            I => \N__20260\
        );

    \I__4581\ : ClkMux
    port map (
            O => \N__20341\,
            I => \N__20257\
        );

    \I__4580\ : Span4Mux_v
    port map (
            O => \N__20336\,
            I => \N__20254\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__20333\,
            I => \N__20251\
        );

    \I__4578\ : IoSpan4Mux
    port map (
            O => \N__20330\,
            I => \N__20248\
        );

    \I__4577\ : Span4Mux_v
    port map (
            O => \N__20325\,
            I => \N__20241\
        );

    \I__4576\ : Span4Mux_v
    port map (
            O => \N__20320\,
            I => \N__20241\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__20317\,
            I => \N__20241\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__20314\,
            I => \N__20238\
        );

    \I__4573\ : Span4Mux_v
    port map (
            O => \N__20305\,
            I => \N__20233\
        );

    \I__4572\ : Span4Mux_h
    port map (
            O => \N__20302\,
            I => \N__20233\
        );

    \I__4571\ : Span4Mux_h
    port map (
            O => \N__20299\,
            I => \N__20228\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__20296\,
            I => \N__20228\
        );

    \I__4569\ : Span4Mux_h
    port map (
            O => \N__20291\,
            I => \N__20223\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__20288\,
            I => \N__20223\
        );

    \I__4567\ : Span4Mux_s2_h
    port map (
            O => \N__20285\,
            I => \N__20216\
        );

    \I__4566\ : Span4Mux_h
    port map (
            O => \N__20282\,
            I => \N__20216\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__20279\,
            I => \N__20216\
        );

    \I__4564\ : Span4Mux_h
    port map (
            O => \N__20274\,
            I => \N__20207\
        );

    \I__4563\ : Span4Mux_v
    port map (
            O => \N__20265\,
            I => \N__20207\
        );

    \I__4562\ : Span4Mux_h
    port map (
            O => \N__20260\,
            I => \N__20207\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__20257\,
            I => \N__20207\
        );

    \I__4560\ : IoSpan4Mux
    port map (
            O => \N__20254\,
            I => \N__20202\
        );

    \I__4559\ : Span4Mux_h
    port map (
            O => \N__20251\,
            I => \N__20199\
        );

    \I__4558\ : IoSpan4Mux
    port map (
            O => \N__20248\,
            I => \N__20192\
        );

    \I__4557\ : IoSpan4Mux
    port map (
            O => \N__20241\,
            I => \N__20192\
        );

    \I__4556\ : IoSpan4Mux
    port map (
            O => \N__20238\,
            I => \N__20192\
        );

    \I__4555\ : Span4Mux_v
    port map (
            O => \N__20233\,
            I => \N__20183\
        );

    \I__4554\ : Span4Mux_v
    port map (
            O => \N__20228\,
            I => \N__20183\
        );

    \I__4553\ : Span4Mux_h
    port map (
            O => \N__20223\,
            I => \N__20183\
        );

    \I__4552\ : Span4Mux_h
    port map (
            O => \N__20216\,
            I => \N__20183\
        );

    \I__4551\ : Sp12to4
    port map (
            O => \N__20207\,
            I => \N__20180\
        );

    \I__4550\ : ClkMux
    port map (
            O => \N__20206\,
            I => \N__20177\
        );

    \I__4549\ : ClkMux
    port map (
            O => \N__20205\,
            I => \N__20174\
        );

    \I__4548\ : Odrv4
    port map (
            O => \N__20202\,
            I => fpga_osc
        );

    \I__4547\ : Odrv4
    port map (
            O => \N__20199\,
            I => fpga_osc
        );

    \I__4546\ : Odrv4
    port map (
            O => \N__20192\,
            I => fpga_osc
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__20183\,
            I => fpga_osc
        );

    \I__4544\ : Odrv12
    port map (
            O => \N__20180\,
            I => fpga_osc
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__20177\,
            I => fpga_osc
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__20174\,
            I => fpga_osc
        );

    \I__4541\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20047\
        );

    \I__4540\ : InMux
    port map (
            O => \N__20158\,
            I => \N__20047\
        );

    \I__4539\ : InMux
    port map (
            O => \N__20157\,
            I => \N__20047\
        );

    \I__4538\ : InMux
    port map (
            O => \N__20156\,
            I => \N__20047\
        );

    \I__4537\ : InMux
    port map (
            O => \N__20155\,
            I => \N__20040\
        );

    \I__4536\ : InMux
    port map (
            O => \N__20154\,
            I => \N__20040\
        );

    \I__4535\ : InMux
    port map (
            O => \N__20153\,
            I => \N__20040\
        );

    \I__4534\ : InMux
    port map (
            O => \N__20152\,
            I => \N__20033\
        );

    \I__4533\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20033\
        );

    \I__4532\ : InMux
    port map (
            O => \N__20150\,
            I => \N__20033\
        );

    \I__4531\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20024\
        );

    \I__4530\ : InMux
    port map (
            O => \N__20148\,
            I => \N__20024\
        );

    \I__4529\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20024\
        );

    \I__4528\ : InMux
    port map (
            O => \N__20146\,
            I => \N__20024\
        );

    \I__4527\ : InMux
    port map (
            O => \N__20145\,
            I => \N__20015\
        );

    \I__4526\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20015\
        );

    \I__4525\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20015\
        );

    \I__4524\ : InMux
    port map (
            O => \N__20142\,
            I => \N__20015\
        );

    \I__4523\ : InMux
    port map (
            O => \N__20141\,
            I => \N__20008\
        );

    \I__4522\ : InMux
    port map (
            O => \N__20140\,
            I => \N__20008\
        );

    \I__4521\ : InMux
    port map (
            O => \N__20139\,
            I => \N__20008\
        );

    \I__4520\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20001\
        );

    \I__4519\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20001\
        );

    \I__4518\ : InMux
    port map (
            O => \N__20136\,
            I => \N__20001\
        );

    \I__4517\ : InMux
    port map (
            O => \N__20135\,
            I => \N__19992\
        );

    \I__4516\ : InMux
    port map (
            O => \N__20134\,
            I => \N__19992\
        );

    \I__4515\ : InMux
    port map (
            O => \N__20133\,
            I => \N__19992\
        );

    \I__4514\ : InMux
    port map (
            O => \N__20132\,
            I => \N__19992\
        );

    \I__4513\ : InMux
    port map (
            O => \N__20131\,
            I => \N__19983\
        );

    \I__4512\ : InMux
    port map (
            O => \N__20130\,
            I => \N__19983\
        );

    \I__4511\ : InMux
    port map (
            O => \N__20129\,
            I => \N__19983\
        );

    \I__4510\ : InMux
    port map (
            O => \N__20128\,
            I => \N__19983\
        );

    \I__4509\ : InMux
    port map (
            O => \N__20127\,
            I => \N__19974\
        );

    \I__4508\ : InMux
    port map (
            O => \N__20126\,
            I => \N__19974\
        );

    \I__4507\ : InMux
    port map (
            O => \N__20125\,
            I => \N__19974\
        );

    \I__4506\ : InMux
    port map (
            O => \N__20124\,
            I => \N__19974\
        );

    \I__4505\ : InMux
    port map (
            O => \N__20123\,
            I => \N__19969\
        );

    \I__4504\ : InMux
    port map (
            O => \N__20122\,
            I => \N__19969\
        );

    \I__4503\ : InMux
    port map (
            O => \N__20121\,
            I => \N__19960\
        );

    \I__4502\ : InMux
    port map (
            O => \N__20120\,
            I => \N__19960\
        );

    \I__4501\ : InMux
    port map (
            O => \N__20119\,
            I => \N__19960\
        );

    \I__4500\ : InMux
    port map (
            O => \N__20118\,
            I => \N__19960\
        );

    \I__4499\ : InMux
    port map (
            O => \N__20117\,
            I => \N__19951\
        );

    \I__4498\ : InMux
    port map (
            O => \N__20116\,
            I => \N__19951\
        );

    \I__4497\ : InMux
    port map (
            O => \N__20115\,
            I => \N__19951\
        );

    \I__4496\ : InMux
    port map (
            O => \N__20114\,
            I => \N__19951\
        );

    \I__4495\ : InMux
    port map (
            O => \N__20113\,
            I => \N__19942\
        );

    \I__4494\ : InMux
    port map (
            O => \N__20112\,
            I => \N__19942\
        );

    \I__4493\ : InMux
    port map (
            O => \N__20111\,
            I => \N__19942\
        );

    \I__4492\ : InMux
    port map (
            O => \N__20110\,
            I => \N__19942\
        );

    \I__4491\ : InMux
    port map (
            O => \N__20109\,
            I => \N__19935\
        );

    \I__4490\ : InMux
    port map (
            O => \N__20108\,
            I => \N__19935\
        );

    \I__4489\ : InMux
    port map (
            O => \N__20107\,
            I => \N__19935\
        );

    \I__4488\ : InMux
    port map (
            O => \N__20106\,
            I => \N__19926\
        );

    \I__4487\ : InMux
    port map (
            O => \N__20105\,
            I => \N__19926\
        );

    \I__4486\ : InMux
    port map (
            O => \N__20104\,
            I => \N__19926\
        );

    \I__4485\ : InMux
    port map (
            O => \N__20103\,
            I => \N__19926\
        );

    \I__4484\ : InMux
    port map (
            O => \N__20102\,
            I => \N__19919\
        );

    \I__4483\ : InMux
    port map (
            O => \N__20101\,
            I => \N__19919\
        );

    \I__4482\ : InMux
    port map (
            O => \N__20100\,
            I => \N__19919\
        );

    \I__4481\ : InMux
    port map (
            O => \N__20099\,
            I => \N__19910\
        );

    \I__4480\ : InMux
    port map (
            O => \N__20098\,
            I => \N__19910\
        );

    \I__4479\ : InMux
    port map (
            O => \N__20097\,
            I => \N__19910\
        );

    \I__4478\ : InMux
    port map (
            O => \N__20096\,
            I => \N__19910\
        );

    \I__4477\ : InMux
    port map (
            O => \N__20095\,
            I => \N__19901\
        );

    \I__4476\ : InMux
    port map (
            O => \N__20094\,
            I => \N__19901\
        );

    \I__4475\ : InMux
    port map (
            O => \N__20093\,
            I => \N__19901\
        );

    \I__4474\ : InMux
    port map (
            O => \N__20092\,
            I => \N__19901\
        );

    \I__4473\ : InMux
    port map (
            O => \N__20091\,
            I => \N__19894\
        );

    \I__4472\ : InMux
    port map (
            O => \N__20090\,
            I => \N__19894\
        );

    \I__4471\ : InMux
    port map (
            O => \N__20089\,
            I => \N__19894\
        );

    \I__4470\ : InMux
    port map (
            O => \N__20088\,
            I => \N__19885\
        );

    \I__4469\ : InMux
    port map (
            O => \N__20087\,
            I => \N__19885\
        );

    \I__4468\ : InMux
    port map (
            O => \N__20086\,
            I => \N__19885\
        );

    \I__4467\ : InMux
    port map (
            O => \N__20085\,
            I => \N__19885\
        );

    \I__4466\ : InMux
    port map (
            O => \N__20084\,
            I => \N__19880\
        );

    \I__4465\ : InMux
    port map (
            O => \N__20083\,
            I => \N__19880\
        );

    \I__4464\ : InMux
    port map (
            O => \N__20082\,
            I => \N__19871\
        );

    \I__4463\ : InMux
    port map (
            O => \N__20081\,
            I => \N__19871\
        );

    \I__4462\ : InMux
    port map (
            O => \N__20080\,
            I => \N__19871\
        );

    \I__4461\ : InMux
    port map (
            O => \N__20079\,
            I => \N__19871\
        );

    \I__4460\ : InMux
    port map (
            O => \N__20078\,
            I => \N__19868\
        );

    \I__4459\ : InMux
    port map (
            O => \N__20077\,
            I => \N__19859\
        );

    \I__4458\ : InMux
    port map (
            O => \N__20076\,
            I => \N__19859\
        );

    \I__4457\ : InMux
    port map (
            O => \N__20075\,
            I => \N__19859\
        );

    \I__4456\ : InMux
    port map (
            O => \N__20074\,
            I => \N__19859\
        );

    \I__4455\ : InMux
    port map (
            O => \N__20073\,
            I => \N__19852\
        );

    \I__4454\ : InMux
    port map (
            O => \N__20072\,
            I => \N__19852\
        );

    \I__4453\ : InMux
    port map (
            O => \N__20071\,
            I => \N__19852\
        );

    \I__4452\ : InMux
    port map (
            O => \N__20070\,
            I => \N__19843\
        );

    \I__4451\ : InMux
    port map (
            O => \N__20069\,
            I => \N__19843\
        );

    \I__4450\ : InMux
    port map (
            O => \N__20068\,
            I => \N__19843\
        );

    \I__4449\ : InMux
    port map (
            O => \N__20067\,
            I => \N__19843\
        );

    \I__4448\ : InMux
    port map (
            O => \N__20066\,
            I => \N__19840\
        );

    \I__4447\ : InMux
    port map (
            O => \N__20065\,
            I => \N__19835\
        );

    \I__4446\ : InMux
    port map (
            O => \N__20064\,
            I => \N__19835\
        );

    \I__4445\ : InMux
    port map (
            O => \N__20063\,
            I => \N__19832\
        );

    \I__4444\ : InMux
    port map (
            O => \N__20062\,
            I => \N__19829\
        );

    \I__4443\ : InMux
    port map (
            O => \N__20061\,
            I => \N__19826\
        );

    \I__4442\ : InMux
    port map (
            O => \N__20060\,
            I => \N__19821\
        );

    \I__4441\ : InMux
    port map (
            O => \N__20059\,
            I => \N__19821\
        );

    \I__4440\ : InMux
    port map (
            O => \N__20058\,
            I => \N__19816\
        );

    \I__4439\ : InMux
    port map (
            O => \N__20057\,
            I => \N__19816\
        );

    \I__4438\ : InMux
    port map (
            O => \N__20056\,
            I => \N__19813\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__20047\,
            I => \N__19803\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__20040\,
            I => \N__19799\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__20033\,
            I => \N__19794\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__20024\,
            I => \N__19791\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__20015\,
            I => \N__19788\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__20008\,
            I => \N__19781\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__20001\,
            I => \N__19778\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__19992\,
            I => \N__19775\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__19983\,
            I => \N__19770\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__19974\,
            I => \N__19767\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__19969\,
            I => \N__19764\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__19960\,
            I => \N__19759\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__19951\,
            I => \N__19756\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__19942\,
            I => \N__19753\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__19935\,
            I => \N__19750\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__19926\,
            I => \N__19746\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__19919\,
            I => \N__19743\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__19910\,
            I => \N__19737\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__19901\,
            I => \N__19734\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__19894\,
            I => \N__19731\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__19885\,
            I => \N__19728\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__19880\,
            I => \N__19725\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__19871\,
            I => \N__19722\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__19868\,
            I => \N__19719\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__19859\,
            I => \N__19716\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__19852\,
            I => \N__19713\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__19843\,
            I => \N__19709\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__19840\,
            I => \N__19706\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__19835\,
            I => \N__19703\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__19832\,
            I => \N__19700\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__19829\,
            I => \N__19697\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__19826\,
            I => \N__19694\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__19821\,
            I => \N__19691\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__19816\,
            I => \N__19688\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__19813\,
            I => \N__19685\
        );

    \I__4402\ : CEMux
    port map (
            O => \N__19812\,
            I => \N__19568\
        );

    \I__4401\ : CEMux
    port map (
            O => \N__19811\,
            I => \N__19568\
        );

    \I__4400\ : CEMux
    port map (
            O => \N__19810\,
            I => \N__19568\
        );

    \I__4399\ : CEMux
    port map (
            O => \N__19809\,
            I => \N__19568\
        );

    \I__4398\ : CEMux
    port map (
            O => \N__19808\,
            I => \N__19568\
        );

    \I__4397\ : CEMux
    port map (
            O => \N__19807\,
            I => \N__19568\
        );

    \I__4396\ : CEMux
    port map (
            O => \N__19806\,
            I => \N__19568\
        );

    \I__4395\ : Glb2LocalMux
    port map (
            O => \N__19803\,
            I => \N__19568\
        );

    \I__4394\ : CEMux
    port map (
            O => \N__19802\,
            I => \N__19568\
        );

    \I__4393\ : Glb2LocalMux
    port map (
            O => \N__19799\,
            I => \N__19568\
        );

    \I__4392\ : CEMux
    port map (
            O => \N__19798\,
            I => \N__19568\
        );

    \I__4391\ : CEMux
    port map (
            O => \N__19797\,
            I => \N__19568\
        );

    \I__4390\ : Glb2LocalMux
    port map (
            O => \N__19794\,
            I => \N__19568\
        );

    \I__4389\ : Glb2LocalMux
    port map (
            O => \N__19791\,
            I => \N__19568\
        );

    \I__4388\ : Glb2LocalMux
    port map (
            O => \N__19788\,
            I => \N__19568\
        );

    \I__4387\ : CEMux
    port map (
            O => \N__19787\,
            I => \N__19568\
        );

    \I__4386\ : CEMux
    port map (
            O => \N__19786\,
            I => \N__19568\
        );

    \I__4385\ : CEMux
    port map (
            O => \N__19785\,
            I => \N__19568\
        );

    \I__4384\ : CEMux
    port map (
            O => \N__19784\,
            I => \N__19568\
        );

    \I__4383\ : Glb2LocalMux
    port map (
            O => \N__19781\,
            I => \N__19568\
        );

    \I__4382\ : Glb2LocalMux
    port map (
            O => \N__19778\,
            I => \N__19568\
        );

    \I__4381\ : Glb2LocalMux
    port map (
            O => \N__19775\,
            I => \N__19568\
        );

    \I__4380\ : CEMux
    port map (
            O => \N__19774\,
            I => \N__19568\
        );

    \I__4379\ : CEMux
    port map (
            O => \N__19773\,
            I => \N__19568\
        );

    \I__4378\ : Glb2LocalMux
    port map (
            O => \N__19770\,
            I => \N__19568\
        );

    \I__4377\ : Glb2LocalMux
    port map (
            O => \N__19767\,
            I => \N__19568\
        );

    \I__4376\ : Glb2LocalMux
    port map (
            O => \N__19764\,
            I => \N__19568\
        );

    \I__4375\ : CEMux
    port map (
            O => \N__19763\,
            I => \N__19568\
        );

    \I__4374\ : CEMux
    port map (
            O => \N__19762\,
            I => \N__19568\
        );

    \I__4373\ : Glb2LocalMux
    port map (
            O => \N__19759\,
            I => \N__19568\
        );

    \I__4372\ : Glb2LocalMux
    port map (
            O => \N__19756\,
            I => \N__19568\
        );

    \I__4371\ : Glb2LocalMux
    port map (
            O => \N__19753\,
            I => \N__19568\
        );

    \I__4370\ : Glb2LocalMux
    port map (
            O => \N__19750\,
            I => \N__19568\
        );

    \I__4369\ : CEMux
    port map (
            O => \N__19749\,
            I => \N__19568\
        );

    \I__4368\ : Glb2LocalMux
    port map (
            O => \N__19746\,
            I => \N__19568\
        );

    \I__4367\ : Glb2LocalMux
    port map (
            O => \N__19743\,
            I => \N__19568\
        );

    \I__4366\ : CEMux
    port map (
            O => \N__19742\,
            I => \N__19568\
        );

    \I__4365\ : CEMux
    port map (
            O => \N__19741\,
            I => \N__19568\
        );

    \I__4364\ : CEMux
    port map (
            O => \N__19740\,
            I => \N__19568\
        );

    \I__4363\ : Glb2LocalMux
    port map (
            O => \N__19737\,
            I => \N__19568\
        );

    \I__4362\ : Glb2LocalMux
    port map (
            O => \N__19734\,
            I => \N__19568\
        );

    \I__4361\ : Glb2LocalMux
    port map (
            O => \N__19731\,
            I => \N__19568\
        );

    \I__4360\ : Glb2LocalMux
    port map (
            O => \N__19728\,
            I => \N__19568\
        );

    \I__4359\ : Glb2LocalMux
    port map (
            O => \N__19725\,
            I => \N__19568\
        );

    \I__4358\ : Glb2LocalMux
    port map (
            O => \N__19722\,
            I => \N__19568\
        );

    \I__4357\ : Glb2LocalMux
    port map (
            O => \N__19719\,
            I => \N__19568\
        );

    \I__4356\ : Glb2LocalMux
    port map (
            O => \N__19716\,
            I => \N__19568\
        );

    \I__4355\ : Glb2LocalMux
    port map (
            O => \N__19713\,
            I => \N__19568\
        );

    \I__4354\ : CEMux
    port map (
            O => \N__19712\,
            I => \N__19568\
        );

    \I__4353\ : Glb2LocalMux
    port map (
            O => \N__19709\,
            I => \N__19568\
        );

    \I__4352\ : Glb2LocalMux
    port map (
            O => \N__19706\,
            I => \N__19568\
        );

    \I__4351\ : Glb2LocalMux
    port map (
            O => \N__19703\,
            I => \N__19568\
        );

    \I__4350\ : Glb2LocalMux
    port map (
            O => \N__19700\,
            I => \N__19568\
        );

    \I__4349\ : Glb2LocalMux
    port map (
            O => \N__19697\,
            I => \N__19568\
        );

    \I__4348\ : Glb2LocalMux
    port map (
            O => \N__19694\,
            I => \N__19568\
        );

    \I__4347\ : Glb2LocalMux
    port map (
            O => \N__19691\,
            I => \N__19568\
        );

    \I__4346\ : Glb2LocalMux
    port map (
            O => \N__19688\,
            I => \N__19568\
        );

    \I__4345\ : Glb2LocalMux
    port map (
            O => \N__19685\,
            I => \N__19568\
        );

    \I__4344\ : GlobalMux
    port map (
            O => \N__19568\,
            I => \N__19565\
        );

    \I__4343\ : gio2CtrlBuf
    port map (
            O => \N__19565\,
            I => \N_65_g\
        );

    \I__4342\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19559\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__19559\,
            I => \N__19556\
        );

    \I__4340\ : Span4Mux_v
    port map (
            O => \N__19556\,
            I => \N__19552\
        );

    \I__4339\ : InMux
    port map (
            O => \N__19555\,
            I => \N__19549\
        );

    \I__4338\ : Span4Mux_v
    port map (
            O => \N__19552\,
            I => \N__19546\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__19549\,
            I => \N__19543\
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__19546\,
            I => vddq_ok
        );

    \I__4335\ : Odrv12
    port map (
            O => \N__19543\,
            I => vddq_ok
        );

    \I__4334\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19535\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__19535\,
            I => v5s_ok
        );

    \I__4332\ : InMux
    port map (
            O => \N__19532\,
            I => \N__19529\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__19529\,
            I => \N__19526\
        );

    \I__4330\ : Span4Mux_s3_h
    port map (
            O => \N__19526\,
            I => \N__19520\
        );

    \I__4329\ : InMux
    port map (
            O => \N__19525\,
            I => \N__19515\
        );

    \I__4328\ : InMux
    port map (
            O => \N__19524\,
            I => \N__19515\
        );

    \I__4327\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19512\
        );

    \I__4326\ : Sp12to4
    port map (
            O => \N__19520\,
            I => \N__19507\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__19515\,
            I => \N__19507\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__19512\,
            I => \N__19504\
        );

    \I__4323\ : Odrv12
    port map (
            O => \N__19507\,
            I => rsmrst_pwrgd_signal
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__19504\,
            I => rsmrst_pwrgd_signal
        );

    \I__4321\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__19496\,
            I => \N__19493\
        );

    \I__4319\ : Span4Mux_v
    port map (
            O => \N__19493\,
            I => \N__19490\
        );

    \I__4318\ : Odrv4
    port map (
            O => \N__19490\,
            I => vccst_cpu_ok
        );

    \I__4317\ : CascadeMux
    port map (
            O => \N__19487\,
            I => \ALL_SYS_PWRGD.m4_0_0_a2_1_cascade_\
        );

    \I__4316\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19481\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__19481\,
            I => \N__19478\
        );

    \I__4314\ : Span12Mux_v
    port map (
            O => \N__19478\,
            I => \N__19475\
        );

    \I__4313\ : Odrv12
    port map (
            O => \N__19475\,
            I => v33s_ok
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__19472\,
            I => \N__19467\
        );

    \I__4311\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19460\
        );

    \I__4310\ : InMux
    port map (
            O => \N__19470\,
            I => \N__19460\
        );

    \I__4309\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19453\
        );

    \I__4308\ : InMux
    port map (
            O => \N__19466\,
            I => \N__19453\
        );

    \I__4307\ : InMux
    port map (
            O => \N__19465\,
            I => \N__19453\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__19460\,
            I => \ALL_SYS_PWRGD.N_245\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__19453\,
            I => \ALL_SYS_PWRGD.N_245\
        );

    \I__4304\ : InMux
    port map (
            O => \N__19448\,
            I => \bfn_11_6_0_\
        );

    \I__4303\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19436\
        );

    \I__4302\ : InMux
    port map (
            O => \N__19444\,
            I => \N__19436\
        );

    \I__4301\ : InMux
    port map (
            O => \N__19443\,
            I => \N__19436\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__19436\,
            I => \N__19427\
        );

    \I__4299\ : InMux
    port map (
            O => \N__19435\,
            I => \N__19418\
        );

    \I__4298\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19418\
        );

    \I__4297\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19418\
        );

    \I__4296\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19418\
        );

    \I__4295\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19413\
        );

    \I__4294\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19413\
        );

    \I__4293\ : Span4Mux_s1_v
    port map (
            O => \N__19427\,
            I => \N__19410\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__19418\,
            I => \N__19407\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__19413\,
            I => \N__19404\
        );

    \I__4290\ : Span4Mux_h
    port map (
            O => \N__19410\,
            I => \N__19401\
        );

    \I__4289\ : Span4Mux_v
    port map (
            O => \N__19407\,
            I => \N__19398\
        );

    \I__4288\ : Span4Mux_h
    port map (
            O => \N__19404\,
            I => \N__19395\
        );

    \I__4287\ : Odrv4
    port map (
            O => \N__19401\,
            I => \COUNTER.un4_counter_7_THRU_CO\
        );

    \I__4286\ : Odrv4
    port map (
            O => \N__19398\,
            I => \COUNTER.un4_counter_7_THRU_CO\
        );

    \I__4285\ : Odrv4
    port map (
            O => \N__19395\,
            I => \COUNTER.un4_counter_7_THRU_CO\
        );

    \I__4284\ : CascadeMux
    port map (
            O => \N__19388\,
            I => \ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa_cascade_\
        );

    \I__4283\ : InMux
    port map (
            O => \N__19385\,
            I => \N__19381\
        );

    \I__4282\ : CascadeMux
    port map (
            O => \N__19384\,
            I => \N__19378\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__19381\,
            I => \N__19375\
        );

    \I__4280\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19372\
        );

    \I__4279\ : Span4Mux_v
    port map (
            O => \N__19375\,
            I => \N__19367\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__19372\,
            I => \N__19367\
        );

    \I__4277\ : Span4Mux_h
    port map (
            O => \N__19367\,
            I => \N__19364\
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__19364\,
            I => \ALL_SYS_PWRGD.un1_curr_state10_0\
        );

    \I__4275\ : CascadeMux
    port map (
            O => \N__19361\,
            I => \N__19357\
        );

    \I__4274\ : InMux
    port map (
            O => \N__19360\,
            I => \N__19353\
        );

    \I__4273\ : InMux
    port map (
            O => \N__19357\,
            I => \N__19348\
        );

    \I__4272\ : InMux
    port map (
            O => \N__19356\,
            I => \N__19348\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__19353\,
            I => \N__19343\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__19348\,
            I => \N__19343\
        );

    \I__4269\ : Span4Mux_v
    port map (
            O => \N__19343\,
            I => \N__19340\
        );

    \I__4268\ : Odrv4
    port map (
            O => \N__19340\,
            I => \ALL_SYS_PWRGD.N_1_i\
        );

    \I__4267\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19334\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__19334\,
            I => \N__19331\
        );

    \I__4265\ : Odrv4
    port map (
            O => \N__19331\,
            I => \ALL_SYS_PWRGD.N_36\
        );

    \I__4264\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19310\
        );

    \I__4263\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19310\
        );

    \I__4262\ : InMux
    port map (
            O => \N__19326\,
            I => \N__19310\
        );

    \I__4261\ : InMux
    port map (
            O => \N__19325\,
            I => \N__19310\
        );

    \I__4260\ : InMux
    port map (
            O => \N__19324\,
            I => \N__19310\
        );

    \I__4259\ : InMux
    port map (
            O => \N__19323\,
            I => \N__19310\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__19310\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_0\
        );

    \I__4257\ : InMux
    port map (
            O => \N__19307\,
            I => \N__19289\
        );

    \I__4256\ : InMux
    port map (
            O => \N__19306\,
            I => \N__19289\
        );

    \I__4255\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19289\
        );

    \I__4254\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19289\
        );

    \I__4253\ : InMux
    port map (
            O => \N__19303\,
            I => \N__19289\
        );

    \I__4252\ : InMux
    port map (
            O => \N__19302\,
            I => \N__19289\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__19289\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_1\
        );

    \I__4250\ : CascadeMux
    port map (
            O => \N__19286\,
            I => \N__19280\
        );

    \I__4249\ : IoInMux
    port map (
            O => \N__19285\,
            I => \N__19277\
        );

    \I__4248\ : IoInMux
    port map (
            O => \N__19284\,
            I => \N__19274\
        );

    \I__4247\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19269\
        );

    \I__4246\ : InMux
    port map (
            O => \N__19280\,
            I => \N__19269\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__19277\,
            I => \N__19266\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__19274\,
            I => \N__19263\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__19269\,
            I => \N__19260\
        );

    \I__4242\ : Span4Mux_s2_v
    port map (
            O => \N__19266\,
            I => \N__19257\
        );

    \I__4241\ : Span4Mux_s1_v
    port map (
            O => \N__19263\,
            I => \N__19254\
        );

    \I__4240\ : Span4Mux_s2_h
    port map (
            O => \N__19260\,
            I => \N__19251\
        );

    \I__4239\ : Span4Mux_v
    port map (
            O => \N__19257\,
            I => \N__19248\
        );

    \I__4238\ : Span4Mux_v
    port map (
            O => \N__19254\,
            I => \N__19245\
        );

    \I__4237\ : Span4Mux_h
    port map (
            O => \N__19251\,
            I => \N__19242\
        );

    \I__4236\ : Span4Mux_h
    port map (
            O => \N__19248\,
            I => \N__19237\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__19245\,
            I => \N__19237\
        );

    \I__4234\ : Span4Mux_h
    port map (
            O => \N__19242\,
            I => \N__19234\
        );

    \I__4233\ : Odrv4
    port map (
            O => \N__19237\,
            I => vccst_pwrgd
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__19234\,
            I => vccst_pwrgd
        );

    \I__4231\ : InMux
    port map (
            O => \N__19229\,
            I => \N__19223\
        );

    \I__4230\ : CascadeMux
    port map (
            O => \N__19228\,
            I => \N__19220\
        );

    \I__4229\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19215\
        );

    \I__4228\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19215\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__19223\,
            I => \N__19212\
        );

    \I__4226\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19209\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__19215\,
            I => \N__19206\
        );

    \I__4224\ : Span4Mux_h
    port map (
            O => \N__19212\,
            I => \N__19203\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__19209\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__4222\ : Odrv4
    port map (
            O => \N__19206\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__4221\ : Odrv4
    port map (
            O => \N__19203\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__4220\ : InMux
    port map (
            O => \N__19196\,
            I => \N__19190\
        );

    \I__4219\ : InMux
    port map (
            O => \N__19195\,
            I => \N__19190\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__4217\ : Span4Mux_v
    port map (
            O => \N__19187\,
            I => \N__19183\
        );

    \I__4216\ : InMux
    port map (
            O => \N__19186\,
            I => \N__19180\
        );

    \I__4215\ : Odrv4
    port map (
            O => \N__19183\,
            I => \RSMRST_PWRGD.N_241\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__19180\,
            I => \RSMRST_PWRGD.N_241\
        );

    \I__4213\ : InMux
    port map (
            O => \N__19175\,
            I => \N__19172\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__19172\,
            I => \N__19169\
        );

    \I__4211\ : Odrv4
    port map (
            O => \N__19169\,
            I => \COUNTER.un4_counter_0_and\
        );

    \I__4210\ : InMux
    port map (
            O => \N__19166\,
            I => \N__19163\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__19163\,
            I => \N__19160\
        );

    \I__4208\ : Span4Mux_v
    port map (
            O => \N__19160\,
            I => \N__19157\
        );

    \I__4207\ : Odrv4
    port map (
            O => \N__19157\,
            I => \COUNTER.un4_counter_1_and\
        );

    \I__4206\ : InMux
    port map (
            O => \N__19154\,
            I => \N__19151\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__19151\,
            I => \N__19148\
        );

    \I__4204\ : Odrv4
    port map (
            O => \N__19148\,
            I => \COUNTER.un4_counter_2_and\
        );

    \I__4203\ : InMux
    port map (
            O => \N__19145\,
            I => \N__19142\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__19142\,
            I => \N__19139\
        );

    \I__4201\ : Odrv12
    port map (
            O => \N__19139\,
            I => \COUNTER.un4_counter_3_and\
        );

    \I__4200\ : InMux
    port map (
            O => \N__19136\,
            I => \N__19133\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__19133\,
            I => \N__19130\
        );

    \I__4198\ : Odrv4
    port map (
            O => \N__19130\,
            I => \COUNTER.un4_counter_4_and\
        );

    \I__4197\ : InMux
    port map (
            O => \N__19127\,
            I => \N__19124\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__19124\,
            I => \N__19121\
        );

    \I__4195\ : Span4Mux_s2_h
    port map (
            O => \N__19121\,
            I => \N__19118\
        );

    \I__4194\ : Odrv4
    port map (
            O => \N__19118\,
            I => \COUNTER.un4_counter_5_and\
        );

    \I__4193\ : InMux
    port map (
            O => \N__19115\,
            I => \N__19112\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__19112\,
            I => \N__19109\
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__19109\,
            I => \COUNTER.un4_counter_6_and\
        );

    \I__4190\ : InMux
    port map (
            O => \N__19106\,
            I => \N__19103\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__19103\,
            I => \N__19100\
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__19100\,
            I => \COUNTER.un4_counter_7_and\
        );

    \I__4187\ : InMux
    port map (
            O => \N__19097\,
            I => \N__19093\
        );

    \I__4186\ : InMux
    port map (
            O => \N__19096\,
            I => \N__19090\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__19093\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__19090\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__19085\,
            I => \N__19081\
        );

    \I__4182\ : InMux
    port map (
            O => \N__19084\,
            I => \N__19078\
        );

    \I__4181\ : InMux
    port map (
            O => \N__19081\,
            I => \N__19075\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__19078\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__19075\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__4178\ : InMux
    port map (
            O => \N__19070\,
            I => \N__19066\
        );

    \I__4177\ : InMux
    port map (
            O => \N__19069\,
            I => \N__19063\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__19066\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__19063\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__4174\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19054\
        );

    \I__4173\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19051\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__19054\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__19051\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__4170\ : InMux
    port map (
            O => \N__19046\,
            I => \N__19042\
        );

    \I__4169\ : InMux
    port map (
            O => \N__19045\,
            I => \N__19039\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__19042\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__19039\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__4166\ : CascadeMux
    port map (
            O => \N__19034\,
            I => \N__19030\
        );

    \I__4165\ : InMux
    port map (
            O => \N__19033\,
            I => \N__19027\
        );

    \I__4164\ : InMux
    port map (
            O => \N__19030\,
            I => \N__19024\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__19027\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__19024\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__4161\ : InMux
    port map (
            O => \N__19019\,
            I => \N__19015\
        );

    \I__4160\ : InMux
    port map (
            O => \N__19018\,
            I => \N__19012\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__19015\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__19012\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__4157\ : InMux
    port map (
            O => \N__19007\,
            I => \N__19003\
        );

    \I__4156\ : InMux
    port map (
            O => \N__19006\,
            I => \N__19000\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__19003\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__19000\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__4153\ : InMux
    port map (
            O => \N__18995\,
            I => \N__18991\
        );

    \I__4152\ : InMux
    port map (
            O => \N__18994\,
            I => \N__18988\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__18991\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__18988\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__18983\,
            I => \N__18979\
        );

    \I__4148\ : InMux
    port map (
            O => \N__18982\,
            I => \N__18976\
        );

    \I__4147\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18973\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__18976\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__18973\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__4144\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18964\
        );

    \I__4143\ : InMux
    port map (
            O => \N__18967\,
            I => \N__18961\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__18964\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__18961\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__4140\ : InMux
    port map (
            O => \N__18956\,
            I => \N__18952\
        );

    \I__4139\ : InMux
    port map (
            O => \N__18955\,
            I => \N__18949\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__18952\,
            I => \N__18946\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__18949\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__18946\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__4135\ : InMux
    port map (
            O => \N__18941\,
            I => \N__18937\
        );

    \I__4134\ : InMux
    port map (
            O => \N__18940\,
            I => \N__18934\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__18937\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__18934\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__4131\ : CascadeMux
    port map (
            O => \N__18929\,
            I => \N__18925\
        );

    \I__4130\ : InMux
    port map (
            O => \N__18928\,
            I => \N__18922\
        );

    \I__4129\ : InMux
    port map (
            O => \N__18925\,
            I => \N__18919\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__18922\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__18919\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__4126\ : InMux
    port map (
            O => \N__18914\,
            I => \N__18910\
        );

    \I__4125\ : InMux
    port map (
            O => \N__18913\,
            I => \N__18907\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__18910\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__18907\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__4122\ : InMux
    port map (
            O => \N__18902\,
            I => \N__18899\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__18899\,
            I => \VPP_VDDQ.un6_count_11\
        );

    \I__4120\ : InMux
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__18893\,
            I => \VPP_VDDQ.un6_count_10\
        );

    \I__4118\ : CascadeMux
    port map (
            O => \N__18890\,
            I => \VPP_VDDQ.un6_count_9_cascade_\
        );

    \I__4117\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__18884\,
            I => \VPP_VDDQ.un6_count_8\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__18881\,
            I => \N__18878\
        );

    \I__4114\ : InMux
    port map (
            O => \N__18878\,
            I => \N__18874\
        );

    \I__4113\ : InMux
    port map (
            O => \N__18877\,
            I => \N__18871\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__18874\,
            I => \N__18868\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__18871\,
            I => \N__18865\
        );

    \I__4110\ : Odrv4
    port map (
            O => \N__18868\,
            I => \VPP_VDDQ.count_esr_RNIRFM64Z0Z_15\
        );

    \I__4109\ : Odrv4
    port map (
            O => \N__18865\,
            I => \VPP_VDDQ.count_esr_RNIRFM64Z0Z_15\
        );

    \I__4108\ : InMux
    port map (
            O => \N__18860\,
            I => \N__18856\
        );

    \I__4107\ : InMux
    port map (
            O => \N__18859\,
            I => \N__18853\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__18856\,
            I => \N__18850\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__18853\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__4104\ : Odrv4
    port map (
            O => \N__18850\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__4103\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18841\
        );

    \I__4102\ : InMux
    port map (
            O => \N__18844\,
            I => \N__18838\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__18841\,
            I => \N__18835\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__18838\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__4099\ : Odrv4
    port map (
            O => \N__18835\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__4098\ : CascadeMux
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__4097\ : InMux
    port map (
            O => \N__18827\,
            I => \N__18823\
        );

    \I__4096\ : InMux
    port map (
            O => \N__18826\,
            I => \N__18820\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__18823\,
            I => \N__18817\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__18820\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__4093\ : Odrv12
    port map (
            O => \N__18817\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__4092\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18808\
        );

    \I__4091\ : InMux
    port map (
            O => \N__18811\,
            I => \N__18805\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__18808\,
            I => \N__18802\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__18805\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__4088\ : Odrv4
    port map (
            O => \N__18802\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__4087\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18793\
        );

    \I__4086\ : InMux
    port map (
            O => \N__18796\,
            I => \N__18790\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__18793\,
            I => \N__18787\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__18790\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__18787\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__4082\ : InMux
    port map (
            O => \N__18782\,
            I => \N__18778\
        );

    \I__4081\ : InMux
    port map (
            O => \N__18781\,
            I => \N__18775\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__18778\,
            I => \N__18772\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__18775\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__4078\ : Odrv4
    port map (
            O => \N__18772\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__18767\,
            I => \N__18763\
        );

    \I__4076\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18760\
        );

    \I__4075\ : InMux
    port map (
            O => \N__18763\,
            I => \N__18757\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__18760\,
            I => \N__18752\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__18757\,
            I => \N__18752\
        );

    \I__4072\ : Odrv4
    port map (
            O => \N__18752\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__4071\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18746\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__18746\,
            I => \N__18742\
        );

    \I__4069\ : InMux
    port map (
            O => \N__18745\,
            I => \N__18739\
        );

    \I__4068\ : Span4Mux_s2_h
    port map (
            O => \N__18742\,
            I => \N__18736\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__18739\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__18736\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__4065\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18728\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__18728\,
            I => \N__18724\
        );

    \I__4063\ : InMux
    port map (
            O => \N__18727\,
            I => \N__18721\
        );

    \I__4062\ : Span4Mux_s2_h
    port map (
            O => \N__18724\,
            I => \N__18718\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__18721\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__4060\ : Odrv4
    port map (
            O => \N__18718\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__4059\ : InMux
    port map (
            O => \N__18713\,
            I => \N__18710\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__18710\,
            I => \N__18706\
        );

    \I__4057\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18703\
        );

    \I__4056\ : Span4Mux_s2_h
    port map (
            O => \N__18706\,
            I => \N__18700\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__18703\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__18700\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__18695\,
            I => \N__18692\
        );

    \I__4052\ : InMux
    port map (
            O => \N__18692\,
            I => \N__18689\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__18689\,
            I => \N__18685\
        );

    \I__4050\ : InMux
    port map (
            O => \N__18688\,
            I => \N__18682\
        );

    \I__4049\ : Span4Mux_s2_h
    port map (
            O => \N__18685\,
            I => \N__18679\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__18682\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__18679\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__4046\ : InMux
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__18671\,
            I => \N__18667\
        );

    \I__4044\ : InMux
    port map (
            O => \N__18670\,
            I => \N__18664\
        );

    \I__4043\ : Span4Mux_s2_h
    port map (
            O => \N__18667\,
            I => \N__18661\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__18664\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__4041\ : Odrv4
    port map (
            O => \N__18661\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__4040\ : InMux
    port map (
            O => \N__18656\,
            I => \N__18653\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__18653\,
            I => \RSMRST_PWRGD.m4_i_i_a2_0_11\
        );

    \I__4038\ : CascadeMux
    port map (
            O => \N__18650\,
            I => \RSMRST_PWRGD.m4_i_i_a2_0_9_cascade_\
        );

    \I__4037\ : InMux
    port map (
            O => \N__18647\,
            I => \N__18643\
        );

    \I__4036\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18640\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__18643\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__18640\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__4033\ : InMux
    port map (
            O => \N__18635\,
            I => \N__18631\
        );

    \I__4032\ : InMux
    port map (
            O => \N__18634\,
            I => \N__18628\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__18631\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__18628\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__4029\ : InMux
    port map (
            O => \N__18623\,
            I => \N__18619\
        );

    \I__4028\ : InMux
    port map (
            O => \N__18622\,
            I => \N__18616\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__18619\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__18616\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__18611\,
            I => \RSMRST_PWRGD.m4_i_i_a2_0_7_cascade_\
        );

    \I__4024\ : InMux
    port map (
            O => \N__18608\,
            I => \N__18604\
        );

    \I__4023\ : InMux
    port map (
            O => \N__18607\,
            I => \N__18601\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__18604\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__18601\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__4020\ : InMux
    port map (
            O => \N__18596\,
            I => \N__18593\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__18593\,
            I => \RSMRST_PWRGD.m4_i_i_a2_0_12\
        );

    \I__4018\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18586\
        );

    \I__4017\ : InMux
    port map (
            O => \N__18589\,
            I => \N__18583\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__18586\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__18583\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__4014\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18574\
        );

    \I__4013\ : InMux
    port map (
            O => \N__18577\,
            I => \N__18571\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__18574\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__18571\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__18566\,
            I => \N__18562\
        );

    \I__4009\ : InMux
    port map (
            O => \N__18565\,
            I => \N__18559\
        );

    \I__4008\ : InMux
    port map (
            O => \N__18562\,
            I => \N__18556\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__18559\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__18556\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__4005\ : InMux
    port map (
            O => \N__18551\,
            I => \N__18547\
        );

    \I__4004\ : InMux
    port map (
            O => \N__18550\,
            I => \N__18544\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__18547\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__18544\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__4001\ : InMux
    port map (
            O => \N__18539\,
            I => \N__18536\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__18536\,
            I => \RSMRST_PWRGD.m4_i_i_a2_0_10\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__18533\,
            I => \RSMRST_PWRGD.N_240_cascade_\
        );

    \I__3998\ : SRMux
    port map (
            O => \N__18530\,
            I => \N__18526\
        );

    \I__3997\ : SRMux
    port map (
            O => \N__18529\,
            I => \N__18523\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__18526\,
            I => \N__18519\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__18523\,
            I => \N__18516\
        );

    \I__3994\ : SRMux
    port map (
            O => \N__18522\,
            I => \N__18513\
        );

    \I__3993\ : Span4Mux_v
    port map (
            O => \N__18519\,
            I => \N__18506\
        );

    \I__3992\ : Span4Mux_v
    port map (
            O => \N__18516\,
            I => \N__18506\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__18513\,
            I => \N__18506\
        );

    \I__3990\ : Sp12to4
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__3989\ : Odrv12
    port map (
            O => \N__18503\,
            I => \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__18500\,
            I => \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0_cascade_\
        );

    \I__3987\ : CEMux
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__18494\,
            I => \RSMRST_PWRGD.N_65_2\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__18491\,
            I => \N__18487\
        );

    \I__3984\ : InMux
    port map (
            O => \N__18490\,
            I => \N__18484\
        );

    \I__3983\ : InMux
    port map (
            O => \N__18487\,
            I => \N__18481\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__18484\,
            I => \N__18476\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__18481\,
            I => \N__18476\
        );

    \I__3980\ : Span4Mux_h
    port map (
            O => \N__18476\,
            I => \N__18473\
        );

    \I__3979\ : Odrv4
    port map (
            O => \N__18473\,
            I => \RSMRST_PWRGD.N_37\
        );

    \I__3978\ : InMux
    port map (
            O => \N__18470\,
            I => \N__18466\
        );

    \I__3977\ : InMux
    port map (
            O => \N__18469\,
            I => \N__18463\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__18466\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__18463\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__3974\ : InMux
    port map (
            O => \N__18458\,
            I => \N__18454\
        );

    \I__3973\ : InMux
    port map (
            O => \N__18457\,
            I => \N__18451\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__18454\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__18451\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__3970\ : InMux
    port map (
            O => \N__18446\,
            I => \POWERLED.un1_count_clk_1_cry_10\
        );

    \I__3969\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18439\
        );

    \I__3968\ : InMux
    port map (
            O => \N__18442\,
            I => \N__18436\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__18439\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__18436\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__3965\ : InMux
    port map (
            O => \N__18431\,
            I => \POWERLED.un1_count_clk_1_cry_11\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__18428\,
            I => \N__18424\
        );

    \I__3963\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18421\
        );

    \I__3962\ : InMux
    port map (
            O => \N__18424\,
            I => \N__18418\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__18421\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__18418\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__3959\ : InMux
    port map (
            O => \N__18413\,
            I => \POWERLED.un1_count_clk_1_cry_12\
        );

    \I__3958\ : InMux
    port map (
            O => \N__18410\,
            I => \N__18406\
        );

    \I__3957\ : InMux
    port map (
            O => \N__18409\,
            I => \N__18403\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__18406\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__18403\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__3954\ : InMux
    port map (
            O => \N__18398\,
            I => \POWERLED.un1_count_clk_1_cry_13\
        );

    \I__3953\ : InMux
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__18392\,
            I => \N__18389\
        );

    \I__3951\ : Span4Mux_v
    port map (
            O => \N__18389\,
            I => \N__18384\
        );

    \I__3950\ : InMux
    port map (
            O => \N__18388\,
            I => \N__18381\
        );

    \I__3949\ : InMux
    port map (
            O => \N__18387\,
            I => \N__18378\
        );

    \I__3948\ : IoSpan4Mux
    port map (
            O => \N__18384\,
            I => \N__18371\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__18381\,
            I => \N__18366\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__18378\,
            I => \N__18366\
        );

    \I__3945\ : InMux
    port map (
            O => \N__18377\,
            I => \N__18363\
        );

    \I__3944\ : InMux
    port map (
            O => \N__18376\,
            I => \N__18360\
        );

    \I__3943\ : InMux
    port map (
            O => \N__18375\,
            I => \N__18357\
        );

    \I__3942\ : IoInMux
    port map (
            O => \N__18374\,
            I => \N__18353\
        );

    \I__3941\ : Span4Mux_s3_h
    port map (
            O => \N__18371\,
            I => \N__18344\
        );

    \I__3940\ : Span4Mux_v
    port map (
            O => \N__18366\,
            I => \N__18344\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__18363\,
            I => \N__18344\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__18360\,
            I => \N__18344\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__18357\,
            I => \N__18341\
        );

    \I__3936\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18338\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__18353\,
            I => \N__18333\
        );

    \I__3934\ : Span4Mux_h
    port map (
            O => \N__18344\,
            I => \N__18328\
        );

    \I__3933\ : Span4Mux_v
    port map (
            O => \N__18341\,
            I => \N__18328\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__18338\,
            I => \N__18325\
        );

    \I__3931\ : InMux
    port map (
            O => \N__18337\,
            I => \N__18322\
        );

    \I__3930\ : InMux
    port map (
            O => \N__18336\,
            I => \N__18319\
        );

    \I__3929\ : Span4Mux_s3_h
    port map (
            O => \N__18333\,
            I => \N__18315\
        );

    \I__3928\ : Span4Mux_v
    port map (
            O => \N__18328\,
            I => \N__18308\
        );

    \I__3927\ : Span4Mux_h
    port map (
            O => \N__18325\,
            I => \N__18308\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__18322\,
            I => \N__18308\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__18319\,
            I => \N__18305\
        );

    \I__3924\ : CascadeMux
    port map (
            O => \N__18318\,
            I => \N__18302\
        );

    \I__3923\ : Span4Mux_v
    port map (
            O => \N__18315\,
            I => \N__18294\
        );

    \I__3922\ : Span4Mux_v
    port map (
            O => \N__18308\,
            I => \N__18294\
        );

    \I__3921\ : Span4Mux_s2_v
    port map (
            O => \N__18305\,
            I => \N__18294\
        );

    \I__3920\ : InMux
    port map (
            O => \N__18302\,
            I => \N__18289\
        );

    \I__3919\ : InMux
    port map (
            O => \N__18301\,
            I => \N__18289\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__18294\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__18289\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3916\ : InMux
    port map (
            O => \N__18284\,
            I => \bfn_9_11_0_\
        );

    \I__3915\ : CascadeMux
    port map (
            O => \N__18281\,
            I => \N__18277\
        );

    \I__3914\ : InMux
    port map (
            O => \N__18280\,
            I => \N__18274\
        );

    \I__3913\ : InMux
    port map (
            O => \N__18277\,
            I => \N__18271\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__18274\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__18271\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__3910\ : CEMux
    port map (
            O => \N__18266\,
            I => \N__18263\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__18263\,
            I => \N__18260\
        );

    \I__3908\ : Span4Mux_v
    port map (
            O => \N__18260\,
            I => \N__18257\
        );

    \I__3907\ : Span4Mux_s2_h
    port map (
            O => \N__18257\,
            I => \N__18254\
        );

    \I__3906\ : Odrv4
    port map (
            O => \N__18254\,
            I => \POWERLED.N_65_0\
        );

    \I__3905\ : SRMux
    port map (
            O => \N__18251\,
            I => \N__18247\
        );

    \I__3904\ : SRMux
    port map (
            O => \N__18250\,
            I => \N__18244\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__18247\,
            I => \N__18240\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__18244\,
            I => \N__18237\
        );

    \I__3901\ : SRMux
    port map (
            O => \N__18243\,
            I => \N__18234\
        );

    \I__3900\ : Span4Mux_v
    port map (
            O => \N__18240\,
            I => \N__18226\
        );

    \I__3899\ : Span4Mux_v
    port map (
            O => \N__18237\,
            I => \N__18226\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__18234\,
            I => \N__18226\
        );

    \I__3897\ : InMux
    port map (
            O => \N__18233\,
            I => \N__18223\
        );

    \I__3896\ : Odrv4
    port map (
            O => \N__18226\,
            I => \POWERLED.count_clk_RNIOH1J11Z0Z_7\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__18223\,
            I => \POWERLED.count_clk_RNIOH1J11Z0Z_7\
        );

    \I__3894\ : InMux
    port map (
            O => \N__18218\,
            I => \N__18214\
        );

    \I__3893\ : InMux
    port map (
            O => \N__18217\,
            I => \N__18211\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__18214\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__18211\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__3890\ : InMux
    port map (
            O => \N__18206\,
            I => \N__18202\
        );

    \I__3889\ : InMux
    port map (
            O => \N__18205\,
            I => \N__18199\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__18202\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__18199\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__18194\,
            I => \N__18190\
        );

    \I__3885\ : InMux
    port map (
            O => \N__18193\,
            I => \N__18187\
        );

    \I__3884\ : InMux
    port map (
            O => \N__18190\,
            I => \N__18184\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__18187\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__18184\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__3881\ : InMux
    port map (
            O => \N__18179\,
            I => \N__18175\
        );

    \I__3880\ : InMux
    port map (
            O => \N__18178\,
            I => \N__18172\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__18175\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__18172\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__3877\ : InMux
    port map (
            O => \N__18167\,
            I => \N__18163\
        );

    \I__3876\ : InMux
    port map (
            O => \N__18166\,
            I => \N__18160\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__18163\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__18160\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__3873\ : InMux
    port map (
            O => \N__18155\,
            I => \N__18151\
        );

    \I__3872\ : InMux
    port map (
            O => \N__18154\,
            I => \N__18148\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__18151\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__18148\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__3869\ : CascadeMux
    port map (
            O => \N__18143\,
            I => \N__18139\
        );

    \I__3868\ : InMux
    port map (
            O => \N__18142\,
            I => \N__18136\
        );

    \I__3867\ : InMux
    port map (
            O => \N__18139\,
            I => \N__18133\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__18136\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__18133\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__3864\ : InMux
    port map (
            O => \N__18128\,
            I => \N__18124\
        );

    \I__3863\ : InMux
    port map (
            O => \N__18127\,
            I => \N__18121\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__18124\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__18121\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__3860\ : InMux
    port map (
            O => \N__18116\,
            I => \N__18111\
        );

    \I__3859\ : InMux
    port map (
            O => \N__18115\,
            I => \N__18106\
        );

    \I__3858\ : InMux
    port map (
            O => \N__18114\,
            I => \N__18106\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__18111\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__18106\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__3855\ : InMux
    port map (
            O => \N__18101\,
            I => \POWERLED.un1_count_clk_1_cry_2\
        );

    \I__3854\ : InMux
    port map (
            O => \N__18098\,
            I => \N__18093\
        );

    \I__3853\ : InMux
    port map (
            O => \N__18097\,
            I => \N__18088\
        );

    \I__3852\ : InMux
    port map (
            O => \N__18096\,
            I => \N__18088\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__18093\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__18088\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__3849\ : InMux
    port map (
            O => \N__18083\,
            I => \POWERLED.un1_count_clk_1_cry_3\
        );

    \I__3848\ : InMux
    port map (
            O => \N__18080\,
            I => \N__18074\
        );

    \I__3847\ : InMux
    port map (
            O => \N__18079\,
            I => \N__18069\
        );

    \I__3846\ : InMux
    port map (
            O => \N__18078\,
            I => \N__18069\
        );

    \I__3845\ : InMux
    port map (
            O => \N__18077\,
            I => \N__18066\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__18074\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__18069\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__18066\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__3841\ : InMux
    port map (
            O => \N__18059\,
            I => \POWERLED.un1_count_clk_1_cry_4\
        );

    \I__3840\ : InMux
    port map (
            O => \N__18056\,
            I => \N__18052\
        );

    \I__3839\ : InMux
    port map (
            O => \N__18055\,
            I => \N__18048\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__18052\,
            I => \N__18045\
        );

    \I__3837\ : InMux
    port map (
            O => \N__18051\,
            I => \N__18041\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__18048\,
            I => \N__18038\
        );

    \I__3835\ : Span4Mux_h
    port map (
            O => \N__18045\,
            I => \N__18035\
        );

    \I__3834\ : InMux
    port map (
            O => \N__18044\,
            I => \N__18032\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__18041\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__3832\ : Odrv4
    port map (
            O => \N__18038\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__3831\ : Odrv4
    port map (
            O => \N__18035\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__18032\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__3829\ : InMux
    port map (
            O => \N__18023\,
            I => \POWERLED.un1_count_clk_1_cry_5\
        );

    \I__3828\ : InMux
    port map (
            O => \N__18020\,
            I => \N__18013\
        );

    \I__3827\ : InMux
    port map (
            O => \N__18019\,
            I => \N__18008\
        );

    \I__3826\ : InMux
    port map (
            O => \N__18018\,
            I => \N__18008\
        );

    \I__3825\ : InMux
    port map (
            O => \N__18017\,
            I => \N__18001\
        );

    \I__3824\ : InMux
    port map (
            O => \N__18016\,
            I => \N__18001\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__18013\,
            I => \N__17997\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__18008\,
            I => \N__17994\
        );

    \I__3821\ : InMux
    port map (
            O => \N__18007\,
            I => \N__17991\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__18006\,
            I => \N__17987\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__18001\,
            I => \N__17984\
        );

    \I__3818\ : InMux
    port map (
            O => \N__18000\,
            I => \N__17981\
        );

    \I__3817\ : Span4Mux_h
    port map (
            O => \N__17997\,
            I => \N__17978\
        );

    \I__3816\ : Span12Mux_s7_v
    port map (
            O => \N__17994\,
            I => \N__17973\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__17991\,
            I => \N__17973\
        );

    \I__3814\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17968\
        );

    \I__3813\ : InMux
    port map (
            O => \N__17987\,
            I => \N__17968\
        );

    \I__3812\ : Span4Mux_h
    port map (
            O => \N__17984\,
            I => \N__17965\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__17981\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__17978\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__3809\ : Odrv12
    port map (
            O => \N__17973\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__17968\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__3807\ : Odrv4
    port map (
            O => \N__17965\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__3806\ : InMux
    port map (
            O => \N__17954\,
            I => \POWERLED.un1_count_clk_1_cry_6\
        );

    \I__3805\ : InMux
    port map (
            O => \N__17951\,
            I => \N__17946\
        );

    \I__3804\ : InMux
    port map (
            O => \N__17950\,
            I => \N__17941\
        );

    \I__3803\ : InMux
    port map (
            O => \N__17949\,
            I => \N__17941\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__17946\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__17941\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__3800\ : InMux
    port map (
            O => \N__17936\,
            I => \bfn_9_10_0_\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17933\,
            I => \N__17927\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17932\,
            I => \N__17920\
        );

    \I__3797\ : InMux
    port map (
            O => \N__17931\,
            I => \N__17920\
        );

    \I__3796\ : InMux
    port map (
            O => \N__17930\,
            I => \N__17920\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__17927\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__17920\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__3793\ : InMux
    port map (
            O => \N__17915\,
            I => \POWERLED.un1_count_clk_1_cry_8\
        );

    \I__3792\ : InMux
    port map (
            O => \N__17912\,
            I => \N__17908\
        );

    \I__3791\ : InMux
    port map (
            O => \N__17911\,
            I => \N__17905\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__17908\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__17905\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__3788\ : InMux
    port map (
            O => \N__17900\,
            I => \POWERLED.un1_count_clk_1_cry_9\
        );

    \I__3787\ : InMux
    port map (
            O => \N__17897\,
            I => \N__17894\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__17894\,
            I => \ALL_SYS_PWRGD.un4_count_9\
        );

    \I__3785\ : SRMux
    port map (
            O => \N__17891\,
            I => \N__17887\
        );

    \I__3784\ : SRMux
    port map (
            O => \N__17890\,
            I => \N__17884\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__17887\,
            I => \N__17880\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__17884\,
            I => \N__17877\
        );

    \I__3781\ : SRMux
    port map (
            O => \N__17883\,
            I => \N__17874\
        );

    \I__3780\ : Span4Mux_v
    port map (
            O => \N__17880\,
            I => \N__17867\
        );

    \I__3779\ : Span4Mux_v
    port map (
            O => \N__17877\,
            I => \N__17867\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__17874\,
            I => \N__17867\
        );

    \I__3777\ : Sp12to4
    port map (
            O => \N__17867\,
            I => \N__17864\
        );

    \I__3776\ : Odrv12
    port map (
            O => \N__17864\,
            I => \ALL_SYS_PWRGD.curr_state_RNIKNST6Z0Z_0\
        );

    \I__3775\ : CascadeMux
    port map (
            O => \N__17861\,
            I => \ALL_SYS_PWRGD.curr_state_RNIKNST6Z0Z_0_cascade_\
        );

    \I__3774\ : CEMux
    port map (
            O => \N__17858\,
            I => \N__17855\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__17855\,
            I => \ALL_SYS_PWRGD.N_65_4\
        );

    \I__3772\ : IoInMux
    port map (
            O => \N__17852\,
            I => \N__17849\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__17849\,
            I => \N__17845\
        );

    \I__3770\ : IoInMux
    port map (
            O => \N__17848\,
            I => \N__17842\
        );

    \I__3769\ : IoSpan4Mux
    port map (
            O => \N__17845\,
            I => \N__17838\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__17842\,
            I => \N__17835\
        );

    \I__3767\ : InMux
    port map (
            O => \N__17841\,
            I => \N__17832\
        );

    \I__3766\ : IoSpan4Mux
    port map (
            O => \N__17838\,
            I => \N__17829\
        );

    \I__3765\ : Span12Mux_s8_h
    port map (
            O => \N__17835\,
            I => \N__17824\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__17832\,
            I => \N__17824\
        );

    \I__3763\ : Odrv4
    port map (
            O => \N__17829\,
            I => slp_susn
        );

    \I__3762\ : Odrv12
    port map (
            O => \N__17824\,
            I => slp_susn
        );

    \I__3761\ : InMux
    port map (
            O => \N__17819\,
            I => \N__17816\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__17816\,
            I => \N__17813\
        );

    \I__3759\ : Span4Mux_v
    port map (
            O => \N__17813\,
            I => \N__17810\
        );

    \I__3758\ : Sp12to4
    port map (
            O => \N__17810\,
            I => \N__17807\
        );

    \I__3757\ : Odrv12
    port map (
            O => \N__17807\,
            I => v5a_ok
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__17804\,
            I => \N__17801\
        );

    \I__3755\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17798\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__17798\,
            I => \N__17795\
        );

    \I__3753\ : Span4Mux_h
    port map (
            O => \N__17795\,
            I => \N__17792\
        );

    \I__3752\ : Span4Mux_v
    port map (
            O => \N__17792\,
            I => \N__17789\
        );

    \I__3751\ : Span4Mux_v
    port map (
            O => \N__17789\,
            I => \N__17786\
        );

    \I__3750\ : Odrv4
    port map (
            O => \N__17786\,
            I => v33a_ok
        );

    \I__3749\ : IoInMux
    port map (
            O => \N__17783\,
            I => \N__17780\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__17780\,
            I => \N__17777\
        );

    \I__3747\ : IoSpan4Mux
    port map (
            O => \N__17777\,
            I => \N__17773\
        );

    \I__3746\ : InMux
    port map (
            O => \N__17776\,
            I => \N__17770\
        );

    \I__3745\ : IoSpan4Mux
    port map (
            O => \N__17773\,
            I => \N__17767\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__17770\,
            I => \N__17764\
        );

    \I__3743\ : Span4Mux_s3_h
    port map (
            O => \N__17767\,
            I => \N__17761\
        );

    \I__3742\ : Sp12to4
    port map (
            O => \N__17764\,
            I => \N__17758\
        );

    \I__3741\ : Sp12to4
    port map (
            O => \N__17761\,
            I => \N__17753\
        );

    \I__3740\ : Span12Mux_s11_v
    port map (
            O => \N__17758\,
            I => \N__17753\
        );

    \I__3739\ : Odrv12
    port map (
            O => \N__17753\,
            I => v1p8a_ok
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__17750\,
            I => \N__17747\
        );

    \I__3737\ : InMux
    port map (
            O => \N__17747\,
            I => \N__17741\
        );

    \I__3736\ : InMux
    port map (
            O => \N__17746\,
            I => \N__17741\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__17741\,
            I => \COUNTER.tmp_i\
        );

    \I__3734\ : InMux
    port map (
            O => \N__17738\,
            I => \N__17734\
        );

    \I__3733\ : IoInMux
    port map (
            O => \N__17737\,
            I => \N__17731\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__17734\,
            I => \N__17728\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__17731\,
            I => \N__17725\
        );

    \I__3730\ : Span4Mux_v
    port map (
            O => \N__17728\,
            I => \N__17722\
        );

    \I__3729\ : Span4Mux_s0_h
    port map (
            O => \N__17725\,
            I => \N__17719\
        );

    \I__3728\ : Span4Mux_h
    port map (
            O => \N__17722\,
            I => \N__17716\
        );

    \I__3727\ : Span4Mux_h
    port map (
            O => \N__17719\,
            I => \N__17713\
        );

    \I__3726\ : Span4Mux_v
    port map (
            O => \N__17716\,
            I => \N__17710\
        );

    \I__3725\ : Span4Mux_h
    port map (
            O => \N__17713\,
            I => \N__17707\
        );

    \I__3724\ : Odrv4
    port map (
            O => \N__17710\,
            I => \tmp_RNIRH3P\
        );

    \I__3723\ : Odrv4
    port map (
            O => \N__17707\,
            I => \tmp_RNIRH3P\
        );

    \I__3722\ : CascadeMux
    port map (
            O => \N__17702\,
            I => \N__17698\
        );

    \I__3721\ : InMux
    port map (
            O => \N__17701\,
            I => \N__17695\
        );

    \I__3720\ : InMux
    port map (
            O => \N__17698\,
            I => \N__17692\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__17695\,
            I => \N__17687\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__17692\,
            I => \N__17687\
        );

    \I__3717\ : Span4Mux_h
    port map (
            O => \N__17687\,
            I => \N__17684\
        );

    \I__3716\ : Odrv4
    port map (
            O => \N__17684\,
            I => \POWERLED.count_clk_1_sqmuxa_5_i\
        );

    \I__3715\ : InMux
    port map (
            O => \N__17681\,
            I => \N__17677\
        );

    \I__3714\ : InMux
    port map (
            O => \N__17680\,
            I => \N__17674\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__17677\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__17674\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__3711\ : InMux
    port map (
            O => \N__17669\,
            I => \N__17663\
        );

    \I__3710\ : InMux
    port map (
            O => \N__17668\,
            I => \N__17656\
        );

    \I__3709\ : InMux
    port map (
            O => \N__17667\,
            I => \N__17656\
        );

    \I__3708\ : InMux
    port map (
            O => \N__17666\,
            I => \N__17656\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__17663\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__17656\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__3705\ : InMux
    port map (
            O => \N__17651\,
            I => \POWERLED.un1_count_clk_1_cry_0\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__17648\,
            I => \N__17644\
        );

    \I__3703\ : InMux
    port map (
            O => \N__17647\,
            I => \N__17640\
        );

    \I__3702\ : InMux
    port map (
            O => \N__17644\,
            I => \N__17637\
        );

    \I__3701\ : InMux
    port map (
            O => \N__17643\,
            I => \N__17634\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__17640\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__17637\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__17634\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__3697\ : InMux
    port map (
            O => \N__17627\,
            I => \POWERLED.un1_count_clk_1_cry_1\
        );

    \I__3696\ : InMux
    port map (
            O => \N__17624\,
            I => \N__17621\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__17621\,
            I => \N__17618\
        );

    \I__3694\ : Span4Mux_v
    port map (
            O => \N__17618\,
            I => \N__17615\
        );

    \I__3693\ : Odrv4
    port map (
            O => \N__17615\,
            I => \COUNTER.counter_1_cry_3_THRU_CO\
        );

    \I__3692\ : InMux
    port map (
            O => \N__17612\,
            I => \N__17608\
        );

    \I__3691\ : CascadeMux
    port map (
            O => \N__17611\,
            I => \N__17604\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__17608\,
            I => \N__17601\
        );

    \I__3689\ : InMux
    port map (
            O => \N__17607\,
            I => \N__17596\
        );

    \I__3688\ : InMux
    port map (
            O => \N__17604\,
            I => \N__17596\
        );

    \I__3687\ : Odrv12
    port map (
            O => \N__17601\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__17596\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__3685\ : InMux
    port map (
            O => \N__17591\,
            I => \N__17587\
        );

    \I__3684\ : CascadeMux
    port map (
            O => \N__17590\,
            I => \N__17584\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__17587\,
            I => \N__17581\
        );

    \I__3682\ : InMux
    port map (
            O => \N__17584\,
            I => \N__17578\
        );

    \I__3681\ : Sp12to4
    port map (
            O => \N__17581\,
            I => \N__17571\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__17578\,
            I => \N__17571\
        );

    \I__3679\ : InMux
    port map (
            O => \N__17577\,
            I => \N__17566\
        );

    \I__3678\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17566\
        );

    \I__3677\ : Odrv12
    port map (
            O => \N__17571\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__17566\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3675\ : InMux
    port map (
            O => \N__17561\,
            I => \N__17558\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__17558\,
            I => \N__17555\
        );

    \I__3673\ : Odrv12
    port map (
            O => \N__17555\,
            I => \COUNTER.counter_1_cry_1_THRU_CO\
        );

    \I__3672\ : InMux
    port map (
            O => \N__17552\,
            I => \N__17549\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__17549\,
            I => \N__17546\
        );

    \I__3670\ : Span4Mux_s1_v
    port map (
            O => \N__17546\,
            I => \N__17541\
        );

    \I__3669\ : InMux
    port map (
            O => \N__17545\,
            I => \N__17536\
        );

    \I__3668\ : InMux
    port map (
            O => \N__17544\,
            I => \N__17536\
        );

    \I__3667\ : Odrv4
    port map (
            O => \N__17541\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__17536\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__3665\ : InMux
    port map (
            O => \N__17531\,
            I => \N__17528\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__17528\,
            I => \N__17525\
        );

    \I__3663\ : Odrv12
    port map (
            O => \N__17525\,
            I => \COUNTER.counter_1_cry_2_THRU_CO\
        );

    \I__3662\ : InMux
    port map (
            O => \N__17522\,
            I => \N__17518\
        );

    \I__3661\ : CascadeMux
    port map (
            O => \N__17521\,
            I => \N__17515\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__17518\,
            I => \N__17511\
        );

    \I__3659\ : InMux
    port map (
            O => \N__17515\,
            I => \N__17506\
        );

    \I__3658\ : InMux
    port map (
            O => \N__17514\,
            I => \N__17506\
        );

    \I__3657\ : Odrv12
    port map (
            O => \N__17511\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__17506\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__3655\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17497\
        );

    \I__3654\ : InMux
    port map (
            O => \N__17500\,
            I => \N__17494\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__17497\,
            I => \ALL_SYS_PWRGD.countZ0Z_7\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__17494\,
            I => \ALL_SYS_PWRGD.countZ0Z_7\
        );

    \I__3651\ : InMux
    port map (
            O => \N__17489\,
            I => \N__17485\
        );

    \I__3650\ : InMux
    port map (
            O => \N__17488\,
            I => \N__17482\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__17485\,
            I => \ALL_SYS_PWRGD.countZ0Z_8\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__17482\,
            I => \ALL_SYS_PWRGD.countZ0Z_8\
        );

    \I__3647\ : CascadeMux
    port map (
            O => \N__17477\,
            I => \N__17473\
        );

    \I__3646\ : InMux
    port map (
            O => \N__17476\,
            I => \N__17470\
        );

    \I__3645\ : InMux
    port map (
            O => \N__17473\,
            I => \N__17467\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__17470\,
            I => \ALL_SYS_PWRGD.countZ0Z_6\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__17467\,
            I => \ALL_SYS_PWRGD.countZ0Z_6\
        );

    \I__3642\ : InMux
    port map (
            O => \N__17462\,
            I => \N__17458\
        );

    \I__3641\ : InMux
    port map (
            O => \N__17461\,
            I => \N__17455\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__17458\,
            I => \ALL_SYS_PWRGD.countZ0Z_4\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__17455\,
            I => \ALL_SYS_PWRGD.countZ0Z_4\
        );

    \I__3638\ : InMux
    port map (
            O => \N__17450\,
            I => \N__17446\
        );

    \I__3637\ : InMux
    port map (
            O => \N__17449\,
            I => \N__17443\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__17446\,
            I => \ALL_SYS_PWRGD.countZ0Z_14\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__17443\,
            I => \ALL_SYS_PWRGD.countZ0Z_14\
        );

    \I__3634\ : InMux
    port map (
            O => \N__17438\,
            I => \N__17434\
        );

    \I__3633\ : InMux
    port map (
            O => \N__17437\,
            I => \N__17431\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__17434\,
            I => \ALL_SYS_PWRGD.countZ0Z_15\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__17431\,
            I => \ALL_SYS_PWRGD.countZ0Z_15\
        );

    \I__3630\ : CascadeMux
    port map (
            O => \N__17426\,
            I => \N__17422\
        );

    \I__3629\ : InMux
    port map (
            O => \N__17425\,
            I => \N__17419\
        );

    \I__3628\ : InMux
    port map (
            O => \N__17422\,
            I => \N__17416\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__17419\,
            I => \ALL_SYS_PWRGD.countZ0Z_13\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__17416\,
            I => \ALL_SYS_PWRGD.countZ0Z_13\
        );

    \I__3625\ : InMux
    port map (
            O => \N__17411\,
            I => \N__17407\
        );

    \I__3624\ : InMux
    port map (
            O => \N__17410\,
            I => \N__17404\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__17407\,
            I => \ALL_SYS_PWRGD.countZ0Z_12\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__17404\,
            I => \ALL_SYS_PWRGD.countZ0Z_12\
        );

    \I__3621\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17396\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__17396\,
            I => \ALL_SYS_PWRGD.un4_count_10\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__17393\,
            I => \ALL_SYS_PWRGD.un4_count_11_cascade_\
        );

    \I__3618\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17387\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__17387\,
            I => \ALL_SYS_PWRGD.un4_count_8\
        );

    \I__3616\ : InMux
    port map (
            O => \N__17384\,
            I => \N__17380\
        );

    \I__3615\ : InMux
    port map (
            O => \N__17383\,
            I => \N__17377\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__17380\,
            I => \ALL_SYS_PWRGD.countZ0Z_1\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__17377\,
            I => \ALL_SYS_PWRGD.countZ0Z_1\
        );

    \I__3612\ : InMux
    port map (
            O => \N__17372\,
            I => \N__17368\
        );

    \I__3611\ : InMux
    port map (
            O => \N__17371\,
            I => \N__17365\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__17368\,
            I => \ALL_SYS_PWRGD.countZ0Z_9\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__17365\,
            I => \ALL_SYS_PWRGD.countZ0Z_9\
        );

    \I__3608\ : CascadeMux
    port map (
            O => \N__17360\,
            I => \N__17356\
        );

    \I__3607\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17353\
        );

    \I__3606\ : InMux
    port map (
            O => \N__17356\,
            I => \N__17350\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__17353\,
            I => \ALL_SYS_PWRGD.countZ0Z_10\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__17350\,
            I => \ALL_SYS_PWRGD.countZ0Z_10\
        );

    \I__3603\ : InMux
    port map (
            O => \N__17345\,
            I => \N__17341\
        );

    \I__3602\ : InMux
    port map (
            O => \N__17344\,
            I => \N__17338\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__17341\,
            I => \ALL_SYS_PWRGD.countZ0Z_0\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__17338\,
            I => \ALL_SYS_PWRGD.countZ0Z_0\
        );

    \I__3599\ : InMux
    port map (
            O => \N__17333\,
            I => \COUNTER.counter_1_cry_27\
        );

    \I__3598\ : InMux
    port map (
            O => \N__17330\,
            I => \COUNTER.counter_1_cry_28\
        );

    \I__3597\ : InMux
    port map (
            O => \N__17327\,
            I => \COUNTER.counter_1_cry_29\
        );

    \I__3596\ : InMux
    port map (
            O => \N__17324\,
            I => \COUNTER.counter_1_cry_30\
        );

    \I__3595\ : InMux
    port map (
            O => \N__17321\,
            I => \N__17317\
        );

    \I__3594\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17314\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__17317\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__17314\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__3591\ : InMux
    port map (
            O => \N__17309\,
            I => \N__17305\
        );

    \I__3590\ : InMux
    port map (
            O => \N__17308\,
            I => \N__17302\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__17305\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__17302\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__17297\,
            I => \N__17293\
        );

    \I__3586\ : InMux
    port map (
            O => \N__17296\,
            I => \N__17290\
        );

    \I__3585\ : InMux
    port map (
            O => \N__17293\,
            I => \N__17287\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__17290\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__17287\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__3582\ : InMux
    port map (
            O => \N__17282\,
            I => \N__17278\
        );

    \I__3581\ : InMux
    port map (
            O => \N__17281\,
            I => \N__17275\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__17278\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__17275\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__3578\ : InMux
    port map (
            O => \N__17270\,
            I => \N__17266\
        );

    \I__3577\ : InMux
    port map (
            O => \N__17269\,
            I => \N__17263\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__17266\,
            I => \ALL_SYS_PWRGD.countZ0Z_5\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__17263\,
            I => \ALL_SYS_PWRGD.countZ0Z_5\
        );

    \I__3574\ : InMux
    port map (
            O => \N__17258\,
            I => \N__17254\
        );

    \I__3573\ : InMux
    port map (
            O => \N__17257\,
            I => \N__17251\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__17254\,
            I => \ALL_SYS_PWRGD.countZ0Z_3\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__17251\,
            I => \ALL_SYS_PWRGD.countZ0Z_3\
        );

    \I__3570\ : CascadeMux
    port map (
            O => \N__17246\,
            I => \N__17242\
        );

    \I__3569\ : InMux
    port map (
            O => \N__17245\,
            I => \N__17239\
        );

    \I__3568\ : InMux
    port map (
            O => \N__17242\,
            I => \N__17236\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__17239\,
            I => \ALL_SYS_PWRGD.countZ0Z_11\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__17236\,
            I => \ALL_SYS_PWRGD.countZ0Z_11\
        );

    \I__3565\ : InMux
    port map (
            O => \N__17231\,
            I => \N__17227\
        );

    \I__3564\ : InMux
    port map (
            O => \N__17230\,
            I => \N__17224\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__17227\,
            I => \ALL_SYS_PWRGD.countZ0Z_2\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__17224\,
            I => \ALL_SYS_PWRGD.countZ0Z_2\
        );

    \I__3561\ : InMux
    port map (
            O => \N__17219\,
            I => \N__17215\
        );

    \I__3560\ : InMux
    port map (
            O => \N__17218\,
            I => \N__17212\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__17215\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__17212\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__3557\ : InMux
    port map (
            O => \N__17207\,
            I => \N__17203\
        );

    \I__3556\ : InMux
    port map (
            O => \N__17206\,
            I => \N__17200\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__17203\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__17200\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__17195\,
            I => \N__17191\
        );

    \I__3552\ : InMux
    port map (
            O => \N__17194\,
            I => \N__17188\
        );

    \I__3551\ : InMux
    port map (
            O => \N__17191\,
            I => \N__17185\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__17188\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__17185\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__3548\ : InMux
    port map (
            O => \N__17180\,
            I => \N__17176\
        );

    \I__3547\ : InMux
    port map (
            O => \N__17179\,
            I => \N__17173\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__17176\,
            I => \N__17170\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__17173\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__17170\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__3543\ : InMux
    port map (
            O => \N__17165\,
            I => \N__17161\
        );

    \I__3542\ : InMux
    port map (
            O => \N__17164\,
            I => \N__17158\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__17161\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__17158\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__3539\ : InMux
    port map (
            O => \N__17153\,
            I => \N__17149\
        );

    \I__3538\ : InMux
    port map (
            O => \N__17152\,
            I => \N__17146\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__17149\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__17146\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__17141\,
            I => \N__17137\
        );

    \I__3534\ : InMux
    port map (
            O => \N__17140\,
            I => \N__17134\
        );

    \I__3533\ : InMux
    port map (
            O => \N__17137\,
            I => \N__17131\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__17134\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__17131\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__3530\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17122\
        );

    \I__3529\ : InMux
    port map (
            O => \N__17125\,
            I => \N__17119\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__17122\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__17119\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__3526\ : InMux
    port map (
            O => \N__17114\,
            I => \COUNTER.counter_1_cry_18\
        );

    \I__3525\ : InMux
    port map (
            O => \N__17111\,
            I => \COUNTER.counter_1_cry_19\
        );

    \I__3524\ : InMux
    port map (
            O => \N__17108\,
            I => \COUNTER.counter_1_cry_20\
        );

    \I__3523\ : InMux
    port map (
            O => \N__17105\,
            I => \COUNTER.counter_1_cry_21\
        );

    \I__3522\ : InMux
    port map (
            O => \N__17102\,
            I => \COUNTER.counter_1_cry_22\
        );

    \I__3521\ : InMux
    port map (
            O => \N__17099\,
            I => \COUNTER.counter_1_cry_23\
        );

    \I__3520\ : InMux
    port map (
            O => \N__17096\,
            I => \bfn_9_4_0_\
        );

    \I__3519\ : InMux
    port map (
            O => \N__17093\,
            I => \COUNTER.counter_1_cry_25\
        );

    \I__3518\ : InMux
    port map (
            O => \N__17090\,
            I => \COUNTER.counter_1_cry_26\
        );

    \I__3517\ : InMux
    port map (
            O => \N__17087\,
            I => \COUNTER.counter_1_cry_9\
        );

    \I__3516\ : InMux
    port map (
            O => \N__17084\,
            I => \COUNTER.counter_1_cry_10\
        );

    \I__3515\ : InMux
    port map (
            O => \N__17081\,
            I => \COUNTER.counter_1_cry_11\
        );

    \I__3514\ : InMux
    port map (
            O => \N__17078\,
            I => \COUNTER.counter_1_cry_12\
        );

    \I__3513\ : InMux
    port map (
            O => \N__17075\,
            I => \COUNTER.counter_1_cry_13\
        );

    \I__3512\ : InMux
    port map (
            O => \N__17072\,
            I => \COUNTER.counter_1_cry_14\
        );

    \I__3511\ : InMux
    port map (
            O => \N__17069\,
            I => \COUNTER.counter_1_cry_15\
        );

    \I__3510\ : InMux
    port map (
            O => \N__17066\,
            I => \bfn_9_3_0_\
        );

    \I__3509\ : InMux
    port map (
            O => \N__17063\,
            I => \COUNTER.counter_1_cry_17\
        );

    \I__3508\ : InMux
    port map (
            O => \N__17060\,
            I => \COUNTER.counter_1_cry_1\
        );

    \I__3507\ : InMux
    port map (
            O => \N__17057\,
            I => \COUNTER.counter_1_cry_2\
        );

    \I__3506\ : InMux
    port map (
            O => \N__17054\,
            I => \COUNTER.counter_1_cry_3\
        );

    \I__3505\ : InMux
    port map (
            O => \N__17051\,
            I => \N__17046\
        );

    \I__3504\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17041\
        );

    \I__3503\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17041\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__17046\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__17041\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__3500\ : InMux
    port map (
            O => \N__17036\,
            I => \N__17033\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__17033\,
            I => \COUNTER.counter_1_cry_4_THRU_CO\
        );

    \I__3498\ : InMux
    port map (
            O => \N__17030\,
            I => \COUNTER.counter_1_cry_4\
        );

    \I__3497\ : CascadeMux
    port map (
            O => \N__17027\,
            I => \N__17023\
        );

    \I__3496\ : InMux
    port map (
            O => \N__17026\,
            I => \N__17019\
        );

    \I__3495\ : InMux
    port map (
            O => \N__17023\,
            I => \N__17014\
        );

    \I__3494\ : InMux
    port map (
            O => \N__17022\,
            I => \N__17014\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__17019\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__17014\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__3491\ : InMux
    port map (
            O => \N__17009\,
            I => \N__17006\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__17006\,
            I => \COUNTER.counter_1_cry_5_THRU_CO\
        );

    \I__3489\ : InMux
    port map (
            O => \N__17003\,
            I => \COUNTER.counter_1_cry_5\
        );

    \I__3488\ : CascadeMux
    port map (
            O => \N__17000\,
            I => \N__16996\
        );

    \I__3487\ : InMux
    port map (
            O => \N__16999\,
            I => \N__16993\
        );

    \I__3486\ : InMux
    port map (
            O => \N__16996\,
            I => \N__16990\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__16993\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__16990\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__3483\ : InMux
    port map (
            O => \N__16985\,
            I => \COUNTER.counter_1_cry_6\
        );

    \I__3482\ : InMux
    port map (
            O => \N__16982\,
            I => \COUNTER.counter_1_cry_7\
        );

    \I__3481\ : InMux
    port map (
            O => \N__16979\,
            I => \bfn_9_2_0_\
        );

    \I__3480\ : InMux
    port map (
            O => \N__16976\,
            I => \VPP_VDDQ.un1_count_1_cry_8\
        );

    \I__3479\ : InMux
    port map (
            O => \N__16973\,
            I => \VPP_VDDQ.un1_count_1_cry_9\
        );

    \I__3478\ : InMux
    port map (
            O => \N__16970\,
            I => \VPP_VDDQ.un1_count_1_cry_10\
        );

    \I__3477\ : InMux
    port map (
            O => \N__16967\,
            I => \VPP_VDDQ.un1_count_1_cry_11\
        );

    \I__3476\ : InMux
    port map (
            O => \N__16964\,
            I => \VPP_VDDQ.un1_count_1_cry_12\
        );

    \I__3475\ : InMux
    port map (
            O => \N__16961\,
            I => \VPP_VDDQ.un1_count_1_cry_13\
        );

    \I__3474\ : InMux
    port map (
            O => \N__16958\,
            I => \bfn_8_16_0_\
        );

    \I__3473\ : CEMux
    port map (
            O => \N__16955\,
            I => \N__16952\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__16952\,
            I => \N__16949\
        );

    \I__3471\ : Odrv4
    port map (
            O => \N__16949\,
            I => \VPP_VDDQ.N_65_1\
        );

    \I__3470\ : SRMux
    port map (
            O => \N__16946\,
            I => \N__16943\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__16943\,
            I => \N__16939\
        );

    \I__3468\ : SRMux
    port map (
            O => \N__16942\,
            I => \N__16936\
        );

    \I__3467\ : Span4Mux_s1_v
    port map (
            O => \N__16939\,
            I => \N__16931\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__16936\,
            I => \N__16931\
        );

    \I__3465\ : Span4Mux_v
    port map (
            O => \N__16931\,
            I => \N__16927\
        );

    \I__3464\ : SRMux
    port map (
            O => \N__16930\,
            I => \N__16924\
        );

    \I__3463\ : Sp12to4
    port map (
            O => \N__16927\,
            I => \N__16918\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__16924\,
            I => \N__16918\
        );

    \I__3461\ : InMux
    port map (
            O => \N__16923\,
            I => \N__16915\
        );

    \I__3460\ : Odrv12
    port map (
            O => \N__16918\,
            I => \VPP_VDDQ.curr_state_RNIGR9S7Z0Z_0\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__16915\,
            I => \VPP_VDDQ.curr_state_RNIGR9S7Z0Z_0\
        );

    \I__3458\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16905\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16909\,
            I => \N__16900\
        );

    \I__3456\ : InMux
    port map (
            O => \N__16908\,
            I => \N__16900\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__16905\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__16900\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__3453\ : InMux
    port map (
            O => \N__16895\,
            I => \N__16891\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__16894\,
            I => \N__16888\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__16891\,
            I => \N__16885\
        );

    \I__3450\ : InMux
    port map (
            O => \N__16888\,
            I => \N__16882\
        );

    \I__3449\ : Odrv4
    port map (
            O => \N__16885\,
            I => \VPP_VDDQ.N_108_i\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__16882\,
            I => \VPP_VDDQ.N_108_i\
        );

    \I__3447\ : InMux
    port map (
            O => \N__16877\,
            I => \VPP_VDDQ.un1_count_1_cry_0\
        );

    \I__3446\ : InMux
    port map (
            O => \N__16874\,
            I => \VPP_VDDQ.un1_count_1_cry_1\
        );

    \I__3445\ : InMux
    port map (
            O => \N__16871\,
            I => \VPP_VDDQ.un1_count_1_cry_2\
        );

    \I__3444\ : InMux
    port map (
            O => \N__16868\,
            I => \VPP_VDDQ.un1_count_1_cry_3\
        );

    \I__3443\ : InMux
    port map (
            O => \N__16865\,
            I => \VPP_VDDQ.un1_count_1_cry_4\
        );

    \I__3442\ : InMux
    port map (
            O => \N__16862\,
            I => \VPP_VDDQ.un1_count_1_cry_5\
        );

    \I__3441\ : InMux
    port map (
            O => \N__16859\,
            I => \VPP_VDDQ.un1_count_1_cry_6\
        );

    \I__3440\ : InMux
    port map (
            O => \N__16856\,
            I => \bfn_8_15_0_\
        );

    \I__3439\ : InMux
    port map (
            O => \N__16853\,
            I => \bfn_8_12_0_\
        );

    \I__3438\ : InMux
    port map (
            O => \N__16850\,
            I => \RSMRST_PWRGD.un1_count_1_cry_8\
        );

    \I__3437\ : InMux
    port map (
            O => \N__16847\,
            I => \RSMRST_PWRGD.un1_count_1_cry_9\
        );

    \I__3436\ : InMux
    port map (
            O => \N__16844\,
            I => \RSMRST_PWRGD.un1_count_1_cry_10\
        );

    \I__3435\ : InMux
    port map (
            O => \N__16841\,
            I => \RSMRST_PWRGD.un1_count_1_cry_11\
        );

    \I__3434\ : InMux
    port map (
            O => \N__16838\,
            I => \RSMRST_PWRGD.un1_count_1_cry_12\
        );

    \I__3433\ : InMux
    port map (
            O => \N__16835\,
            I => \RSMRST_PWRGD.un1_count_1_cry_13\
        );

    \I__3432\ : InMux
    port map (
            O => \N__16832\,
            I => \bfn_8_13_0_\
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__16829\,
            I => \POWERLED.count_off_1_sqmuxa_i_a6_0_1_cascade_\
        );

    \I__3430\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16822\
        );

    \I__3429\ : InMux
    port map (
            O => \N__16825\,
            I => \N__16819\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__16822\,
            I => \POWERLED.N_136\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__16819\,
            I => \POWERLED.N_136\
        );

    \I__3426\ : InMux
    port map (
            O => \N__16814\,
            I => \N__16811\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__16811\,
            I => \N__16808\
        );

    \I__3424\ : Odrv4
    port map (
            O => \N__16808\,
            I => \POWERLED.count_off_1_sqmuxa_i_a6_0_3\
        );

    \I__3423\ : InMux
    port map (
            O => \N__16805\,
            I => \RSMRST_PWRGD.un1_count_1_cry_0\
        );

    \I__3422\ : InMux
    port map (
            O => \N__16802\,
            I => \RSMRST_PWRGD.un1_count_1_cry_1\
        );

    \I__3421\ : InMux
    port map (
            O => \N__16799\,
            I => \RSMRST_PWRGD.un1_count_1_cry_2\
        );

    \I__3420\ : InMux
    port map (
            O => \N__16796\,
            I => \RSMRST_PWRGD.un1_count_1_cry_3\
        );

    \I__3419\ : InMux
    port map (
            O => \N__16793\,
            I => \RSMRST_PWRGD.un1_count_1_cry_4\
        );

    \I__3418\ : InMux
    port map (
            O => \N__16790\,
            I => \RSMRST_PWRGD.un1_count_1_cry_5\
        );

    \I__3417\ : InMux
    port map (
            O => \N__16787\,
            I => \RSMRST_PWRGD.un1_count_1_cry_6\
        );

    \I__3416\ : InMux
    port map (
            O => \N__16784\,
            I => \N__16781\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__16781\,
            I => \N__16778\
        );

    \I__3414\ : Odrv4
    port map (
            O => \N__16778\,
            I => \POWERLED.N_366_1\
        );

    \I__3413\ : InMux
    port map (
            O => \N__16775\,
            I => \N__16762\
        );

    \I__3412\ : InMux
    port map (
            O => \N__16774\,
            I => \N__16762\
        );

    \I__3411\ : InMux
    port map (
            O => \N__16773\,
            I => \N__16762\
        );

    \I__3410\ : InMux
    port map (
            O => \N__16772\,
            I => \N__16753\
        );

    \I__3409\ : InMux
    port map (
            O => \N__16771\,
            I => \N__16746\
        );

    \I__3408\ : InMux
    port map (
            O => \N__16770\,
            I => \N__16746\
        );

    \I__3407\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16746\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__16762\,
            I => \N__16743\
        );

    \I__3405\ : InMux
    port map (
            O => \N__16761\,
            I => \N__16740\
        );

    \I__3404\ : InMux
    port map (
            O => \N__16760\,
            I => \N__16732\
        );

    \I__3403\ : InMux
    port map (
            O => \N__16759\,
            I => \N__16723\
        );

    \I__3402\ : InMux
    port map (
            O => \N__16758\,
            I => \N__16723\
        );

    \I__3401\ : InMux
    port map (
            O => \N__16757\,
            I => \N__16723\
        );

    \I__3400\ : InMux
    port map (
            O => \N__16756\,
            I => \N__16723\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__16753\,
            I => \N__16720\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__16746\,
            I => \N__16717\
        );

    \I__3397\ : Span4Mux_v
    port map (
            O => \N__16743\,
            I => \N__16712\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__16740\,
            I => \N__16712\
        );

    \I__3395\ : InMux
    port map (
            O => \N__16739\,
            I => \N__16709\
        );

    \I__3394\ : InMux
    port map (
            O => \N__16738\,
            I => \N__16700\
        );

    \I__3393\ : InMux
    port map (
            O => \N__16737\,
            I => \N__16700\
        );

    \I__3392\ : InMux
    port map (
            O => \N__16736\,
            I => \N__16700\
        );

    \I__3391\ : InMux
    port map (
            O => \N__16735\,
            I => \N__16700\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__16732\,
            I => \N__16697\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__16723\,
            I => \N__16692\
        );

    \I__3388\ : Span4Mux_h
    port map (
            O => \N__16720\,
            I => \N__16692\
        );

    \I__3387\ : Span4Mux_h
    port map (
            O => \N__16717\,
            I => \N__16687\
        );

    \I__3386\ : Span4Mux_h
    port map (
            O => \N__16712\,
            I => \N__16687\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__16709\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__16700\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__16697\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__3382\ : Odrv4
    port map (
            O => \N__16692\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__3381\ : Odrv4
    port map (
            O => \N__16687\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__3380\ : InMux
    port map (
            O => \N__16676\,
            I => \N__16673\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__16673\,
            I => \N__16669\
        );

    \I__3378\ : CascadeMux
    port map (
            O => \N__16672\,
            I => \N__16666\
        );

    \I__3377\ : Span4Mux_h
    port map (
            O => \N__16669\,
            I => \N__16663\
        );

    \I__3376\ : InMux
    port map (
            O => \N__16666\,
            I => \N__16660\
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__16663\,
            I => \POWERLED.N_177_5\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__16660\,
            I => \POWERLED.N_177_5\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__16655\,
            I => \POWERLED.count_clk_0_sqmuxa_5_0_o2_0_0_cascade_\
        );

    \I__3372\ : InMux
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__3370\ : Span4Mux_v
    port map (
            O => \N__16646\,
            I => \N__16642\
        );

    \I__3369\ : InMux
    port map (
            O => \N__16645\,
            I => \N__16639\
        );

    \I__3368\ : Odrv4
    port map (
            O => \N__16642\,
            I => \POWERLED.N_141\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__16639\,
            I => \POWERLED.N_141\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__16634\,
            I => \POWERLED.N_136_cascade_\
        );

    \I__3365\ : InMux
    port map (
            O => \N__16631\,
            I => \N__16624\
        );

    \I__3364\ : InMux
    port map (
            O => \N__16630\,
            I => \N__16624\
        );

    \I__3363\ : InMux
    port map (
            O => \N__16629\,
            I => \N__16620\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__16624\,
            I => \N__16617\
        );

    \I__3361\ : InMux
    port map (
            O => \N__16623\,
            I => \N__16614\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__16620\,
            I => \POWERLED.N_146\
        );

    \I__3359\ : Odrv4
    port map (
            O => \N__16617\,
            I => \POWERLED.N_146\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__16614\,
            I => \POWERLED.N_146\
        );

    \I__3357\ : InMux
    port map (
            O => \N__16607\,
            I => \N__16604\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__16604\,
            I => \N__16601\
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__16601\,
            I => \POWERLED.count_clk_0_sqmuxa_5_0_a6_1\
        );

    \I__3354\ : InMux
    port map (
            O => \N__16598\,
            I => \N__16595\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__16595\,
            I => \POWERLED.count_clk_0_sqmuxa_5_0_o2_4\
        );

    \I__3352\ : IoInMux
    port map (
            O => \N__16592\,
            I => \N__16587\
        );

    \I__3351\ : CascadeMux
    port map (
            O => \N__16591\,
            I => \N__16584\
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__16590\,
            I => \N__16578\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__16587\,
            I => \N__16574\
        );

    \I__3348\ : InMux
    port map (
            O => \N__16584\,
            I => \N__16567\
        );

    \I__3347\ : InMux
    port map (
            O => \N__16583\,
            I => \N__16567\
        );

    \I__3346\ : InMux
    port map (
            O => \N__16582\,
            I => \N__16567\
        );

    \I__3345\ : InMux
    port map (
            O => \N__16581\,
            I => \N__16564\
        );

    \I__3344\ : InMux
    port map (
            O => \N__16578\,
            I => \N__16561\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__16577\,
            I => \N__16558\
        );

    \I__3342\ : IoSpan4Mux
    port map (
            O => \N__16574\,
            I => \N__16553\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__16567\,
            I => \N__16546\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__16564\,
            I => \N__16546\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__16561\,
            I => \N__16546\
        );

    \I__3338\ : InMux
    port map (
            O => \N__16558\,
            I => \N__16543\
        );

    \I__3337\ : InMux
    port map (
            O => \N__16557\,
            I => \N__16538\
        );

    \I__3336\ : InMux
    port map (
            O => \N__16556\,
            I => \N__16538\
        );

    \I__3335\ : Span4Mux_s2_h
    port map (
            O => \N__16553\,
            I => \N__16534\
        );

    \I__3334\ : Span4Mux_v
    port map (
            O => \N__16546\,
            I => \N__16531\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__16543\,
            I => \N__16528\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__16538\,
            I => \N__16525\
        );

    \I__3331\ : InMux
    port map (
            O => \N__16537\,
            I => \N__16522\
        );

    \I__3330\ : Span4Mux_h
    port map (
            O => \N__16534\,
            I => \N__16517\
        );

    \I__3329\ : Span4Mux_v
    port map (
            O => \N__16531\,
            I => \N__16517\
        );

    \I__3328\ : Sp12to4
    port map (
            O => \N__16528\,
            I => \N__16510\
        );

    \I__3327\ : Sp12to4
    port map (
            O => \N__16525\,
            I => \N__16510\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__16522\,
            I => \N__16510\
        );

    \I__3325\ : Sp12to4
    port map (
            O => \N__16517\,
            I => \N__16505\
        );

    \I__3324\ : Span12Mux_v
    port map (
            O => \N__16510\,
            I => \N__16505\
        );

    \I__3323\ : Odrv12
    port map (
            O => \N__16505\,
            I => gpio_fpga_soc_4
        );

    \I__3322\ : InMux
    port map (
            O => \N__16502\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_12\
        );

    \I__3321\ : InMux
    port map (
            O => \N__16499\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_13\
        );

    \I__3320\ : InMux
    port map (
            O => \N__16496\,
            I => \bfn_8_7_0_\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__16493\,
            I => \N__16490\
        );

    \I__3318\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16486\
        );

    \I__3317\ : InMux
    port map (
            O => \N__16489\,
            I => \N__16483\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__16486\,
            I => \N__16480\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__16483\,
            I => \N__16477\
        );

    \I__3314\ : Span4Mux_h
    port map (
            O => \N__16480\,
            I => \N__16474\
        );

    \I__3313\ : Odrv4
    port map (
            O => \N__16477\,
            I => \POWERLED.dutycycle_RNIO18NZ0Z_9\
        );

    \I__3312\ : Odrv4
    port map (
            O => \N__16474\,
            I => \POWERLED.dutycycle_RNIO18NZ0Z_9\
        );

    \I__3311\ : CascadeMux
    port map (
            O => \N__16469\,
            I => \N__16462\
        );

    \I__3310\ : InMux
    port map (
            O => \N__16468\,
            I => \N__16453\
        );

    \I__3309\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16453\
        );

    \I__3308\ : CascadeMux
    port map (
            O => \N__16466\,
            I => \N__16449\
        );

    \I__3307\ : InMux
    port map (
            O => \N__16465\,
            I => \N__16445\
        );

    \I__3306\ : InMux
    port map (
            O => \N__16462\,
            I => \N__16442\
        );

    \I__3305\ : InMux
    port map (
            O => \N__16461\,
            I => \N__16439\
        );

    \I__3304\ : InMux
    port map (
            O => \N__16460\,
            I => \N__16434\
        );

    \I__3303\ : InMux
    port map (
            O => \N__16459\,
            I => \N__16434\
        );

    \I__3302\ : InMux
    port map (
            O => \N__16458\,
            I => \N__16431\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__16453\,
            I => \N__16428\
        );

    \I__3300\ : InMux
    port map (
            O => \N__16452\,
            I => \N__16425\
        );

    \I__3299\ : InMux
    port map (
            O => \N__16449\,
            I => \N__16420\
        );

    \I__3298\ : InMux
    port map (
            O => \N__16448\,
            I => \N__16420\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__16445\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__16442\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__16439\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__16434\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__16431\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__3292\ : Odrv12
    port map (
            O => \N__16428\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__16425\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__16420\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__16403\,
            I => \N__16399\
        );

    \I__3288\ : CascadeMux
    port map (
            O => \N__16402\,
            I => \N__16390\
        );

    \I__3287\ : InMux
    port map (
            O => \N__16399\,
            I => \N__16381\
        );

    \I__3286\ : InMux
    port map (
            O => \N__16398\,
            I => \N__16381\
        );

    \I__3285\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16381\
        );

    \I__3284\ : InMux
    port map (
            O => \N__16396\,
            I => \N__16378\
        );

    \I__3283\ : InMux
    port map (
            O => \N__16395\,
            I => \N__16375\
        );

    \I__3282\ : InMux
    port map (
            O => \N__16394\,
            I => \N__16372\
        );

    \I__3281\ : InMux
    port map (
            O => \N__16393\,
            I => \N__16367\
        );

    \I__3280\ : InMux
    port map (
            O => \N__16390\,
            I => \N__16367\
        );

    \I__3279\ : InMux
    port map (
            O => \N__16389\,
            I => \N__16362\
        );

    \I__3278\ : InMux
    port map (
            O => \N__16388\,
            I => \N__16362\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__16381\,
            I => \N__16359\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__16378\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__16375\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__16372\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__16367\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__16362\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__3271\ : Odrv4
    port map (
            O => \N__16359\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__3270\ : CascadeMux
    port map (
            O => \N__16346\,
            I => \N__16340\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__16345\,
            I => \N__16336\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__16344\,
            I => \N__16331\
        );

    \I__3267\ : InMux
    port map (
            O => \N__16343\,
            I => \N__16326\
        );

    \I__3266\ : InMux
    port map (
            O => \N__16340\,
            I => \N__16323\
        );

    \I__3265\ : InMux
    port map (
            O => \N__16339\,
            I => \N__16318\
        );

    \I__3264\ : InMux
    port map (
            O => \N__16336\,
            I => \N__16318\
        );

    \I__3263\ : InMux
    port map (
            O => \N__16335\,
            I => \N__16315\
        );

    \I__3262\ : InMux
    port map (
            O => \N__16334\,
            I => \N__16312\
        );

    \I__3261\ : InMux
    port map (
            O => \N__16331\,
            I => \N__16305\
        );

    \I__3260\ : InMux
    port map (
            O => \N__16330\,
            I => \N__16305\
        );

    \I__3259\ : InMux
    port map (
            O => \N__16329\,
            I => \N__16305\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__16326\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__16323\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__16318\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__16315\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__16312\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__16305\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__3252\ : CascadeMux
    port map (
            O => \N__16292\,
            I => \N__16289\
        );

    \I__3251\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16276\
        );

    \I__3250\ : InMux
    port map (
            O => \N__16288\,
            I => \N__16276\
        );

    \I__3249\ : InMux
    port map (
            O => \N__16287\,
            I => \N__16273\
        );

    \I__3248\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16268\
        );

    \I__3247\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16268\
        );

    \I__3246\ : InMux
    port map (
            O => \N__16284\,
            I => \N__16265\
        );

    \I__3245\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16258\
        );

    \I__3244\ : InMux
    port map (
            O => \N__16282\,
            I => \N__16258\
        );

    \I__3243\ : InMux
    port map (
            O => \N__16281\,
            I => \N__16258\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__16276\,
            I => \N__16255\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__16273\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__16268\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__16265\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__16258\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__16255\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__16244\,
            I => \N__16239\
        );

    \I__3235\ : InMux
    port map (
            O => \N__16243\,
            I => \N__16232\
        );

    \I__3234\ : InMux
    port map (
            O => \N__16242\,
            I => \N__16228\
        );

    \I__3233\ : InMux
    port map (
            O => \N__16239\,
            I => \N__16225\
        );

    \I__3232\ : InMux
    port map (
            O => \N__16238\,
            I => \N__16222\
        );

    \I__3231\ : InMux
    port map (
            O => \N__16237\,
            I => \N__16219\
        );

    \I__3230\ : InMux
    port map (
            O => \N__16236\,
            I => \N__16216\
        );

    \I__3229\ : InMux
    port map (
            O => \N__16235\,
            I => \N__16213\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__16232\,
            I => \N__16210\
        );

    \I__3227\ : InMux
    port map (
            O => \N__16231\,
            I => \N__16207\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__16228\,
            I => \N__16204\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__16225\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__16222\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__16219\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__16216\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__16213\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__16210\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__16207\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__16204\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__16187\,
            I => \N__16181\
        );

    \I__3216\ : InMux
    port map (
            O => \N__16186\,
            I => \N__16177\
        );

    \I__3215\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16174\
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__16184\,
            I => \N__16169\
        );

    \I__3213\ : InMux
    port map (
            O => \N__16181\,
            I => \N__16164\
        );

    \I__3212\ : InMux
    port map (
            O => \N__16180\,
            I => \N__16161\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__16177\,
            I => \N__16156\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__16174\,
            I => \N__16156\
        );

    \I__3209\ : InMux
    port map (
            O => \N__16173\,
            I => \N__16149\
        );

    \I__3208\ : InMux
    port map (
            O => \N__16172\,
            I => \N__16149\
        );

    \I__3207\ : InMux
    port map (
            O => \N__16169\,
            I => \N__16149\
        );

    \I__3206\ : InMux
    port map (
            O => \N__16168\,
            I => \N__16146\
        );

    \I__3205\ : InMux
    port map (
            O => \N__16167\,
            I => \N__16143\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__16164\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__16161\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__3202\ : Odrv4
    port map (
            O => \N__16156\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__16149\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__16146\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__16143\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__16130\,
            I => \N__16125\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__16129\,
            I => \N__16122\
        );

    \I__3196\ : InMux
    port map (
            O => \N__16128\,
            I => \N__16119\
        );

    \I__3195\ : InMux
    port map (
            O => \N__16125\,
            I => \N__16112\
        );

    \I__3194\ : InMux
    port map (
            O => \N__16122\,
            I => \N__16109\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__16119\,
            I => \N__16106\
        );

    \I__3192\ : InMux
    port map (
            O => \N__16118\,
            I => \N__16103\
        );

    \I__3191\ : InMux
    port map (
            O => \N__16117\,
            I => \N__16098\
        );

    \I__3190\ : InMux
    port map (
            O => \N__16116\,
            I => \N__16098\
        );

    \I__3189\ : InMux
    port map (
            O => \N__16115\,
            I => \N__16095\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__16112\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__16109\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__16106\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__16103\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__16098\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__16095\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3182\ : InMux
    port map (
            O => \N__16082\,
            I => \N__16077\
        );

    \I__3181\ : InMux
    port map (
            O => \N__16081\,
            I => \N__16074\
        );

    \I__3180\ : InMux
    port map (
            O => \N__16080\,
            I => \N__16069\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__16077\,
            I => \N__16062\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__16074\,
            I => \N__16059\
        );

    \I__3177\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16056\
        );

    \I__3176\ : InMux
    port map (
            O => \N__16072\,
            I => \N__16053\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__16069\,
            I => \N__16050\
        );

    \I__3174\ : InMux
    port map (
            O => \N__16068\,
            I => \N__16043\
        );

    \I__3173\ : InMux
    port map (
            O => \N__16067\,
            I => \N__16043\
        );

    \I__3172\ : InMux
    port map (
            O => \N__16066\,
            I => \N__16043\
        );

    \I__3171\ : InMux
    port map (
            O => \N__16065\,
            I => \N__16040\
        );

    \I__3170\ : Span4Mux_h
    port map (
            O => \N__16062\,
            I => \N__16035\
        );

    \I__3169\ : Span4Mux_h
    port map (
            O => \N__16059\,
            I => \N__16035\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__16056\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__16053\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3166\ : Odrv4
    port map (
            O => \N__16050\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__16043\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__16040\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3163\ : Odrv4
    port map (
            O => \N__16035\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__3162\ : InMux
    port map (
            O => \N__16022\,
            I => \N__16019\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__16019\,
            I => \POWERLED.un2_slp_s3n_2_0_o2_3_7\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__16016\,
            I => \POWERLED.un2_slp_s3n_2_0_o2_3_8_cascade_\
        );

    \I__3159\ : InMux
    port map (
            O => \N__16013\,
            I => \N__16010\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__16010\,
            I => \N__16007\
        );

    \I__3157\ : Span4Mux_v
    port map (
            O => \N__16007\,
            I => \N__16004\
        );

    \I__3156\ : Odrv4
    port map (
            O => \N__16004\,
            I => \POWERLED.un2_slp_s3n_2_0_o2_3_6\
        );

    \I__3155\ : InMux
    port map (
            O => \N__16001\,
            I => \N__15993\
        );

    \I__3154\ : InMux
    port map (
            O => \N__16000\,
            I => \N__15990\
        );

    \I__3153\ : InMux
    port map (
            O => \N__15999\,
            I => \N__15981\
        );

    \I__3152\ : InMux
    port map (
            O => \N__15998\,
            I => \N__15981\
        );

    \I__3151\ : InMux
    port map (
            O => \N__15997\,
            I => \N__15981\
        );

    \I__3150\ : InMux
    port map (
            O => \N__15996\,
            I => \N__15981\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__15993\,
            I => \N__15978\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__15990\,
            I => \N__15975\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__15981\,
            I => \N__15972\
        );

    \I__3146\ : Span4Mux_h
    port map (
            O => \N__15978\,
            I => \N__15969\
        );

    \I__3145\ : Span4Mux_h
    port map (
            O => \N__15975\,
            I => \N__15966\
        );

    \I__3144\ : Span4Mux_h
    port map (
            O => \N__15972\,
            I => \N__15963\
        );

    \I__3143\ : Odrv4
    port map (
            O => \N__15969\,
            I => \POWERLED.N_112\
        );

    \I__3142\ : Odrv4
    port map (
            O => \N__15966\,
            I => \POWERLED.N_112\
        );

    \I__3141\ : Odrv4
    port map (
            O => \N__15963\,
            I => \POWERLED.N_112\
        );

    \I__3140\ : InMux
    port map (
            O => \N__15956\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_3\
        );

    \I__3139\ : InMux
    port map (
            O => \N__15953\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_4\
        );

    \I__3138\ : InMux
    port map (
            O => \N__15950\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_5\
        );

    \I__3137\ : InMux
    port map (
            O => \N__15947\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_6\
        );

    \I__3136\ : InMux
    port map (
            O => \N__15944\,
            I => \bfn_8_6_0_\
        );

    \I__3135\ : InMux
    port map (
            O => \N__15941\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_8\
        );

    \I__3134\ : InMux
    port map (
            O => \N__15938\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_9\
        );

    \I__3133\ : InMux
    port map (
            O => \N__15935\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_10\
        );

    \I__3132\ : InMux
    port map (
            O => \N__15932\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_11\
        );

    \I__3131\ : InMux
    port map (
            O => \N__15929\,
            I => \N__15926\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__15926\,
            I => \N__15923\
        );

    \I__3129\ : Span4Mux_h
    port map (
            O => \N__15923\,
            I => \N__15920\
        );

    \I__3128\ : Odrv4
    port map (
            O => \N__15920\,
            I => \HDA_STRAP.count_RNO_0Z0Z_6\
        );

    \I__3127\ : CascadeMux
    port map (
            O => \N__15917\,
            I => \N__15911\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__15916\,
            I => \N__15908\
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__15915\,
            I => \N__15905\
        );

    \I__3124\ : InMux
    port map (
            O => \N__15914\,
            I => \N__15896\
        );

    \I__3123\ : InMux
    port map (
            O => \N__15911\,
            I => \N__15891\
        );

    \I__3122\ : InMux
    port map (
            O => \N__15908\,
            I => \N__15891\
        );

    \I__3121\ : InMux
    port map (
            O => \N__15905\,
            I => \N__15886\
        );

    \I__3120\ : InMux
    port map (
            O => \N__15904\,
            I => \N__15886\
        );

    \I__3119\ : InMux
    port map (
            O => \N__15903\,
            I => \N__15883\
        );

    \I__3118\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15880\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__15901\,
            I => \N__15876\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__15900\,
            I => \N__15873\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__15899\,
            I => \N__15869\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__15896\,
            I => \N__15864\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__15891\,
            I => \N__15855\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__15886\,
            I => \N__15855\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__15883\,
            I => \N__15855\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__15880\,
            I => \N__15855\
        );

    \I__3109\ : InMux
    port map (
            O => \N__15879\,
            I => \N__15852\
        );

    \I__3108\ : InMux
    port map (
            O => \N__15876\,
            I => \N__15849\
        );

    \I__3107\ : InMux
    port map (
            O => \N__15873\,
            I => \N__15846\
        );

    \I__3106\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15839\
        );

    \I__3105\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15839\
        );

    \I__3104\ : InMux
    port map (
            O => \N__15868\,
            I => \N__15839\
        );

    \I__3103\ : InMux
    port map (
            O => \N__15867\,
            I => \N__15836\
        );

    \I__3102\ : Span4Mux_v
    port map (
            O => \N__15864\,
            I => \N__15829\
        );

    \I__3101\ : Span4Mux_v
    port map (
            O => \N__15855\,
            I => \N__15829\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__15852\,
            I => \N__15829\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__15849\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__15846\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__15839\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__15836\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__3095\ : Odrv4
    port map (
            O => \N__15829\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__15818\,
            I => \N__15815\
        );

    \I__3093\ : InMux
    port map (
            O => \N__15815\,
            I => \N__15804\
        );

    \I__3092\ : InMux
    port map (
            O => \N__15814\,
            I => \N__15795\
        );

    \I__3091\ : InMux
    port map (
            O => \N__15813\,
            I => \N__15795\
        );

    \I__3090\ : InMux
    port map (
            O => \N__15812\,
            I => \N__15795\
        );

    \I__3089\ : InMux
    port map (
            O => \N__15811\,
            I => \N__15795\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15810\,
            I => \N__15792\
        );

    \I__3087\ : InMux
    port map (
            O => \N__15809\,
            I => \N__15789\
        );

    \I__3086\ : InMux
    port map (
            O => \N__15808\,
            I => \N__15782\
        );

    \I__3085\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15782\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__15804\,
            I => \N__15779\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__15795\,
            I => \N__15770\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__15792\,
            I => \N__15770\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__15789\,
            I => \N__15770\
        );

    \I__3080\ : InMux
    port map (
            O => \N__15788\,
            I => \N__15767\
        );

    \I__3079\ : InMux
    port map (
            O => \N__15787\,
            I => \N__15764\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__15782\,
            I => \N__15761\
        );

    \I__3077\ : Span4Mux_h
    port map (
            O => \N__15779\,
            I => \N__15758\
        );

    \I__3076\ : InMux
    port map (
            O => \N__15778\,
            I => \N__15753\
        );

    \I__3075\ : InMux
    port map (
            O => \N__15777\,
            I => \N__15753\
        );

    \I__3074\ : Span4Mux_s2_v
    port map (
            O => \N__15770\,
            I => \N__15750\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__15767\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__15764\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3071\ : Odrv4
    port map (
            O => \N__15761\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3070\ : Odrv4
    port map (
            O => \N__15758\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__15753\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__15750\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__3067\ : InMux
    port map (
            O => \N__15737\,
            I => \N__15729\
        );

    \I__3066\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15729\
        );

    \I__3065\ : InMux
    port map (
            O => \N__15735\,
            I => \N__15726\
        );

    \I__3064\ : InMux
    port map (
            O => \N__15734\,
            I => \N__15718\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__15729\,
            I => \N__15715\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__15726\,
            I => \N__15712\
        );

    \I__3061\ : InMux
    port map (
            O => \N__15725\,
            I => \N__15703\
        );

    \I__3060\ : InMux
    port map (
            O => \N__15724\,
            I => \N__15703\
        );

    \I__3059\ : InMux
    port map (
            O => \N__15723\,
            I => \N__15703\
        );

    \I__3058\ : InMux
    port map (
            O => \N__15722\,
            I => \N__15703\
        );

    \I__3057\ : InMux
    port map (
            O => \N__15721\,
            I => \N__15700\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__15718\,
            I => \N__15693\
        );

    \I__3055\ : Span4Mux_s1_v
    port map (
            O => \N__15715\,
            I => \N__15693\
        );

    \I__3054\ : Span4Mux_v
    port map (
            O => \N__15712\,
            I => \N__15693\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__15703\,
            I => \HDA_STRAP.count_RNIB5IA5Z0Z_0\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__15700\,
            I => \HDA_STRAP.count_RNIB5IA5Z0Z_0\
        );

    \I__3051\ : Odrv4
    port map (
            O => \N__15693\,
            I => \HDA_STRAP.count_RNIB5IA5Z0Z_0\
        );

    \I__3050\ : InMux
    port map (
            O => \N__15686\,
            I => \N__15683\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__15683\,
            I => \N__15680\
        );

    \I__3048\ : Span4Mux_s1_v
    port map (
            O => \N__15680\,
            I => \N__15676\
        );

    \I__3047\ : InMux
    port map (
            O => \N__15679\,
            I => \N__15673\
        );

    \I__3046\ : Odrv4
    port map (
            O => \N__15676\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__15673\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__3044\ : InMux
    port map (
            O => \N__15668\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_0\
        );

    \I__3043\ : InMux
    port map (
            O => \N__15665\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_1\
        );

    \I__3042\ : InMux
    port map (
            O => \N__15662\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_2\
        );

    \I__3041\ : InMux
    port map (
            O => \N__15659\,
            I => \N__15656\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__15656\,
            I => \N__15653\
        );

    \I__3039\ : Span4Mux_v
    port map (
            O => \N__15653\,
            I => \N__15640\
        );

    \I__3038\ : InMux
    port map (
            O => \N__15652\,
            I => \N__15637\
        );

    \I__3037\ : InMux
    port map (
            O => \N__15651\,
            I => \N__15632\
        );

    \I__3036\ : InMux
    port map (
            O => \N__15650\,
            I => \N__15625\
        );

    \I__3035\ : InMux
    port map (
            O => \N__15649\,
            I => \N__15625\
        );

    \I__3034\ : InMux
    port map (
            O => \N__15648\,
            I => \N__15625\
        );

    \I__3033\ : InMux
    port map (
            O => \N__15647\,
            I => \N__15622\
        );

    \I__3032\ : InMux
    port map (
            O => \N__15646\,
            I => \N__15617\
        );

    \I__3031\ : InMux
    port map (
            O => \N__15645\,
            I => \N__15617\
        );

    \I__3030\ : InMux
    port map (
            O => \N__15644\,
            I => \N__15612\
        );

    \I__3029\ : InMux
    port map (
            O => \N__15643\,
            I => \N__15612\
        );

    \I__3028\ : Span4Mux_h
    port map (
            O => \N__15640\,
            I => \N__15607\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__15637\,
            I => \N__15607\
        );

    \I__3026\ : InMux
    port map (
            O => \N__15636\,
            I => \N__15602\
        );

    \I__3025\ : InMux
    port map (
            O => \N__15635\,
            I => \N__15602\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__15632\,
            I => \N__15597\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__15625\,
            I => \N__15597\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__15622\,
            I => \N_55\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__15617\,
            I => \N_55\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__15612\,
            I => \N_55\
        );

    \I__3019\ : Odrv4
    port map (
            O => \N__15607\,
            I => \N_55\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__15602\,
            I => \N_55\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__15597\,
            I => \N_55\
        );

    \I__3016\ : InMux
    port map (
            O => \N__15584\,
            I => \N__15576\
        );

    \I__3015\ : InMux
    port map (
            O => \N__15583\,
            I => \N__15576\
        );

    \I__3014\ : InMux
    port map (
            O => \N__15582\,
            I => \N__15571\
        );

    \I__3013\ : InMux
    port map (
            O => \N__15581\,
            I => \N__15571\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__15576\,
            I => \VPP_VDDQ.N_238\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__15571\,
            I => \VPP_VDDQ.N_238\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__15566\,
            I => \VPP_VDDQ.N_238_cascade_\
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__15563\,
            I => \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\
        );

    \I__3008\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15557\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__15557\,
            I => \VPP_VDDQ.G_127_0\
        );

    \I__3006\ : InMux
    port map (
            O => \N__15554\,
            I => \N__15550\
        );

    \I__3005\ : InMux
    port map (
            O => \N__15553\,
            I => \N__15547\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__15550\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__15547\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__3002\ : InMux
    port map (
            O => \N__15542\,
            I => \N__15532\
        );

    \I__3001\ : InMux
    port map (
            O => \N__15541\,
            I => \N__15532\
        );

    \I__3000\ : InMux
    port map (
            O => \N__15540\,
            I => \N__15529\
        );

    \I__2999\ : InMux
    port map (
            O => \N__15539\,
            I => \N__15526\
        );

    \I__2998\ : InMux
    port map (
            O => \N__15538\,
            I => \N__15521\
        );

    \I__2997\ : InMux
    port map (
            O => \N__15537\,
            I => \N__15521\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__15532\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__15529\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__15526\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__15521\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__2992\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15504\
        );

    \I__2991\ : InMux
    port map (
            O => \N__15511\,
            I => \N__15501\
        );

    \I__2990\ : InMux
    port map (
            O => \N__15510\,
            I => \N__15498\
        );

    \I__2989\ : InMux
    port map (
            O => \N__15509\,
            I => \N__15491\
        );

    \I__2988\ : InMux
    port map (
            O => \N__15508\,
            I => \N__15491\
        );

    \I__2987\ : InMux
    port map (
            O => \N__15507\,
            I => \N__15491\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__15504\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__15501\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__15498\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__15491\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__15482\,
            I => \N__15479\
        );

    \I__2981\ : InMux
    port map (
            O => \N__15479\,
            I => \N__15476\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__15476\,
            I => \N__15472\
        );

    \I__2979\ : InMux
    port map (
            O => \N__15475\,
            I => \N__15469\
        );

    \I__2978\ : Odrv4
    port map (
            O => \N__15472\,
            I => \VPP_VDDQ.N_128\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__15469\,
            I => \VPP_VDDQ.N_128\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__15464\,
            I => \VPP_VDDQ.N_154_cascade_\
        );

    \I__2975\ : InMux
    port map (
            O => \N__15461\,
            I => \N__15458\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__15458\,
            I => \POWERLED.count_clk_1_sqmuxa_5_0_1\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__15455\,
            I => \POWERLED.N_127_cascade_\
        );

    \I__2972\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15449\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__15449\,
            I => \POWERLED.count_clk_1_sqmuxa_5_0_0\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__15446\,
            I => \N__15442\
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__15445\,
            I => \N__15439\
        );

    \I__2968\ : InMux
    port map (
            O => \N__15442\,
            I => \N__15435\
        );

    \I__2967\ : InMux
    port map (
            O => \N__15439\,
            I => \N__15432\
        );

    \I__2966\ : InMux
    port map (
            O => \N__15438\,
            I => \N__15429\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__15435\,
            I => \POWERLED.N_88\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__15432\,
            I => \POWERLED.N_88\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__15429\,
            I => \POWERLED.N_88\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__15422\,
            I => \POWERLED.dutycycle_3_sqmuxa_1_i_0_1_1_cascade_\
        );

    \I__2961\ : InMux
    port map (
            O => \N__15419\,
            I => \N__15415\
        );

    \I__2960\ : InMux
    port map (
            O => \N__15418\,
            I => \N__15412\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__15415\,
            I => \POWERLED.N_200_2\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__15412\,
            I => \POWERLED.N_200_2\
        );

    \I__2957\ : InMux
    port map (
            O => \N__15407\,
            I => \N__15404\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__15404\,
            I => \POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_1\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__15401\,
            I => \POWERLED.N_366_1_cascade_\
        );

    \I__2954\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15395\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__15395\,
            I => \POWERLED.N_251\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__15392\,
            I => \N__15389\
        );

    \I__2951\ : InMux
    port map (
            O => \N__15389\,
            I => \N__15385\
        );

    \I__2950\ : InMux
    port map (
            O => \N__15388\,
            I => \N__15382\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__15385\,
            I => \N__15377\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__15382\,
            I => \N__15377\
        );

    \I__2947\ : Odrv12
    port map (
            O => \N__15377\,
            I => \POWERLED.dutycycle\
        );

    \I__2946\ : InMux
    port map (
            O => \N__15374\,
            I => \N__15369\
        );

    \I__2945\ : InMux
    port map (
            O => \N__15373\,
            I => \N__15364\
        );

    \I__2944\ : InMux
    port map (
            O => \N__15372\,
            I => \N__15364\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__15369\,
            I => \POWERLED.N_243\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__15364\,
            I => \POWERLED.N_243\
        );

    \I__2941\ : InMux
    port map (
            O => \N__15359\,
            I => \N__15352\
        );

    \I__2940\ : InMux
    port map (
            O => \N__15358\,
            I => \N__15347\
        );

    \I__2939\ : InMux
    port map (
            O => \N__15357\,
            I => \N__15340\
        );

    \I__2938\ : InMux
    port map (
            O => \N__15356\,
            I => \N__15340\
        );

    \I__2937\ : InMux
    port map (
            O => \N__15355\,
            I => \N__15340\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__15352\,
            I => \N__15337\
        );

    \I__2935\ : InMux
    port map (
            O => \N__15351\,
            I => \N__15334\
        );

    \I__2934\ : InMux
    port map (
            O => \N__15350\,
            I => \N__15331\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__15347\,
            I => \N__15326\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__15340\,
            I => \N__15326\
        );

    \I__2931\ : Span4Mux_h
    port map (
            O => \N__15337\,
            I => \N__15323\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__15334\,
            I => \N__15318\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__15331\,
            I => \N__15318\
        );

    \I__2928\ : Span4Mux_h
    port map (
            O => \N__15326\,
            I => \N__15315\
        );

    \I__2927\ : Sp12to4
    port map (
            O => \N__15323\,
            I => \N__15310\
        );

    \I__2926\ : Span12Mux_s8_h
    port map (
            O => \N__15318\,
            I => \N__15310\
        );

    \I__2925\ : Span4Mux_v
    port map (
            O => \N__15315\,
            I => \N__15307\
        );

    \I__2924\ : Odrv12
    port map (
            O => \N__15310\,
            I => slp_s4n
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__15307\,
            I => slp_s4n
        );

    \I__2922\ : InMux
    port map (
            O => \N__15302\,
            I => \N__15295\
        );

    \I__2921\ : InMux
    port map (
            O => \N__15301\,
            I => \N__15290\
        );

    \I__2920\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15286\
        );

    \I__2919\ : InMux
    port map (
            O => \N__15299\,
            I => \N__15283\
        );

    \I__2918\ : InMux
    port map (
            O => \N__15298\,
            I => \N__15279\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__15295\,
            I => \N__15276\
        );

    \I__2916\ : InMux
    port map (
            O => \N__15294\,
            I => \N__15273\
        );

    \I__2915\ : InMux
    port map (
            O => \N__15293\,
            I => \N__15270\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__15290\,
            I => \N__15267\
        );

    \I__2913\ : InMux
    port map (
            O => \N__15289\,
            I => \N__15264\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__15286\,
            I => \N__15259\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__15283\,
            I => \N__15259\
        );

    \I__2910\ : InMux
    port map (
            O => \N__15282\,
            I => \N__15255\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__15279\,
            I => \N__15252\
        );

    \I__2908\ : Span4Mux_v
    port map (
            O => \N__15276\,
            I => \N__15241\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__15273\,
            I => \N__15241\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__15270\,
            I => \N__15241\
        );

    \I__2905\ : Span4Mux_v
    port map (
            O => \N__15267\,
            I => \N__15241\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__15264\,
            I => \N__15241\
        );

    \I__2903\ : Span4Mux_h
    port map (
            O => \N__15259\,
            I => \N__15238\
        );

    \I__2902\ : InMux
    port map (
            O => \N__15258\,
            I => \N__15235\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__15255\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__15252\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__2899\ : Odrv4
    port map (
            O => \N__15241\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__15238\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__15235\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__15224\,
            I => \N__15217\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__15223\,
            I => \N__15213\
        );

    \I__2894\ : InMux
    port map (
            O => \N__15222\,
            I => \N__15205\
        );

    \I__2893\ : InMux
    port map (
            O => \N__15221\,
            I => \N__15202\
        );

    \I__2892\ : InMux
    port map (
            O => \N__15220\,
            I => \N__15199\
        );

    \I__2891\ : InMux
    port map (
            O => \N__15217\,
            I => \N__15190\
        );

    \I__2890\ : InMux
    port map (
            O => \N__15216\,
            I => \N__15190\
        );

    \I__2889\ : InMux
    port map (
            O => \N__15213\,
            I => \N__15190\
        );

    \I__2888\ : InMux
    port map (
            O => \N__15212\,
            I => \N__15190\
        );

    \I__2887\ : InMux
    port map (
            O => \N__15211\,
            I => \N__15185\
        );

    \I__2886\ : InMux
    port map (
            O => \N__15210\,
            I => \N__15185\
        );

    \I__2885\ : InMux
    port map (
            O => \N__15209\,
            I => \N__15180\
        );

    \I__2884\ : InMux
    port map (
            O => \N__15208\,
            I => \N__15180\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__15205\,
            I => \N__15171\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__15202\,
            I => \N__15171\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__15199\,
            I => \N__15171\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__15190\,
            I => \N__15171\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__15185\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__15180\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__15171\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__2876\ : InMux
    port map (
            O => \N__15164\,
            I => \N__15158\
        );

    \I__2875\ : InMux
    port map (
            O => \N__15163\,
            I => \N__15152\
        );

    \I__2874\ : InMux
    port map (
            O => \N__15162\,
            I => \N__15152\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__15161\,
            I => \N__15149\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__15158\,
            I => \N__15144\
        );

    \I__2871\ : InMux
    port map (
            O => \N__15157\,
            I => \N__15141\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__15152\,
            I => \N__15138\
        );

    \I__2869\ : InMux
    port map (
            O => \N__15149\,
            I => \N__15134\
        );

    \I__2868\ : InMux
    port map (
            O => \N__15148\,
            I => \N__15131\
        );

    \I__2867\ : InMux
    port map (
            O => \N__15147\,
            I => \N__15128\
        );

    \I__2866\ : Span4Mux_v
    port map (
            O => \N__15144\,
            I => \N__15123\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__15141\,
            I => \N__15123\
        );

    \I__2864\ : Span4Mux_h
    port map (
            O => \N__15138\,
            I => \N__15120\
        );

    \I__2863\ : InMux
    port map (
            O => \N__15137\,
            I => \N__15117\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__15134\,
            I => \POWERLED.count_off_RNIIKVR3Z0Z_10\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__15131\,
            I => \POWERLED.count_off_RNIIKVR3Z0Z_10\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__15128\,
            I => \POWERLED.count_off_RNIIKVR3Z0Z_10\
        );

    \I__2859\ : Odrv4
    port map (
            O => \N__15123\,
            I => \POWERLED.count_off_RNIIKVR3Z0Z_10\
        );

    \I__2858\ : Odrv4
    port map (
            O => \N__15120\,
            I => \POWERLED.count_off_RNIIKVR3Z0Z_10\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__15117\,
            I => \POWERLED.count_off_RNIIKVR3Z0Z_10\
        );

    \I__2856\ : InMux
    port map (
            O => \N__15104\,
            I => \N__15101\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__15101\,
            I => \POWERLED.N_148\
        );

    \I__2854\ : InMux
    port map (
            O => \N__15098\,
            I => \N__15094\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__15097\,
            I => \N__15087\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__15094\,
            I => \N__15080\
        );

    \I__2851\ : InMux
    port map (
            O => \N__15093\,
            I => \N__15077\
        );

    \I__2850\ : InMux
    port map (
            O => \N__15092\,
            I => \N__15070\
        );

    \I__2849\ : InMux
    port map (
            O => \N__15091\,
            I => \N__15070\
        );

    \I__2848\ : InMux
    port map (
            O => \N__15090\,
            I => \N__15070\
        );

    \I__2847\ : InMux
    port map (
            O => \N__15087\,
            I => \N__15065\
        );

    \I__2846\ : InMux
    port map (
            O => \N__15086\,
            I => \N__15065\
        );

    \I__2845\ : InMux
    port map (
            O => \N__15085\,
            I => \N__15058\
        );

    \I__2844\ : InMux
    port map (
            O => \N__15084\,
            I => \N__15058\
        );

    \I__2843\ : InMux
    port map (
            O => \N__15083\,
            I => \N__15058\
        );

    \I__2842\ : Span4Mux_h
    port map (
            O => \N__15080\,
            I => \N__15050\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__15077\,
            I => \N__15050\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__15070\,
            I => \N__15050\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__15065\,
            I => \N__15047\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__15058\,
            I => \N__15044\
        );

    \I__2837\ : InMux
    port map (
            O => \N__15057\,
            I => \N__15041\
        );

    \I__2836\ : Span4Mux_v
    port map (
            O => \N__15050\,
            I => \N__15038\
        );

    \I__2835\ : Span4Mux_v
    port map (
            O => \N__15047\,
            I => \N__15031\
        );

    \I__2834\ : Span4Mux_v
    port map (
            O => \N__15044\,
            I => \N__15031\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__15041\,
            I => \N__15031\
        );

    \I__2832\ : Span4Mux_h
    port map (
            O => \N__15038\,
            I => \N__15026\
        );

    \I__2831\ : Span4Mux_h
    port map (
            O => \N__15031\,
            I => \N__15026\
        );

    \I__2830\ : Odrv4
    port map (
            O => \N__15026\,
            I => slp_s3n
        );

    \I__2829\ : IoInMux
    port map (
            O => \N__15023\,
            I => \N__15020\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__15020\,
            I => \N__15016\
        );

    \I__2827\ : InMux
    port map (
            O => \N__15019\,
            I => \N__15013\
        );

    \I__2826\ : Span4Mux_s2_h
    port map (
            O => \N__15016\,
            I => \N__15007\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__15013\,
            I => \N__15004\
        );

    \I__2824\ : InMux
    port map (
            O => \N__15012\,
            I => \N__14999\
        );

    \I__2823\ : InMux
    port map (
            O => \N__15011\,
            I => \N__14994\
        );

    \I__2822\ : InMux
    port map (
            O => \N__15010\,
            I => \N__14994\
        );

    \I__2821\ : Span4Mux_h
    port map (
            O => \N__15007\,
            I => \N__14991\
        );

    \I__2820\ : Span4Mux_v
    port map (
            O => \N__15004\,
            I => \N__14988\
        );

    \I__2819\ : InMux
    port map (
            O => \N__15003\,
            I => \N__14983\
        );

    \I__2818\ : InMux
    port map (
            O => \N__15002\,
            I => \N__14983\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__14999\,
            I => \N__14978\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__14994\,
            I => \N__14978\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__14991\,
            I => vccst_en
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__14988\,
            I => vccst_en
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__14983\,
            I => vccst_en
        );

    \I__2812\ : Odrv4
    port map (
            O => \N__14978\,
            I => vccst_en
        );

    \I__2811\ : IoInMux
    port map (
            O => \N__14969\,
            I => \N__14966\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__14966\,
            I => \N__14963\
        );

    \I__2809\ : Odrv12
    port map (
            O => \N__14963\,
            I => vpp_en
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__14960\,
            I => \POWERLED.N_203_cascade_\
        );

    \I__2807\ : CascadeMux
    port map (
            O => \N__14957\,
            I => \POWERLED.N_251_cascade_\
        );

    \I__2806\ : InMux
    port map (
            O => \N__14954\,
            I => \N__14951\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__14951\,
            I => \POWERLED.un2_slp_s3n_2_0_1_0\
        );

    \I__2804\ : InMux
    port map (
            O => \N__14948\,
            I => \N__14945\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__14945\,
            I => \POWERLED.count_clk_139_tz_0\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__14942\,
            I => \POWERLED.un2_slp_s3n_2_0_cascade_\
        );

    \I__2801\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14936\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__14936\,
            I => \POWERLED.N_246\
        );

    \I__2799\ : InMux
    port map (
            O => \N__14933\,
            I => \N__14930\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__14930\,
            I => \N__14927\
        );

    \I__2797\ : Span4Mux_h
    port map (
            O => \N__14927\,
            I => \N__14923\
        );

    \I__2796\ : InMux
    port map (
            O => \N__14926\,
            I => \N__14920\
        );

    \I__2795\ : Odrv4
    port map (
            O => \N__14923\,
            I => \POWERLED.N_205\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__14920\,
            I => \POWERLED.N_205\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__14915\,
            I => \POWERLED.un2_slp_s3n_2_0_a6_3_0_cascade_\
        );

    \I__2792\ : InMux
    port map (
            O => \N__14912\,
            I => \N__14909\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__14909\,
            I => \POWERLED.un2_slp_s3n_2_0_1\
        );

    \I__2790\ : InMux
    port map (
            O => \N__14906\,
            I => \N__14903\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__14903\,
            I => \N__14898\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__14902\,
            I => \N__14894\
        );

    \I__2787\ : InMux
    port map (
            O => \N__14901\,
            I => \N__14891\
        );

    \I__2786\ : Span4Mux_h
    port map (
            O => \N__14898\,
            I => \N__14888\
        );

    \I__2785\ : InMux
    port map (
            O => \N__14897\,
            I => \N__14885\
        );

    \I__2784\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14882\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__14891\,
            I => \N__14879\
        );

    \I__2782\ : Odrv4
    port map (
            O => \N__14888\,
            I => \POWERLED.N_127\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__14885\,
            I => \POWERLED.N_127\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__14882\,
            I => \POWERLED.N_127\
        );

    \I__2779\ : Odrv4
    port map (
            O => \N__14879\,
            I => \POWERLED.N_127\
        );

    \I__2778\ : InMux
    port map (
            O => \N__14870\,
            I => \POWERLED.dutycycle_cry_9\
        );

    \I__2777\ : InMux
    port map (
            O => \N__14867\,
            I => \POWERLED.dutycycle_cry_10\
        );

    \I__2776\ : InMux
    port map (
            O => \N__14864\,
            I => \POWERLED.dutycycle_cry_11\
        );

    \I__2775\ : InMux
    port map (
            O => \N__14861\,
            I => \POWERLED.dutycycle_cry_12\
        );

    \I__2774\ : InMux
    port map (
            O => \N__14858\,
            I => \POWERLED.dutycycle_cry_13\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__14855\,
            I => \N__14845\
        );

    \I__2772\ : CascadeMux
    port map (
            O => \N__14854\,
            I => \N__14841\
        );

    \I__2771\ : CascadeMux
    port map (
            O => \N__14853\,
            I => \N__14837\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__14852\,
            I => \N__14833\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__14851\,
            I => \N__14829\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__14850\,
            I => \N__14825\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__14849\,
            I => \N__14821\
        );

    \I__2766\ : InMux
    port map (
            O => \N__14848\,
            I => \N__14805\
        );

    \I__2765\ : InMux
    port map (
            O => \N__14845\,
            I => \N__14805\
        );

    \I__2764\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14805\
        );

    \I__2763\ : InMux
    port map (
            O => \N__14841\,
            I => \N__14805\
        );

    \I__2762\ : InMux
    port map (
            O => \N__14840\,
            I => \N__14805\
        );

    \I__2761\ : InMux
    port map (
            O => \N__14837\,
            I => \N__14805\
        );

    \I__2760\ : InMux
    port map (
            O => \N__14836\,
            I => \N__14805\
        );

    \I__2759\ : InMux
    port map (
            O => \N__14833\,
            I => \N__14787\
        );

    \I__2758\ : InMux
    port map (
            O => \N__14832\,
            I => \N__14787\
        );

    \I__2757\ : InMux
    port map (
            O => \N__14829\,
            I => \N__14787\
        );

    \I__2756\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14787\
        );

    \I__2755\ : InMux
    port map (
            O => \N__14825\,
            I => \N__14787\
        );

    \I__2754\ : InMux
    port map (
            O => \N__14824\,
            I => \N__14787\
        );

    \I__2753\ : InMux
    port map (
            O => \N__14821\,
            I => \N__14787\
        );

    \I__2752\ : InMux
    port map (
            O => \N__14820\,
            I => \N__14787\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__14805\,
            I => \N__14784\
        );

    \I__2750\ : InMux
    port map (
            O => \N__14804\,
            I => \N__14781\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__14787\,
            I => \N__14778\
        );

    \I__2748\ : Span4Mux_h
    port map (
            O => \N__14784\,
            I => \N__14775\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__14781\,
            I => \POWERLED.N_177\
        );

    \I__2746\ : Odrv4
    port map (
            O => \N__14778\,
            I => \POWERLED.N_177\
        );

    \I__2745\ : Odrv4
    port map (
            O => \N__14775\,
            I => \POWERLED.N_177\
        );

    \I__2744\ : InMux
    port map (
            O => \N__14768\,
            I => \bfn_7_9_0_\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__14765\,
            I => \POWERLED.N_246_cascade_\
        );

    \I__2742\ : InMux
    port map (
            O => \N__14762\,
            I => \N__14759\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__14759\,
            I => \POWERLED.N_203_4\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__14756\,
            I => \POWERLED.N_203_4_cascade_\
        );

    \I__2739\ : InMux
    port map (
            O => \N__14753\,
            I => \N__14748\
        );

    \I__2738\ : InMux
    port map (
            O => \N__14752\,
            I => \N__14745\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__14751\,
            I => \N__14742\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__14748\,
            I => \N__14737\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__14745\,
            I => \N__14733\
        );

    \I__2734\ : InMux
    port map (
            O => \N__14742\,
            I => \N__14730\
        );

    \I__2733\ : CascadeMux
    port map (
            O => \N__14741\,
            I => \N__14727\
        );

    \I__2732\ : CascadeMux
    port map (
            O => \N__14740\,
            I => \N__14723\
        );

    \I__2731\ : Span4Mux_v
    port map (
            O => \N__14737\,
            I => \N__14719\
        );

    \I__2730\ : InMux
    port map (
            O => \N__14736\,
            I => \N__14716\
        );

    \I__2729\ : Span4Mux_v
    port map (
            O => \N__14733\,
            I => \N__14713\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__14730\,
            I => \N__14710\
        );

    \I__2727\ : InMux
    port map (
            O => \N__14727\,
            I => \N__14707\
        );

    \I__2726\ : InMux
    port map (
            O => \N__14726\,
            I => \N__14704\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14723\,
            I => \N__14701\
        );

    \I__2724\ : InMux
    port map (
            O => \N__14722\,
            I => \N__14698\
        );

    \I__2723\ : Span4Mux_v
    port map (
            O => \N__14719\,
            I => \N__14693\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__14716\,
            I => \N__14693\
        );

    \I__2721\ : Span4Mux_h
    port map (
            O => \N__14713\,
            I => \N__14688\
        );

    \I__2720\ : Span4Mux_h
    port map (
            O => \N__14710\,
            I => \N__14688\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__14707\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__14704\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__14701\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__14698\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__2715\ : Odrv4
    port map (
            O => \N__14693\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__2714\ : Odrv4
    port map (
            O => \N__14688\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__2713\ : InMux
    port map (
            O => \N__14675\,
            I => \N__14672\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__14672\,
            I => \POWERLED.dutycycle_s_2\
        );

    \I__2711\ : InMux
    port map (
            O => \N__14669\,
            I => \POWERLED.dutycycle_cry_1\
        );

    \I__2710\ : InMux
    port map (
            O => \N__14666\,
            I => \N__14662\
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__14665\,
            I => \N__14659\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__14662\,
            I => \N__14655\
        );

    \I__2707\ : InMux
    port map (
            O => \N__14659\,
            I => \N__14651\
        );

    \I__2706\ : InMux
    port map (
            O => \N__14658\,
            I => \N__14648\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__14655\,
            I => \N__14641\
        );

    \I__2704\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14638\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__14651\,
            I => \N__14633\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__14648\,
            I => \N__14633\
        );

    \I__2701\ : InMux
    port map (
            O => \N__14647\,
            I => \N__14630\
        );

    \I__2700\ : InMux
    port map (
            O => \N__14646\,
            I => \N__14625\
        );

    \I__2699\ : InMux
    port map (
            O => \N__14645\,
            I => \N__14625\
        );

    \I__2698\ : InMux
    port map (
            O => \N__14644\,
            I => \N__14622\
        );

    \I__2697\ : Odrv4
    port map (
            O => \N__14641\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__14638\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__14633\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__14630\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__14625\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__14622\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__2691\ : InMux
    port map (
            O => \N__14609\,
            I => \POWERLED.dutycycle_cry_2\
        );

    \I__2690\ : InMux
    port map (
            O => \N__14606\,
            I => \N__14598\
        );

    \I__2689\ : InMux
    port map (
            O => \N__14605\,
            I => \N__14593\
        );

    \I__2688\ : InMux
    port map (
            O => \N__14604\,
            I => \N__14593\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__14603\,
            I => \N__14590\
        );

    \I__2686\ : InMux
    port map (
            O => \N__14602\,
            I => \N__14587\
        );

    \I__2685\ : InMux
    port map (
            O => \N__14601\,
            I => \N__14582\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__14598\,
            I => \N__14579\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__14593\,
            I => \N__14576\
        );

    \I__2682\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14573\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__14587\,
            I => \N__14570\
        );

    \I__2680\ : InMux
    port map (
            O => \N__14586\,
            I => \N__14565\
        );

    \I__2679\ : InMux
    port map (
            O => \N__14585\,
            I => \N__14565\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__14582\,
            I => \N__14560\
        );

    \I__2677\ : Span4Mux_h
    port map (
            O => \N__14579\,
            I => \N__14560\
        );

    \I__2676\ : Span4Mux_h
    port map (
            O => \N__14576\,
            I => \N__14557\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__14573\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__2674\ : Odrv4
    port map (
            O => \N__14570\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__14565\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__2672\ : Odrv4
    port map (
            O => \N__14560\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__2671\ : Odrv4
    port map (
            O => \N__14557\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__2670\ : InMux
    port map (
            O => \N__14546\,
            I => \POWERLED.dutycycle_cry_3\
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__14543\,
            I => \N__14539\
        );

    \I__2668\ : InMux
    port map (
            O => \N__14542\,
            I => \N__14536\
        );

    \I__2667\ : InMux
    port map (
            O => \N__14539\,
            I => \N__14533\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__14536\,
            I => \N__14527\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__14533\,
            I => \N__14524\
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__14532\,
            I => \N__14520\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__14531\,
            I => \N__14517\
        );

    \I__2662\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14514\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__14527\,
            I => \N__14511\
        );

    \I__2660\ : Span4Mux_h
    port map (
            O => \N__14524\,
            I => \N__14508\
        );

    \I__2659\ : InMux
    port map (
            O => \N__14523\,
            I => \N__14505\
        );

    \I__2658\ : InMux
    port map (
            O => \N__14520\,
            I => \N__14500\
        );

    \I__2657\ : InMux
    port map (
            O => \N__14517\,
            I => \N__14500\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__14514\,
            I => \N__14497\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__14511\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__2654\ : Odrv4
    port map (
            O => \N__14508\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__14505\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__14500\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__2651\ : Odrv4
    port map (
            O => \N__14497\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__2650\ : InMux
    port map (
            O => \N__14486\,
            I => \N__14482\
        );

    \I__2649\ : InMux
    port map (
            O => \N__14485\,
            I => \N__14479\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__14482\,
            I => \N__14476\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__14479\,
            I => \N__14473\
        );

    \I__2646\ : Span4Mux_h
    port map (
            O => \N__14476\,
            I => \N__14470\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__14473\,
            I => \N__14467\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__14470\,
            I => \POWERLED.dutycycle_s_5\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__14467\,
            I => \POWERLED.dutycycle_s_5\
        );

    \I__2642\ : InMux
    port map (
            O => \N__14462\,
            I => \POWERLED.dutycycle_cry_4\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__14459\,
            I => \N__14456\
        );

    \I__2640\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14451\
        );

    \I__2639\ : InMux
    port map (
            O => \N__14455\,
            I => \N__14446\
        );

    \I__2638\ : InMux
    port map (
            O => \N__14454\,
            I => \N__14446\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__14451\,
            I => \N__14437\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__14446\,
            I => \N__14437\
        );

    \I__2635\ : InMux
    port map (
            O => \N__14445\,
            I => \N__14434\
        );

    \I__2634\ : InMux
    port map (
            O => \N__14444\,
            I => \N__14427\
        );

    \I__2633\ : InMux
    port map (
            O => \N__14443\,
            I => \N__14427\
        );

    \I__2632\ : InMux
    port map (
            O => \N__14442\,
            I => \N__14427\
        );

    \I__2631\ : Span4Mux_v
    port map (
            O => \N__14437\,
            I => \N__14424\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__14434\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__14427\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__14424\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__2627\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14411\
        );

    \I__2626\ : InMux
    port map (
            O => \N__14416\,
            I => \N__14411\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__14411\,
            I => \N__14408\
        );

    \I__2624\ : Span4Mux_h
    port map (
            O => \N__14408\,
            I => \N__14405\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__14405\,
            I => \POWERLED.dutycycle_s_6\
        );

    \I__2622\ : InMux
    port map (
            O => \N__14402\,
            I => \POWERLED.dutycycle_cry_5\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__14399\,
            I => \N__14389\
        );

    \I__2620\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14386\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__14397\,
            I => \N__14382\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__14396\,
            I => \N__14379\
        );

    \I__2617\ : InMux
    port map (
            O => \N__14395\,
            I => \N__14374\
        );

    \I__2616\ : InMux
    port map (
            O => \N__14394\,
            I => \N__14374\
        );

    \I__2615\ : InMux
    port map (
            O => \N__14393\,
            I => \N__14370\
        );

    \I__2614\ : InMux
    port map (
            O => \N__14392\,
            I => \N__14365\
        );

    \I__2613\ : InMux
    port map (
            O => \N__14389\,
            I => \N__14365\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__14386\,
            I => \N__14362\
        );

    \I__2611\ : InMux
    port map (
            O => \N__14385\,
            I => \N__14357\
        );

    \I__2610\ : InMux
    port map (
            O => \N__14382\,
            I => \N__14357\
        );

    \I__2609\ : InMux
    port map (
            O => \N__14379\,
            I => \N__14354\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__14374\,
            I => \N__14351\
        );

    \I__2607\ : InMux
    port map (
            O => \N__14373\,
            I => \N__14348\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__14370\,
            I => \N__14343\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__14365\,
            I => \N__14343\
        );

    \I__2604\ : Span4Mux_v
    port map (
            O => \N__14362\,
            I => \N__14338\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__14357\,
            I => \N__14338\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__14354\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__2601\ : Odrv4
    port map (
            O => \N__14351\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__14348\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__2599\ : Odrv4
    port map (
            O => \N__14343\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__14338\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__2597\ : InMux
    port map (
            O => \N__14327\,
            I => \bfn_7_8_0_\
        );

    \I__2596\ : InMux
    port map (
            O => \N__14324\,
            I => \POWERLED.dutycycle_cry_7\
        );

    \I__2595\ : InMux
    port map (
            O => \N__14321\,
            I => \POWERLED.dutycycle_cry_8\
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__14318\,
            I => \POWERLED.un1_dutycycle_1_39_0_cascade_\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__14315\,
            I => \N__14312\
        );

    \I__2592\ : InMux
    port map (
            O => \N__14312\,
            I => \N__14309\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__14309\,
            I => \POWERLED.dutycycle_RNI34C41Z0Z_8\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__14306\,
            I => \N__14301\
        );

    \I__2589\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14296\
        );

    \I__2588\ : InMux
    port map (
            O => \N__14304\,
            I => \N__14296\
        );

    \I__2587\ : InMux
    port map (
            O => \N__14301\,
            I => \N__14293\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__14296\,
            I => \N__14290\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__14293\,
            I => \N__14285\
        );

    \I__2584\ : Span4Mux_h
    port map (
            O => \N__14290\,
            I => \N__14285\
        );

    \I__2583\ : Span4Mux_v
    port map (
            O => \N__14285\,
            I => \N__14282\
        );

    \I__2582\ : Odrv4
    port map (
            O => \N__14282\,
            I => \POWERLED.N_117\
        );

    \I__2581\ : InMux
    port map (
            O => \N__14279\,
            I => \N__14275\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__14278\,
            I => \N__14272\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__14275\,
            I => \N__14269\
        );

    \I__2578\ : InMux
    port map (
            O => \N__14272\,
            I => \N__14266\
        );

    \I__2577\ : Odrv12
    port map (
            O => \N__14269\,
            I => \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__14266\,
            I => \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5\
        );

    \I__2575\ : InMux
    port map (
            O => \N__14261\,
            I => \N__14258\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__14258\,
            I => \POWERLED.dutycycle_RNIK4I81Z0Z_6\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__14255\,
            I => \N__14252\
        );

    \I__2572\ : InMux
    port map (
            O => \N__14252\,
            I => \N__14249\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__14249\,
            I => \N__14246\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__14246\,
            I => \POWERLED.dutycycle_lm_0_1_2\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__14243\,
            I => \N__14240\
        );

    \I__2568\ : InMux
    port map (
            O => \N__14240\,
            I => \N__14236\
        );

    \I__2567\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14233\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__14236\,
            I => \N__14230\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__14233\,
            I => \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6\
        );

    \I__2564\ : Odrv4
    port map (
            O => \N__14230\,
            I => \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6\
        );

    \I__2563\ : InMux
    port map (
            O => \N__14225\,
            I => \N__14222\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__14222\,
            I => \POWERLED.dutycycle_RNIQAI81Z0Z_4\
        );

    \I__2561\ : InMux
    port map (
            O => \N__14219\,
            I => \N__14216\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__14216\,
            I => \POWERLED.dutycycle_RNIOQLJZ0Z_4\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__14213\,
            I => \N__14210\
        );

    \I__2558\ : InMux
    port map (
            O => \N__14210\,
            I => \N__14206\
        );

    \I__2557\ : InMux
    port map (
            O => \N__14209\,
            I => \N__14203\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__14206\,
            I => \N__14200\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__14203\,
            I => \N__14197\
        );

    \I__2554\ : Span4Mux_v
    port map (
            O => \N__14200\,
            I => \N__14191\
        );

    \I__2553\ : Span4Mux_h
    port map (
            O => \N__14197\,
            I => \N__14188\
        );

    \I__2552\ : InMux
    port map (
            O => \N__14196\,
            I => \N__14185\
        );

    \I__2551\ : InMux
    port map (
            O => \N__14195\,
            I => \N__14182\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__14194\,
            I => \N__14179\
        );

    \I__2549\ : Span4Mux_h
    port map (
            O => \N__14191\,
            I => \N__14174\
        );

    \I__2548\ : Span4Mux_v
    port map (
            O => \N__14188\,
            I => \N__14169\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__14185\,
            I => \N__14169\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__14182\,
            I => \N__14166\
        );

    \I__2545\ : InMux
    port map (
            O => \N__14179\,
            I => \N__14163\
        );

    \I__2544\ : InMux
    port map (
            O => \N__14178\,
            I => \N__14160\
        );

    \I__2543\ : InMux
    port map (
            O => \N__14177\,
            I => \N__14157\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__14174\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__14169\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__14166\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__14163\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__14160\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__14157\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__2536\ : InMux
    port map (
            O => \N__14144\,
            I => \N__14141\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__14141\,
            I => \N__14138\
        );

    \I__2534\ : Span4Mux_v
    port map (
            O => \N__14138\,
            I => \N__14135\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__14135\,
            I => \POWERLED.dutycycle_s_0\
        );

    \I__2532\ : InMux
    port map (
            O => \N__14132\,
            I => \POWERLED.dutycycle_cry_c_0_THRU_CO\
        );

    \I__2531\ : InMux
    port map (
            O => \N__14129\,
            I => \N__14124\
        );

    \I__2530\ : InMux
    port map (
            O => \N__14128\,
            I => \N__14120\
        );

    \I__2529\ : InMux
    port map (
            O => \N__14127\,
            I => \N__14116\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__14124\,
            I => \N__14113\
        );

    \I__2527\ : InMux
    port map (
            O => \N__14123\,
            I => \N__14107\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__14120\,
            I => \N__14104\
        );

    \I__2525\ : InMux
    port map (
            O => \N__14119\,
            I => \N__14101\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__14116\,
            I => \N__14098\
        );

    \I__2523\ : Span4Mux_v
    port map (
            O => \N__14113\,
            I => \N__14095\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__14112\,
            I => \N__14092\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__14111\,
            I => \N__14089\
        );

    \I__2520\ : CascadeMux
    port map (
            O => \N__14110\,
            I => \N__14085\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__14107\,
            I => \N__14082\
        );

    \I__2518\ : Span4Mux_v
    port map (
            O => \N__14104\,
            I => \N__14077\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__14101\,
            I => \N__14077\
        );

    \I__2516\ : Span4Mux_v
    port map (
            O => \N__14098\,
            I => \N__14072\
        );

    \I__2515\ : Span4Mux_h
    port map (
            O => \N__14095\,
            I => \N__14072\
        );

    \I__2514\ : InMux
    port map (
            O => \N__14092\,
            I => \N__14067\
        );

    \I__2513\ : InMux
    port map (
            O => \N__14089\,
            I => \N__14067\
        );

    \I__2512\ : InMux
    port map (
            O => \N__14088\,
            I => \N__14062\
        );

    \I__2511\ : InMux
    port map (
            O => \N__14085\,
            I => \N__14062\
        );

    \I__2510\ : Odrv12
    port map (
            O => \N__14082\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__2509\ : Odrv4
    port map (
            O => \N__14077\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__2508\ : Odrv4
    port map (
            O => \N__14072\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__14067\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__14062\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__2505\ : InMux
    port map (
            O => \N__14051\,
            I => \N__14048\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__14048\,
            I => \N__14045\
        );

    \I__2503\ : Span4Mux_h
    port map (
            O => \N__14045\,
            I => \N__14042\
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__14042\,
            I => \POWERLED.dutycycle_s_1\
        );

    \I__2501\ : InMux
    port map (
            O => \N__14039\,
            I => \POWERLED.dutycycle_cry_0\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__14036\,
            I => \N__14033\
        );

    \I__2499\ : InMux
    port map (
            O => \N__14033\,
            I => \N__14030\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__14030\,
            I => \N__14027\
        );

    \I__2497\ : Odrv12
    port map (
            O => \N__14027\,
            I => \HDA_STRAP.curr_state_RNO_0Z0Z_2\
        );

    \I__2496\ : CascadeMux
    port map (
            O => \N__14024\,
            I => \N__14021\
        );

    \I__2495\ : InMux
    port map (
            O => \N__14021\,
            I => \N__14018\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__14018\,
            I => \HDA_STRAP.count_RNO_0Z0Z_10\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__14015\,
            I => \N__14012\
        );

    \I__2492\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14008\
        );

    \I__2491\ : InMux
    port map (
            O => \N__14011\,
            I => \N__14005\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__14008\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__14005\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__2488\ : InMux
    port map (
            O => \N__14000\,
            I => \N__13997\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__13997\,
            I => \HDA_STRAP.count_RNO_0Z0Z_16\
        );

    \I__2486\ : InMux
    port map (
            O => \N__13994\,
            I => \N__13990\
        );

    \I__2485\ : InMux
    port map (
            O => \N__13993\,
            I => \N__13987\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__13990\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__13987\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__2482\ : InMux
    port map (
            O => \N__13982\,
            I => \N__13979\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__13979\,
            I => \HDA_STRAP.count_RNO_0Z0Z_17\
        );

    \I__2480\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13972\
        );

    \I__2479\ : InMux
    port map (
            O => \N__13975\,
            I => \N__13969\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__13972\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__13969\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__2476\ : InMux
    port map (
            O => \N__13964\,
            I => \N__13961\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__13961\,
            I => \HDA_STRAP.count_RNO_0Z0Z_8\
        );

    \I__2474\ : InMux
    port map (
            O => \N__13958\,
            I => \N__13954\
        );

    \I__2473\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13951\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__13954\,
            I => \HDA_STRAP.countZ0Z_8\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__13951\,
            I => \HDA_STRAP.countZ0Z_8\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__13946\,
            I => \N__13943\
        );

    \I__2469\ : InMux
    port map (
            O => \N__13943\,
            I => \N__13940\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__13940\,
            I => \POWERLED.dutycycle_RNI31MG_0Z0Z_12\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__13937\,
            I => \N__13934\
        );

    \I__2466\ : InMux
    port map (
            O => \N__13934\,
            I => \N__13931\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__13931\,
            I => \POWERLED.dutycycle_RNI31MGZ0Z_12\
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__13928\,
            I => \N__13924\
        );

    \I__2463\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13921\
        );

    \I__2462\ : InMux
    port map (
            O => \N__13924\,
            I => \N__13918\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__13921\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__13918\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\
        );

    \I__2459\ : InMux
    port map (
            O => \N__13913\,
            I => \N__13909\
        );

    \I__2458\ : InMux
    port map (
            O => \N__13912\,
            I => \N__13906\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__13909\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__13906\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__2455\ : InMux
    port map (
            O => \N__13901\,
            I => \N__13897\
        );

    \I__2454\ : InMux
    port map (
            O => \N__13900\,
            I => \N__13894\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__13897\,
            I => \HDA_STRAP.countZ0Z_1\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__13894\,
            I => \HDA_STRAP.countZ0Z_1\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__13889\,
            I => \N__13885\
        );

    \I__2450\ : InMux
    port map (
            O => \N__13888\,
            I => \N__13882\
        );

    \I__2449\ : InMux
    port map (
            O => \N__13885\,
            I => \N__13879\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__13882\,
            I => \HDA_STRAP.countZ0Z_3\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__13879\,
            I => \HDA_STRAP.countZ0Z_3\
        );

    \I__2446\ : InMux
    port map (
            O => \N__13874\,
            I => \N__13870\
        );

    \I__2445\ : InMux
    port map (
            O => \N__13873\,
            I => \N__13867\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__13870\,
            I => \N__13862\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__13867\,
            I => \N__13862\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__13862\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__2441\ : InMux
    port map (
            O => \N__13859\,
            I => \N__13855\
        );

    \I__2440\ : InMux
    port map (
            O => \N__13858\,
            I => \N__13852\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__13855\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__13852\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__2437\ : CascadeMux
    port map (
            O => \N__13847\,
            I => \N__13843\
        );

    \I__2436\ : InMux
    port map (
            O => \N__13846\,
            I => \N__13840\
        );

    \I__2435\ : InMux
    port map (
            O => \N__13843\,
            I => \N__13837\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__13840\,
            I => \HDA_STRAP.countZ0Z_15\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__13837\,
            I => \HDA_STRAP.countZ0Z_15\
        );

    \I__2432\ : InMux
    port map (
            O => \N__13832\,
            I => \N__13828\
        );

    \I__2431\ : InMux
    port map (
            O => \N__13831\,
            I => \N__13825\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__13828\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__13825\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__13820\,
            I => \HDA_STRAP.un4_count_9_cascade_\
        );

    \I__2427\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13813\
        );

    \I__2426\ : InMux
    port map (
            O => \N__13816\,
            I => \N__13810\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__13813\,
            I => \HDA_STRAP.countZ0Z_13\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__13810\,
            I => \HDA_STRAP.countZ0Z_13\
        );

    \I__2423\ : InMux
    port map (
            O => \N__13805\,
            I => \N__13801\
        );

    \I__2422\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13798\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__13801\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__13798\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__2419\ : InMux
    port map (
            O => \N__13793\,
            I => \N__13789\
        );

    \I__2418\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13786\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__13789\,
            I => \HDA_STRAP.countZ0Z_5\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__13786\,
            I => \HDA_STRAP.countZ0Z_5\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__13781\,
            I => \N__13777\
        );

    \I__2414\ : InMux
    port map (
            O => \N__13780\,
            I => \N__13774\
        );

    \I__2413\ : InMux
    port map (
            O => \N__13777\,
            I => \N__13771\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__13774\,
            I => \HDA_STRAP.countZ0Z_9\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__13771\,
            I => \HDA_STRAP.countZ0Z_9\
        );

    \I__2410\ : InMux
    port map (
            O => \N__13766\,
            I => \N__13762\
        );

    \I__2409\ : InMux
    port map (
            O => \N__13765\,
            I => \N__13759\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__13762\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__13759\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__2406\ : InMux
    port map (
            O => \N__13754\,
            I => \N__13750\
        );

    \I__2405\ : InMux
    port map (
            O => \N__13753\,
            I => \N__13747\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__13750\,
            I => \N__13744\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__13747\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__13744\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__2401\ : InMux
    port map (
            O => \N__13739\,
            I => \N__13736\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__13736\,
            I => \HDA_STRAP.un4_count_12\
        );

    \I__2399\ : InMux
    port map (
            O => \N__13733\,
            I => \N__13730\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__13730\,
            I => \HDA_STRAP.un4_count_11\
        );

    \I__2397\ : CascadeMux
    port map (
            O => \N__13727\,
            I => \HDA_STRAP.un4_count_10_cascade_\
        );

    \I__2396\ : InMux
    port map (
            O => \N__13724\,
            I => \N__13721\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__13721\,
            I => \HDA_STRAP.un4_count_13\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__13718\,
            I => \HDA_STRAP.count_RNIB5IA5Z0Z_0_cascade_\
        );

    \I__2393\ : CascadeMux
    port map (
            O => \N__13715\,
            I => \POWERLED.N_208_cascade_\
        );

    \I__2392\ : InMux
    port map (
            O => \N__13712\,
            I => \N__13709\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__13709\,
            I => \POWERLED.func_state_ns_i_0_1_1\
        );

    \I__2390\ : InMux
    port map (
            O => \N__13706\,
            I => \N__13703\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__13703\,
            I => \N__13695\
        );

    \I__2388\ : InMux
    port map (
            O => \N__13702\,
            I => \N__13690\
        );

    \I__2387\ : InMux
    port map (
            O => \N__13701\,
            I => \N__13690\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__13700\,
            I => \N__13687\
        );

    \I__2385\ : CascadeMux
    port map (
            O => \N__13699\,
            I => \N__13684\
        );

    \I__2384\ : InMux
    port map (
            O => \N__13698\,
            I => \N__13680\
        );

    \I__2383\ : Span4Mux_h
    port map (
            O => \N__13695\,
            I => \N__13677\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__13690\,
            I => \N__13674\
        );

    \I__2381\ : InMux
    port map (
            O => \N__13687\,
            I => \N__13667\
        );

    \I__2380\ : InMux
    port map (
            O => \N__13684\,
            I => \N__13667\
        );

    \I__2379\ : InMux
    port map (
            O => \N__13683\,
            I => \N__13667\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__13680\,
            I => \POWERLED.N_222\
        );

    \I__2377\ : Odrv4
    port map (
            O => \N__13677\,
            I => \POWERLED.N_222\
        );

    \I__2376\ : Odrv4
    port map (
            O => \N__13674\,
            I => \POWERLED.N_222\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__13667\,
            I => \POWERLED.N_222\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__13658\,
            I => \POWERLED.N_222_cascade_\
        );

    \I__2373\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13649\
        );

    \I__2372\ : InMux
    port map (
            O => \N__13654\,
            I => \N__13649\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__13649\,
            I => \POWERLED.N_228\
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__13646\,
            I => \POWERLED.N_211_cascade_\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__13643\,
            I => \N__13640\
        );

    \I__2368\ : InMux
    port map (
            O => \N__13640\,
            I => \N__13637\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__13637\,
            I => \POWERLED.func_state_ns_i_0_0_1\
        );

    \I__2366\ : InMux
    port map (
            O => \N__13634\,
            I => \N__13631\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__13631\,
            I => \POWERLED.N_179\
        );

    \I__2364\ : InMux
    port map (
            O => \N__13628\,
            I => \N__13625\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__13625\,
            I => \POWERLED.N_178\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__13622\,
            I => \N__13619\
        );

    \I__2361\ : InMux
    port map (
            O => \N__13619\,
            I => \N__13616\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__13616\,
            I => \N__13613\
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__13613\,
            I => \POWERLED.N_180\
        );

    \I__2358\ : InMux
    port map (
            O => \N__13610\,
            I => \N__13607\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__13607\,
            I => \N__13603\
        );

    \I__2356\ : InMux
    port map (
            O => \N__13606\,
            I => \N__13600\
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__13603\,
            I => \POWERLED.N_250\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__13600\,
            I => \POWERLED.N_250\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__13595\,
            I => \N__13590\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__13594\,
            I => \N__13587\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__13593\,
            I => \N__13583\
        );

    \I__2350\ : InMux
    port map (
            O => \N__13590\,
            I => \N__13576\
        );

    \I__2349\ : InMux
    port map (
            O => \N__13587\,
            I => \N__13576\
        );

    \I__2348\ : InMux
    port map (
            O => \N__13586\,
            I => \N__13576\
        );

    \I__2347\ : InMux
    port map (
            O => \N__13583\,
            I => \N__13573\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__13576\,
            I => \N__13570\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__13573\,
            I => \N__13567\
        );

    \I__2344\ : Span4Mux_h
    port map (
            O => \N__13570\,
            I => \N__13564\
        );

    \I__2343\ : Span4Mux_v
    port map (
            O => \N__13567\,
            I => \N__13561\
        );

    \I__2342\ : Odrv4
    port map (
            O => \N__13564\,
            I => \POWERLED.N_213\
        );

    \I__2341\ : Odrv4
    port map (
            O => \N__13561\,
            I => \POWERLED.N_213\
        );

    \I__2340\ : InMux
    port map (
            O => \N__13556\,
            I => \N__13550\
        );

    \I__2339\ : InMux
    port map (
            O => \N__13555\,
            I => \N__13550\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__13550\,
            I => \N__13545\
        );

    \I__2337\ : InMux
    port map (
            O => \N__13549\,
            I => \N__13540\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13548\,
            I => \N__13540\
        );

    \I__2335\ : Span4Mux_v
    port map (
            O => \N__13545\,
            I => \N__13535\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__13540\,
            I => \N__13535\
        );

    \I__2333\ : Odrv4
    port map (
            O => \N__13535\,
            I => \POWERLED.N_234\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__13532\,
            I => \POWERLED.N_218_cascade_\
        );

    \I__2331\ : InMux
    port map (
            O => \N__13529\,
            I => \N__13525\
        );

    \I__2330\ : InMux
    port map (
            O => \N__13528\,
            I => \N__13522\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__13525\,
            I => \N__13518\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__13522\,
            I => \N__13514\
        );

    \I__2327\ : InMux
    port map (
            O => \N__13521\,
            I => \N__13511\
        );

    \I__2326\ : Span4Mux_v
    port map (
            O => \N__13518\,
            I => \N__13508\
        );

    \I__2325\ : InMux
    port map (
            O => \N__13517\,
            I => \N__13505\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__13514\,
            I => \POWERLED.N_248\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__13511\,
            I => \POWERLED.N_248\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__13508\,
            I => \POWERLED.N_248\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__13505\,
            I => \POWERLED.N_248\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__13496\,
            I => \POWERLED.N_88_cascade_\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__13493\,
            I => \N__13490\
        );

    \I__2318\ : InMux
    port map (
            O => \N__13490\,
            I => \N__13487\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__13487\,
            I => \N__13484\
        );

    \I__2316\ : Odrv12
    port map (
            O => \N__13484\,
            I => \POWERLED.dutycycle_RNIC8C11Z0Z_15\
        );

    \I__2315\ : InMux
    port map (
            O => \N__13481\,
            I => \N__13478\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__13478\,
            I => \N__13475\
        );

    \I__2313\ : Span4Mux_h
    port map (
            O => \N__13475\,
            I => \N__13472\
        );

    \I__2312\ : Odrv4
    port map (
            O => \N__13472\,
            I => \POWERLED.dutycycle_RNI73C11Z0Z_15\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__13469\,
            I => \N__13466\
        );

    \I__2310\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13463\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__13463\,
            I => \POWERLED.N_368_0_i_i_a6_0\
        );

    \I__2308\ : CascadeMux
    port map (
            O => \N__13460\,
            I => \POWERLED.N_207_cascade_\
        );

    \I__2307\ : CascadeMux
    port map (
            O => \N__13457\,
            I => \N__13453\
        );

    \I__2306\ : InMux
    port map (
            O => \N__13456\,
            I => \N__13450\
        );

    \I__2305\ : InMux
    port map (
            O => \N__13453\,
            I => \N__13447\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__13450\,
            I => \POWERLED.N_48\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__13447\,
            I => \POWERLED.N_48\
        );

    \I__2302\ : CascadeMux
    port map (
            O => \N__13442\,
            I => \N__13439\
        );

    \I__2301\ : InMux
    port map (
            O => \N__13439\,
            I => \N__13436\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__13436\,
            I => \POWERLED.N_149\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__13433\,
            I => \POWERLED.N_149_cascade_\
        );

    \I__2298\ : InMux
    port map (
            O => \N__13430\,
            I => \N__13426\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__13429\,
            I => \N__13423\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__13426\,
            I => \N__13418\
        );

    \I__2295\ : InMux
    port map (
            O => \N__13423\,
            I => \N__13411\
        );

    \I__2294\ : InMux
    port map (
            O => \N__13422\,
            I => \N__13411\
        );

    \I__2293\ : InMux
    port map (
            O => \N__13421\,
            I => \N__13411\
        );

    \I__2292\ : Span4Mux_v
    port map (
            O => \N__13418\,
            I => \N__13406\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__13411\,
            I => \N__13406\
        );

    \I__2290\ : Span4Mux_h
    port map (
            O => \N__13406\,
            I => \N__13403\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__13403\,
            I => \POWERLED.N_214\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__13400\,
            I => \N__13397\
        );

    \I__2287\ : InMux
    port map (
            O => \N__13397\,
            I => \N__13394\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__13394\,
            I => \N__13391\
        );

    \I__2285\ : Odrv4
    port map (
            O => \N__13391\,
            I => \POWERLED.dutycycle_RNI2V0PZ0Z_10\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__13388\,
            I => \POWERLED.dutycycle_RNI2V0PZ0Z_10_cascade_\
        );

    \I__2283\ : InMux
    port map (
            O => \N__13385\,
            I => \N__13382\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__13382\,
            I => \N__13379\
        );

    \I__2281\ : Odrv4
    port map (
            O => \N__13379\,
            I => \POWERLED.dutycycle_RNI712I1Z0Z_15\
        );

    \I__2280\ : InMux
    port map (
            O => \N__13376\,
            I => \N__13373\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__13373\,
            I => \N__13370\
        );

    \I__2278\ : Odrv4
    port map (
            O => \N__13370\,
            I => \POWERLED.dutycycle_RNIQ09G1Z0Z_10\
        );

    \I__2277\ : InMux
    port map (
            O => \N__13367\,
            I => \N__13363\
        );

    \I__2276\ : InMux
    port map (
            O => \N__13366\,
            I => \N__13360\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__13363\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__13360\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__2273\ : InMux
    port map (
            O => \N__13355\,
            I => \N__13351\
        );

    \I__2272\ : InMux
    port map (
            O => \N__13354\,
            I => \N__13348\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__13351\,
            I => \N__13345\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__13348\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__13345\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__13340\,
            I => \N__13336\
        );

    \I__2267\ : InMux
    port map (
            O => \N__13339\,
            I => \N__13333\
        );

    \I__2266\ : InMux
    port map (
            O => \N__13336\,
            I => \N__13330\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__13333\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__13330\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__2263\ : InMux
    port map (
            O => \N__13325\,
            I => \N__13321\
        );

    \I__2262\ : InMux
    port map (
            O => \N__13324\,
            I => \N__13318\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__13321\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__13318\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__2259\ : InMux
    port map (
            O => \N__13313\,
            I => \N__13310\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__13310\,
            I => \N__13307\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__13307\,
            I => \POWERLED.func_state_ns_0_a2_8_0\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__13304\,
            I => \POWERLED.un1_dutycycle_1_44_0_cascade_\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__13301\,
            I => \N__13298\
        );

    \I__2254\ : InMux
    port map (
            O => \N__13298\,
            I => \N__13295\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__13295\,
            I => \N__13292\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__13292\,
            I => \POWERLED.dutycycle_RNIF3561Z0Z_9\
        );

    \I__2251\ : InMux
    port map (
            O => \N__13289\,
            I => \N__13286\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__13286\,
            I => \POWERLED.dutycycle_RNIE4FLZ0Z_9\
        );

    \I__2249\ : InMux
    port map (
            O => \N__13283\,
            I => \N__13280\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__13280\,
            I => \POWERLED.dutycycle_RNI53MGZ0Z_14\
        );

    \I__2247\ : InMux
    port map (
            O => \N__13277\,
            I => \N__13274\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__13274\,
            I => \POWERLED.dutycycle_RNI84C11Z0Z_14\
        );

    \I__2245\ : InMux
    port map (
            O => \N__13271\,
            I => \N__13268\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__13268\,
            I => \POWERLED.dutycycle_RNIB1FLZ0Z_8\
        );

    \I__2243\ : CascadeMux
    port map (
            O => \N__13265\,
            I => \N__13262\
        );

    \I__2242\ : InMux
    port map (
            O => \N__13262\,
            I => \N__13259\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__13259\,
            I => \POWERLED.dutycycle_RNI75MGZ0Z_15\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__13256\,
            I => \POWERLED.un1_dutycycle_1_34_0_cascade_\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__13253\,
            I => \POWERLED.un1_dutycycle_1_axb_8_cascade_\
        );

    \I__2238\ : InMux
    port map (
            O => \N__13250\,
            I => \N__13247\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__13247\,
            I => \N__13243\
        );

    \I__2236\ : InMux
    port map (
            O => \N__13246\,
            I => \N__13240\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__13243\,
            I => \POWERLED.dutycycle_fast_RNILMLMZ0Z_6\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__13240\,
            I => \POWERLED.dutycycle_fast_RNILMLMZ0Z_6\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__13235\,
            I => \N__13232\
        );

    \I__2232\ : InMux
    port map (
            O => \N__13232\,
            I => \N__13229\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__13226\,
            I => \POWERLED.dutycycle_RNIJL1R1Z0Z_6\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__13223\,
            I => \N__13219\
        );

    \I__2228\ : InMux
    port map (
            O => \N__13222\,
            I => \N__13215\
        );

    \I__2227\ : InMux
    port map (
            O => \N__13219\,
            I => \N__13212\
        );

    \I__2226\ : InMux
    port map (
            O => \N__13218\,
            I => \N__13209\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__13215\,
            I => \POWERLED.dutycycle_fastZ0Z_6\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__13212\,
            I => \POWERLED.dutycycle_fastZ0Z_6\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__13209\,
            I => \POWERLED.dutycycle_fastZ0Z_6\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__13202\,
            I => \N__13199\
        );

    \I__2221\ : InMux
    port map (
            O => \N__13199\,
            I => \N__13195\
        );

    \I__2220\ : InMux
    port map (
            O => \N__13198\,
            I => \N__13192\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__13195\,
            I => \N__13189\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__13192\,
            I => \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__13189\,
            I => \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6\
        );

    \I__2216\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13180\
        );

    \I__2215\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13177\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__13180\,
            I => \N__13174\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__13177\,
            I => \N__13171\
        );

    \I__2212\ : Span4Mux_h
    port map (
            O => \N__13174\,
            I => \N__13168\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__13171\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__13168\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__2209\ : InMux
    port map (
            O => \N__13163\,
            I => \POWERLED.un1_dutycycle_1_cry_10\
        );

    \I__2208\ : InMux
    port map (
            O => \N__13160\,
            I => \N__13157\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__13157\,
            I => \N__13153\
        );

    \I__2206\ : InMux
    port map (
            O => \N__13156\,
            I => \N__13150\
        );

    \I__2205\ : Span4Mux_v
    port map (
            O => \N__13153\,
            I => \N__13147\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__13150\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__13147\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__2202\ : InMux
    port map (
            O => \N__13142\,
            I => \POWERLED.un1_dutycycle_1_cry_11\
        );

    \I__2201\ : InMux
    port map (
            O => \N__13139\,
            I => \N__13136\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__13136\,
            I => \N__13132\
        );

    \I__2199\ : InMux
    port map (
            O => \N__13135\,
            I => \N__13129\
        );

    \I__2198\ : Span4Mux_h
    port map (
            O => \N__13132\,
            I => \N__13126\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__13129\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__13126\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__2195\ : InMux
    port map (
            O => \N__13121\,
            I => \POWERLED.un1_dutycycle_1_cry_12\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__13118\,
            I => \N__13115\
        );

    \I__2193\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13111\
        );

    \I__2192\ : InMux
    port map (
            O => \N__13114\,
            I => \N__13108\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__13111\,
            I => \N__13105\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__13108\,
            I => \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__13105\,
            I => \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1\
        );

    \I__2188\ : InMux
    port map (
            O => \N__13100\,
            I => \POWERLED.un1_dutycycle_1_cry_13\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__13097\,
            I => \N__13092\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__13096\,
            I => \N__13089\
        );

    \I__2185\ : InMux
    port map (
            O => \N__13095\,
            I => \N__13079\
        );

    \I__2184\ : InMux
    port map (
            O => \N__13092\,
            I => \N__13079\
        );

    \I__2183\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13079\
        );

    \I__2182\ : InMux
    port map (
            O => \N__13088\,
            I => \N__13079\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__13079\,
            I => \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1\
        );

    \I__2180\ : InMux
    port map (
            O => \N__13076\,
            I => \POWERLED.un1_dutycycle_1_cry_14\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__13073\,
            I => \N__13070\
        );

    \I__2178\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13061\
        );

    \I__2177\ : InMux
    port map (
            O => \N__13069\,
            I => \N__13061\
        );

    \I__2176\ : InMux
    port map (
            O => \N__13068\,
            I => \N__13061\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__13061\,
            I => \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71\
        );

    \I__2174\ : InMux
    port map (
            O => \N__13058\,
            I => \bfn_6_7_0_\
        );

    \I__2173\ : InMux
    port map (
            O => \N__13055\,
            I => \POWERLED.CO2\
        );

    \I__2172\ : InMux
    port map (
            O => \N__13052\,
            I => \N__13046\
        );

    \I__2171\ : InMux
    port map (
            O => \N__13051\,
            I => \N__13046\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__13046\,
            I => \POWERLED.CO2_THRU_CO\
        );

    \I__2169\ : InMux
    port map (
            O => \N__13043\,
            I => \N__13038\
        );

    \I__2168\ : InMux
    port map (
            O => \N__13042\,
            I => \N__13035\
        );

    \I__2167\ : InMux
    port map (
            O => \N__13041\,
            I => \N__13032\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__13038\,
            I => \POWERLED.dutycycle_fastZ0Z_5\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__13035\,
            I => \POWERLED.dutycycle_fastZ0Z_5\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__13032\,
            I => \POWERLED.dutycycle_fastZ0Z_5\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__13025\,
            I => \N__13022\
        );

    \I__2162\ : InMux
    port map (
            O => \N__13022\,
            I => \N__13018\
        );

    \I__2161\ : InMux
    port map (
            O => \N__13021\,
            I => \N__13015\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__13018\,
            I => \N__13012\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__13015\,
            I => \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5\
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__13012\,
            I => \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5\
        );

    \I__2157\ : InMux
    port map (
            O => \N__13007\,
            I => \N__13003\
        );

    \I__2156\ : InMux
    port map (
            O => \N__13006\,
            I => \N__13000\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__13003\,
            I => \N__12997\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__13000\,
            I => \N__12992\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__12997\,
            I => \N__12992\
        );

    \I__2152\ : Span4Mux_v
    port map (
            O => \N__12992\,
            I => \N__12989\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__12989\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__2150\ : InMux
    port map (
            O => \N__12986\,
            I => \POWERLED.un1_dutycycle_1_cry_2\
        );

    \I__2149\ : InMux
    port map (
            O => \N__12983\,
            I => \N__12980\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__12980\,
            I => \N__12976\
        );

    \I__2147\ : InMux
    port map (
            O => \N__12979\,
            I => \N__12973\
        );

    \I__2146\ : Span4Mux_h
    port map (
            O => \N__12976\,
            I => \N__12968\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__12973\,
            I => \N__12968\
        );

    \I__2144\ : Span4Mux_v
    port map (
            O => \N__12968\,
            I => \N__12965\
        );

    \I__2143\ : Odrv4
    port map (
            O => \N__12965\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__2142\ : InMux
    port map (
            O => \N__12962\,
            I => \POWERLED.un1_dutycycle_1_cry_3\
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__12959\,
            I => \N__12956\
        );

    \I__2140\ : InMux
    port map (
            O => \N__12956\,
            I => \N__12953\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__12953\,
            I => \POWERLED.dutycycle_RNIEJ021Z0Z_4\
        );

    \I__2138\ : InMux
    port map (
            O => \N__12950\,
            I => \N__12946\
        );

    \I__2137\ : InMux
    port map (
            O => \N__12949\,
            I => \N__12943\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__12946\,
            I => \N__12940\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__12943\,
            I => \N__12935\
        );

    \I__2134\ : Span4Mux_s1_h
    port map (
            O => \N__12940\,
            I => \N__12935\
        );

    \I__2133\ : Span4Mux_h
    port map (
            O => \N__12935\,
            I => \N__12932\
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__12932\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__2131\ : InMux
    port map (
            O => \N__12929\,
            I => \POWERLED.un1_dutycycle_1_cry_4\
        );

    \I__2130\ : InMux
    port map (
            O => \N__12926\,
            I => \N__12923\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__12923\,
            I => \N__12920\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__12920\,
            I => \POWERLED.dutycycle_RNI6NI81Z0Z_5\
        );

    \I__2127\ : InMux
    port map (
            O => \N__12917\,
            I => \N__12913\
        );

    \I__2126\ : InMux
    port map (
            O => \N__12916\,
            I => \N__12910\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__12913\,
            I => \N__12907\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__12910\,
            I => \N__12904\
        );

    \I__2123\ : Span4Mux_v
    port map (
            O => \N__12907\,
            I => \N__12899\
        );

    \I__2122\ : Span4Mux_s1_h
    port map (
            O => \N__12904\,
            I => \N__12899\
        );

    \I__2121\ : Span4Mux_h
    port map (
            O => \N__12899\,
            I => \N__12896\
        );

    \I__2120\ : Odrv4
    port map (
            O => \N__12896\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__2119\ : InMux
    port map (
            O => \N__12893\,
            I => \POWERLED.un1_dutycycle_1_cry_5\
        );

    \I__2118\ : InMux
    port map (
            O => \N__12890\,
            I => \N__12887\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__12887\,
            I => \N__12884\
        );

    \I__2116\ : Span4Mux_h
    port map (
            O => \N__12884\,
            I => \N__12881\
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__12881\,
            I => \POWERLED.dutycycle_RNIJNBA1Z0Z_6\
        );

    \I__2114\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12875\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__12875\,
            I => \N__12871\
        );

    \I__2112\ : InMux
    port map (
            O => \N__12874\,
            I => \N__12868\
        );

    \I__2111\ : Span4Mux_v
    port map (
            O => \N__12871\,
            I => \N__12865\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__12868\,
            I => \N__12862\
        );

    \I__2109\ : Span4Mux_v
    port map (
            O => \N__12865\,
            I => \N__12857\
        );

    \I__2108\ : Span4Mux_s1_h
    port map (
            O => \N__12862\,
            I => \N__12857\
        );

    \I__2107\ : Span4Mux_h
    port map (
            O => \N__12857\,
            I => \N__12854\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__12854\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__2105\ : InMux
    port map (
            O => \N__12851\,
            I => \POWERLED.un1_dutycycle_1_cry_6\
        );

    \I__2104\ : InMux
    port map (
            O => \N__12848\,
            I => \N__12844\
        );

    \I__2103\ : InMux
    port map (
            O => \N__12847\,
            I => \N__12841\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__12844\,
            I => \N__12838\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__12841\,
            I => \N__12835\
        );

    \I__2100\ : Span4Mux_v
    port map (
            O => \N__12838\,
            I => \N__12832\
        );

    \I__2099\ : Span4Mux_h
    port map (
            O => \N__12835\,
            I => \N__12829\
        );

    \I__2098\ : Span4Mux_h
    port map (
            O => \N__12832\,
            I => \N__12826\
        );

    \I__2097\ : Odrv4
    port map (
            O => \N__12829\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__2096\ : Odrv4
    port map (
            O => \N__12826\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__2095\ : InMux
    port map (
            O => \N__12821\,
            I => \bfn_6_6_0_\
        );

    \I__2094\ : InMux
    port map (
            O => \N__12818\,
            I => \N__12815\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__12815\,
            I => \N__12812\
        );

    \I__2092\ : Span4Mux_v
    port map (
            O => \N__12812\,
            I => \N__12808\
        );

    \I__2091\ : InMux
    port map (
            O => \N__12811\,
            I => \N__12805\
        );

    \I__2090\ : Span4Mux_h
    port map (
            O => \N__12808\,
            I => \N__12802\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__12805\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__2088\ : Odrv4
    port map (
            O => \N__12802\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__2087\ : InMux
    port map (
            O => \N__12797\,
            I => \POWERLED.un1_dutycycle_1_cry_8\
        );

    \I__2086\ : InMux
    port map (
            O => \N__12794\,
            I => \N__12790\
        );

    \I__2085\ : InMux
    port map (
            O => \N__12793\,
            I => \N__12787\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__12790\,
            I => \N__12784\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__12787\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__2082\ : Odrv12
    port map (
            O => \N__12784\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__2081\ : InMux
    port map (
            O => \N__12779\,
            I => \POWERLED.un1_dutycycle_1_cry_9\
        );

    \I__2080\ : InMux
    port map (
            O => \N__12776\,
            I => \HDA_STRAP.un1_count_1_cry_11\
        );

    \I__2079\ : InMux
    port map (
            O => \N__12773\,
            I => \HDA_STRAP.un1_count_1_cry_12\
        );

    \I__2078\ : InMux
    port map (
            O => \N__12770\,
            I => \HDA_STRAP.un1_count_1_cry_13\
        );

    \I__2077\ : InMux
    port map (
            O => \N__12767\,
            I => \HDA_STRAP.un1_count_1_cry_14\
        );

    \I__2076\ : InMux
    port map (
            O => \N__12764\,
            I => \bfn_6_3_0_\
        );

    \I__2075\ : InMux
    port map (
            O => \N__12761\,
            I => \HDA_STRAP.un1_count_1_cry_16\
        );

    \I__2074\ : InMux
    port map (
            O => \N__12758\,
            I => \N__12754\
        );

    \I__2073\ : InMux
    port map (
            O => \N__12757\,
            I => \N__12751\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__12754\,
            I => \N__12746\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__12751\,
            I => \N__12746\
        );

    \I__2070\ : Span12Mux_s11_v
    port map (
            O => \N__12746\,
            I => \N__12743\
        );

    \I__2069\ : Odrv12
    port map (
            O => \N__12743\,
            I => \POWERLED.un1_dutycycle_1_axb_0\
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__12740\,
            I => \N__12737\
        );

    \I__2067\ : InMux
    port map (
            O => \N__12737\,
            I => \N__12734\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__12734\,
            I => \POWERLED.un1_dutycycle_1_axb_1\
        );

    \I__2065\ : InMux
    port map (
            O => \N__12731\,
            I => \N__12727\
        );

    \I__2064\ : InMux
    port map (
            O => \N__12730\,
            I => \N__12724\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__12727\,
            I => \N__12721\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__12724\,
            I => \N__12718\
        );

    \I__2061\ : Span4Mux_v
    port map (
            O => \N__12721\,
            I => \N__12715\
        );

    \I__2060\ : Span12Mux_s11_v
    port map (
            O => \N__12718\,
            I => \N__12712\
        );

    \I__2059\ : Odrv4
    port map (
            O => \N__12715\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__2058\ : Odrv12
    port map (
            O => \N__12712\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__2057\ : InMux
    port map (
            O => \N__12707\,
            I => \POWERLED.un1_dutycycle_1_cry_0\
        );

    \I__2056\ : InMux
    port map (
            O => \N__12704\,
            I => \N__12701\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__12701\,
            I => \POWERLED.dutycycle_RNI16B71Z0Z_5\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__12698\,
            I => \N__12694\
        );

    \I__2053\ : InMux
    port map (
            O => \N__12697\,
            I => \N__12691\
        );

    \I__2052\ : InMux
    port map (
            O => \N__12694\,
            I => \N__12688\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__12691\,
            I => \POWERLED.dutycycle_RNIFHLJZ0Z_0\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__12688\,
            I => \POWERLED.dutycycle_RNIFHLJZ0Z_0\
        );

    \I__2049\ : InMux
    port map (
            O => \N__12683\,
            I => \N__12679\
        );

    \I__2048\ : InMux
    port map (
            O => \N__12682\,
            I => \N__12676\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__12679\,
            I => \N__12671\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__12676\,
            I => \N__12671\
        );

    \I__2045\ : Span4Mux_v
    port map (
            O => \N__12671\,
            I => \N__12668\
        );

    \I__2044\ : Span4Mux_h
    port map (
            O => \N__12668\,
            I => \N__12665\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__12665\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__2042\ : InMux
    port map (
            O => \N__12662\,
            I => \POWERLED.un1_dutycycle_1_cry_1\
        );

    \I__2041\ : InMux
    port map (
            O => \N__12659\,
            I => \HDA_STRAP.un1_count_1_cry_2\
        );

    \I__2040\ : InMux
    port map (
            O => \N__12656\,
            I => \HDA_STRAP.un1_count_1_cry_3\
        );

    \I__2039\ : InMux
    port map (
            O => \N__12653\,
            I => \HDA_STRAP.un1_count_1_cry_4\
        );

    \I__2038\ : InMux
    port map (
            O => \N__12650\,
            I => \HDA_STRAP.un1_count_1_cry_5\
        );

    \I__2037\ : InMux
    port map (
            O => \N__12647\,
            I => \HDA_STRAP.un1_count_1_cry_6\
        );

    \I__2036\ : InMux
    port map (
            O => \N__12644\,
            I => \bfn_6_2_0_\
        );

    \I__2035\ : InMux
    port map (
            O => \N__12641\,
            I => \HDA_STRAP.un1_count_1_cry_8\
        );

    \I__2034\ : InMux
    port map (
            O => \N__12638\,
            I => \HDA_STRAP.un1_count_1_cry_9\
        );

    \I__2033\ : InMux
    port map (
            O => \N__12635\,
            I => \N__12632\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__12632\,
            I => \HDA_STRAP.count_RNO_0Z0Z_11\
        );

    \I__2031\ : InMux
    port map (
            O => \N__12629\,
            I => \HDA_STRAP.un1_count_1_cry_10\
        );

    \I__2030\ : InMux
    port map (
            O => \N__12626\,
            I => \N__12623\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__12623\,
            I => \N__12617\
        );

    \I__2028\ : InMux
    port map (
            O => \N__12622\,
            I => \N__12614\
        );

    \I__2027\ : InMux
    port map (
            O => \N__12621\,
            I => \N__12609\
        );

    \I__2026\ : InMux
    port map (
            O => \N__12620\,
            I => \N__12609\
        );

    \I__2025\ : Span4Mux_h
    port map (
            O => \N__12617\,
            I => \N__12606\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__12614\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__12609\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__2022\ : Odrv4
    port map (
            O => \N__12606\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__2021\ : InMux
    port map (
            O => \N__12599\,
            I => \POWERLED.un1_count_1_cry_12\
        );

    \I__2020\ : InMux
    port map (
            O => \N__12596\,
            I => \N__12593\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__12593\,
            I => \N__12587\
        );

    \I__2018\ : InMux
    port map (
            O => \N__12592\,
            I => \N__12584\
        );

    \I__2017\ : InMux
    port map (
            O => \N__12591\,
            I => \N__12581\
        );

    \I__2016\ : InMux
    port map (
            O => \N__12590\,
            I => \N__12578\
        );

    \I__2015\ : Span4Mux_h
    port map (
            O => \N__12587\,
            I => \N__12575\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__12584\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__12581\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__12578\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__12575\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__2010\ : InMux
    port map (
            O => \N__12566\,
            I => \POWERLED.un1_count_1_cry_13\
        );

    \I__2009\ : InMux
    port map (
            O => \N__12563\,
            I => \bfn_5_16_0_\
        );

    \I__2008\ : InMux
    port map (
            O => \N__12560\,
            I => \N__12557\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__12557\,
            I => \N__12553\
        );

    \I__2006\ : InMux
    port map (
            O => \N__12556\,
            I => \N__12548\
        );

    \I__2005\ : Span4Mux_h
    port map (
            O => \N__12553\,
            I => \N__12545\
        );

    \I__2004\ : InMux
    port map (
            O => \N__12552\,
            I => \N__12540\
        );

    \I__2003\ : InMux
    port map (
            O => \N__12551\,
            I => \N__12540\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__12548\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__2001\ : Odrv4
    port map (
            O => \N__12545\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__12540\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__1999\ : CEMux
    port map (
            O => \N__12533\,
            I => \N__12530\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__12530\,
            I => \N__12527\
        );

    \I__1997\ : Odrv12
    port map (
            O => \N__12527\,
            I => \POWERLED.N_65_5\
        );

    \I__1996\ : SRMux
    port map (
            O => \N__12524\,
            I => \N__12521\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__12521\,
            I => \N__12516\
        );

    \I__1994\ : SRMux
    port map (
            O => \N__12520\,
            I => \N__12511\
        );

    \I__1993\ : SRMux
    port map (
            O => \N__12519\,
            I => \N__12508\
        );

    \I__1992\ : Span4Mux_h
    port map (
            O => \N__12516\,
            I => \N__12505\
        );

    \I__1991\ : SRMux
    port map (
            O => \N__12515\,
            I => \N__12502\
        );

    \I__1990\ : InMux
    port map (
            O => \N__12514\,
            I => \N__12499\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__12511\,
            I => \POWERLED.curr_state_RNI75RB5Z0Z_0\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__12508\,
            I => \POWERLED.curr_state_RNI75RB5Z0Z_0\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__12505\,
            I => \POWERLED.curr_state_RNI75RB5Z0Z_0\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__12502\,
            I => \POWERLED.curr_state_RNI75RB5Z0Z_0\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__12499\,
            I => \POWERLED.curr_state_RNI75RB5Z0Z_0\
        );

    \I__1984\ : InMux
    port map (
            O => \N__12488\,
            I => \N__12485\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__12485\,
            I => \HDA_STRAP.count_RNO_0Z0Z_0\
        );

    \I__1982\ : InMux
    port map (
            O => \N__12482\,
            I => \HDA_STRAP.un1_count_1_cry_0\
        );

    \I__1981\ : InMux
    port map (
            O => \N__12479\,
            I => \HDA_STRAP.un1_count_1_cry_1\
        );

    \I__1980\ : InMux
    port map (
            O => \N__12476\,
            I => \N__12473\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__12473\,
            I => \N__12469\
        );

    \I__1978\ : InMux
    port map (
            O => \N__12472\,
            I => \N__12464\
        );

    \I__1977\ : Span4Mux_h
    port map (
            O => \N__12469\,
            I => \N__12461\
        );

    \I__1976\ : InMux
    port map (
            O => \N__12468\,
            I => \N__12456\
        );

    \I__1975\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12456\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__12464\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__12461\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__12456\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__1971\ : InMux
    port map (
            O => \N__12449\,
            I => \POWERLED.un1_count_1_cry_3\
        );

    \I__1970\ : InMux
    port map (
            O => \N__12446\,
            I => \N__12443\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__12443\,
            I => \N__12437\
        );

    \I__1968\ : InMux
    port map (
            O => \N__12442\,
            I => \N__12434\
        );

    \I__1967\ : InMux
    port map (
            O => \N__12441\,
            I => \N__12429\
        );

    \I__1966\ : InMux
    port map (
            O => \N__12440\,
            I => \N__12429\
        );

    \I__1965\ : Span4Mux_v
    port map (
            O => \N__12437\,
            I => \N__12426\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__12434\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__12429\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__12426\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1961\ : InMux
    port map (
            O => \N__12419\,
            I => \POWERLED.un1_count_1_cry_4\
        );

    \I__1960\ : InMux
    port map (
            O => \N__12416\,
            I => \N__12413\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__12413\,
            I => \N__12407\
        );

    \I__1958\ : InMux
    port map (
            O => \N__12412\,
            I => \N__12404\
        );

    \I__1957\ : InMux
    port map (
            O => \N__12411\,
            I => \N__12399\
        );

    \I__1956\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12399\
        );

    \I__1955\ : Span4Mux_h
    port map (
            O => \N__12407\,
            I => \N__12396\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__12404\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__12399\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__12396\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__1951\ : InMux
    port map (
            O => \N__12389\,
            I => \POWERLED.un1_count_1_cry_5\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__12386\,
            I => \N__12381\
        );

    \I__1949\ : InMux
    port map (
            O => \N__12385\,
            I => \N__12378\
        );

    \I__1948\ : InMux
    port map (
            O => \N__12384\,
            I => \N__12372\
        );

    \I__1947\ : InMux
    port map (
            O => \N__12381\,
            I => \N__12372\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__12378\,
            I => \N__12369\
        );

    \I__1945\ : InMux
    port map (
            O => \N__12377\,
            I => \N__12366\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__12372\,
            I => \N__12361\
        );

    \I__1943\ : Span4Mux_v
    port map (
            O => \N__12369\,
            I => \N__12361\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__12366\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__12361\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__1940\ : InMux
    port map (
            O => \N__12356\,
            I => \POWERLED.un1_count_1_cry_6\
        );

    \I__1939\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12349\
        );

    \I__1938\ : InMux
    port map (
            O => \N__12352\,
            I => \N__12344\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__12349\,
            I => \N__12341\
        );

    \I__1936\ : InMux
    port map (
            O => \N__12348\,
            I => \N__12336\
        );

    \I__1935\ : InMux
    port map (
            O => \N__12347\,
            I => \N__12336\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__12344\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__1933\ : Odrv4
    port map (
            O => \N__12341\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__12336\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__1931\ : InMux
    port map (
            O => \N__12329\,
            I => \POWERLED.un1_count_1_cry_7\
        );

    \I__1930\ : InMux
    port map (
            O => \N__12326\,
            I => \N__12322\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__12325\,
            I => \N__12317\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__12322\,
            I => \N__12314\
        );

    \I__1927\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12311\
        );

    \I__1926\ : InMux
    port map (
            O => \N__12320\,
            I => \N__12308\
        );

    \I__1925\ : InMux
    port map (
            O => \N__12317\,
            I => \N__12305\
        );

    \I__1924\ : Span4Mux_v
    port map (
            O => \N__12314\,
            I => \N__12302\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__12311\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__12308\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__12305\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1920\ : Odrv4
    port map (
            O => \N__12302\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1919\ : InMux
    port map (
            O => \N__12293\,
            I => \bfn_5_15_0_\
        );

    \I__1918\ : InMux
    port map (
            O => \N__12290\,
            I => \N__12287\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__12287\,
            I => \N__12283\
        );

    \I__1916\ : InMux
    port map (
            O => \N__12286\,
            I => \N__12278\
        );

    \I__1915\ : Span4Mux_v
    port map (
            O => \N__12283\,
            I => \N__12275\
        );

    \I__1914\ : InMux
    port map (
            O => \N__12282\,
            I => \N__12270\
        );

    \I__1913\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12270\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__12278\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__1911\ : Odrv4
    port map (
            O => \N__12275\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__12270\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__1909\ : InMux
    port map (
            O => \N__12263\,
            I => \POWERLED.un1_count_1_cry_9\
        );

    \I__1908\ : InMux
    port map (
            O => \N__12260\,
            I => \N__12257\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__12257\,
            I => \N__12251\
        );

    \I__1906\ : InMux
    port map (
            O => \N__12256\,
            I => \N__12248\
        );

    \I__1905\ : InMux
    port map (
            O => \N__12255\,
            I => \N__12245\
        );

    \I__1904\ : InMux
    port map (
            O => \N__12254\,
            I => \N__12242\
        );

    \I__1903\ : Span4Mux_h
    port map (
            O => \N__12251\,
            I => \N__12239\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__12248\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__12245\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__12242\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__1899\ : Odrv4
    port map (
            O => \N__12239\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__1898\ : InMux
    port map (
            O => \N__12230\,
            I => \POWERLED.un1_count_1_cry_10\
        );

    \I__1897\ : InMux
    port map (
            O => \N__12227\,
            I => \N__12224\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__12224\,
            I => \N__12218\
        );

    \I__1895\ : InMux
    port map (
            O => \N__12223\,
            I => \N__12215\
        );

    \I__1894\ : InMux
    port map (
            O => \N__12222\,
            I => \N__12212\
        );

    \I__1893\ : InMux
    port map (
            O => \N__12221\,
            I => \N__12209\
        );

    \I__1892\ : Span4Mux_h
    port map (
            O => \N__12218\,
            I => \N__12206\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__12215\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__12212\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__12209\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__12206\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__1887\ : InMux
    port map (
            O => \N__12197\,
            I => \POWERLED.un1_count_1_cry_11\
        );

    \I__1886\ : InMux
    port map (
            O => \N__12194\,
            I => \N__12190\
        );

    \I__1885\ : InMux
    port map (
            O => \N__12193\,
            I => \N__12187\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__12190\,
            I => \N__12184\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__12187\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__12184\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__1881\ : InMux
    port map (
            O => \N__12179\,
            I => \N__12175\
        );

    \I__1880\ : InMux
    port map (
            O => \N__12178\,
            I => \N__12172\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__12175\,
            I => \N__12169\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__12172\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__1877\ : Odrv4
    port map (
            O => \N__12169\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__12164\,
            I => \N__12160\
        );

    \I__1875\ : InMux
    port map (
            O => \N__12163\,
            I => \N__12157\
        );

    \I__1874\ : InMux
    port map (
            O => \N__12160\,
            I => \N__12154\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__12157\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__12154\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__1871\ : InMux
    port map (
            O => \N__12149\,
            I => \N__12145\
        );

    \I__1870\ : InMux
    port map (
            O => \N__12148\,
            I => \N__12142\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__12145\,
            I => \N__12139\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__12142\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__1867\ : Odrv4
    port map (
            O => \N__12139\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__1866\ : InMux
    port map (
            O => \N__12134\,
            I => \N__12131\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__12131\,
            I => \POWERLED.func_state_ns_0_a2_11_0\
        );

    \I__1864\ : InMux
    port map (
            O => \N__12128\,
            I => \N__12125\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__12125\,
            I => \POWERLED.func_state_ns_0_a2_10_0\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__12122\,
            I => \POWERLED.func_state_ns_0_a2_9_0_cascade_\
        );

    \I__1861\ : InMux
    port map (
            O => \N__12119\,
            I => \N__12105\
        );

    \I__1860\ : InMux
    port map (
            O => \N__12118\,
            I => \N__12098\
        );

    \I__1859\ : InMux
    port map (
            O => \N__12117\,
            I => \N__12098\
        );

    \I__1858\ : InMux
    port map (
            O => \N__12116\,
            I => \N__12098\
        );

    \I__1857\ : InMux
    port map (
            O => \N__12115\,
            I => \N__12089\
        );

    \I__1856\ : InMux
    port map (
            O => \N__12114\,
            I => \N__12089\
        );

    \I__1855\ : InMux
    port map (
            O => \N__12113\,
            I => \N__12089\
        );

    \I__1854\ : InMux
    port map (
            O => \N__12112\,
            I => \N__12089\
        );

    \I__1853\ : InMux
    port map (
            O => \N__12111\,
            I => \N__12080\
        );

    \I__1852\ : InMux
    port map (
            O => \N__12110\,
            I => \N__12080\
        );

    \I__1851\ : InMux
    port map (
            O => \N__12109\,
            I => \N__12080\
        );

    \I__1850\ : InMux
    port map (
            O => \N__12108\,
            I => \N__12080\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__12105\,
            I => \N__12075\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__12098\,
            I => \N__12075\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__12089\,
            I => \POWERLED.count_off_0_sqmuxa\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__12080\,
            I => \POWERLED.count_off_0_sqmuxa\
        );

    \I__1845\ : Odrv12
    port map (
            O => \N__12075\,
            I => \POWERLED.count_off_0_sqmuxa\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__12068\,
            I => \POWERLED.count_off_0_sqmuxa_cascade_\
        );

    \I__1843\ : InMux
    port map (
            O => \N__12065\,
            I => \N__12059\
        );

    \I__1842\ : InMux
    port map (
            O => \N__12064\,
            I => \N__12052\
        );

    \I__1841\ : InMux
    port map (
            O => \N__12063\,
            I => \N__12052\
        );

    \I__1840\ : InMux
    port map (
            O => \N__12062\,
            I => \N__12052\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__12059\,
            I => \N__12049\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__12052\,
            I => \N__12046\
        );

    \I__1837\ : Odrv4
    port map (
            O => \N__12049\,
            I => \POWERLED.N_85_1\
        );

    \I__1836\ : Odrv12
    port map (
            O => \N__12046\,
            I => \POWERLED.N_85_1\
        );

    \I__1835\ : InMux
    port map (
            O => \N__12041\,
            I => \N__12035\
        );

    \I__1834\ : InMux
    port map (
            O => \N__12040\,
            I => \N__12030\
        );

    \I__1833\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12030\
        );

    \I__1832\ : InMux
    port map (
            O => \N__12038\,
            I => \N__12027\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__12035\,
            I => \N__12024\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__12030\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__12027\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__1828\ : Odrv4
    port map (
            O => \N__12024\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__1827\ : InMux
    port map (
            O => \N__12017\,
            I => \N__12012\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__12016\,
            I => \N__12009\
        );

    \I__1825\ : InMux
    port map (
            O => \N__12015\,
            I => \N__12006\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__12012\,
            I => \N__12003\
        );

    \I__1823\ : InMux
    port map (
            O => \N__12009\,
            I => \N__12000\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__12006\,
            I => \N__11995\
        );

    \I__1821\ : Span4Mux_s2_h
    port map (
            O => \N__12003\,
            I => \N__11995\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__12000\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__1819\ : Odrv4
    port map (
            O => \N__11995\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__1818\ : InMux
    port map (
            O => \N__11990\,
            I => \N__11987\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__11987\,
            I => \N__11983\
        );

    \I__1816\ : InMux
    port map (
            O => \N__11986\,
            I => \N__11978\
        );

    \I__1815\ : Span4Mux_v
    port map (
            O => \N__11983\,
            I => \N__11975\
        );

    \I__1814\ : InMux
    port map (
            O => \N__11982\,
            I => \N__11970\
        );

    \I__1813\ : InMux
    port map (
            O => \N__11981\,
            I => \N__11970\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__11978\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__11975\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__11970\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__1809\ : InMux
    port map (
            O => \N__11963\,
            I => \POWERLED.un1_count_1_cry_1\
        );

    \I__1808\ : InMux
    port map (
            O => \N__11960\,
            I => \N__11957\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__11957\,
            I => \N__11953\
        );

    \I__1806\ : InMux
    port map (
            O => \N__11956\,
            I => \N__11948\
        );

    \I__1805\ : Span4Mux_h
    port map (
            O => \N__11953\,
            I => \N__11945\
        );

    \I__1804\ : InMux
    port map (
            O => \N__11952\,
            I => \N__11940\
        );

    \I__1803\ : InMux
    port map (
            O => \N__11951\,
            I => \N__11940\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__11948\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__11945\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__11940\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__1799\ : InMux
    port map (
            O => \N__11933\,
            I => \POWERLED.un1_count_1_cry_2\
        );

    \I__1798\ : InMux
    port map (
            O => \N__11930\,
            I => \POWERLED.un1_count_off_1_cry_8\
        );

    \I__1797\ : InMux
    port map (
            O => \N__11927\,
            I => \POWERLED.un1_count_off_1_cry_9\
        );

    \I__1796\ : InMux
    port map (
            O => \N__11924\,
            I => \POWERLED.un1_count_off_1_cry_10\
        );

    \I__1795\ : InMux
    port map (
            O => \N__11921\,
            I => \POWERLED.un1_count_off_1_cry_11\
        );

    \I__1794\ : InMux
    port map (
            O => \N__11918\,
            I => \POWERLED.un1_count_off_1_cry_12\
        );

    \I__1793\ : InMux
    port map (
            O => \N__11915\,
            I => \POWERLED.un1_count_off_1_cry_13\
        );

    \I__1792\ : InMux
    port map (
            O => \N__11912\,
            I => \POWERLED.un1_count_off_1_cry_14\
        );

    \I__1791\ : InMux
    port map (
            O => \N__11909\,
            I => \N__11905\
        );

    \I__1790\ : InMux
    port map (
            O => \N__11908\,
            I => \N__11902\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__11905\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__11902\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__1787\ : InMux
    port map (
            O => \N__11897\,
            I => \N__11893\
        );

    \I__1786\ : InMux
    port map (
            O => \N__11896\,
            I => \N__11890\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__11893\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__11890\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__11885\,
            I => \N__11881\
        );

    \I__1782\ : InMux
    port map (
            O => \N__11884\,
            I => \N__11878\
        );

    \I__1781\ : InMux
    port map (
            O => \N__11881\,
            I => \N__11875\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__11878\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__11875\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__1778\ : InMux
    port map (
            O => \N__11870\,
            I => \N__11866\
        );

    \I__1777\ : InMux
    port map (
            O => \N__11869\,
            I => \N__11863\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__11866\,
            I => \N__11860\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__11863\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__11860\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__1773\ : InMux
    port map (
            O => \N__11855\,
            I => \N__11851\
        );

    \I__1772\ : InMux
    port map (
            O => \N__11854\,
            I => \N__11848\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__11851\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__11848\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__1769\ : InMux
    port map (
            O => \N__11843\,
            I => \N__11839\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11842\,
            I => \N__11836\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__11839\,
            I => \N__11833\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__11836\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__11833\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__11828\,
            I => \N__11824\
        );

    \I__1763\ : InMux
    port map (
            O => \N__11827\,
            I => \N__11821\
        );

    \I__1762\ : InMux
    port map (
            O => \N__11824\,
            I => \N__11818\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__11821\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__11818\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__1759\ : InMux
    port map (
            O => \N__11813\,
            I => \N__11809\
        );

    \I__1758\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11806\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__11809\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__11806\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__1755\ : InMux
    port map (
            O => \N__11801\,
            I => \POWERLED.un1_count_off_1_cry_0\
        );

    \I__1754\ : InMux
    port map (
            O => \N__11798\,
            I => \POWERLED.un1_count_off_1_cry_1\
        );

    \I__1753\ : InMux
    port map (
            O => \N__11795\,
            I => \POWERLED.un1_count_off_1_cry_2\
        );

    \I__1752\ : InMux
    port map (
            O => \N__11792\,
            I => \POWERLED.un1_count_off_1_cry_3\
        );

    \I__1751\ : InMux
    port map (
            O => \N__11789\,
            I => \POWERLED.un1_count_off_1_cry_4\
        );

    \I__1750\ : InMux
    port map (
            O => \N__11786\,
            I => \POWERLED.un1_count_off_1_cry_5\
        );

    \I__1749\ : InMux
    port map (
            O => \N__11783\,
            I => \POWERLED.un1_count_off_1_cry_6\
        );

    \I__1748\ : InMux
    port map (
            O => \N__11780\,
            I => \bfn_5_10_0_\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__11777\,
            I => \N__11774\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11774\,
            I => \N__11771\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__11771\,
            I => \POWERLED.un1_dutycycle_1_i_29\
        );

    \I__1744\ : InMux
    port map (
            O => \N__11768\,
            I => \N__11765\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__11765\,
            I => \N__11762\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__11762\,
            I => \POWERLED.mult1_un61_sum_i\
        );

    \I__1741\ : InMux
    port map (
            O => \N__11759\,
            I => \N__11756\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__11756\,
            I => \POWERLED.mult1_un54_sum_i\
        );

    \I__1739\ : InMux
    port map (
            O => \N__11753\,
            I => \N__11750\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__11750\,
            I => \N__11747\
        );

    \I__1737\ : Odrv12
    port map (
            O => \N__11747\,
            I => \POWERLED.mult1_un75_sum_i\
        );

    \I__1736\ : InMux
    port map (
            O => \N__11744\,
            I => \N__11738\
        );

    \I__1735\ : InMux
    port map (
            O => \N__11743\,
            I => \N__11738\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__11738\,
            I => \N__11735\
        );

    \I__1733\ : Span4Mux_h
    port map (
            O => \N__11735\,
            I => \N__11732\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__11732\,
            I => \POWERLED.N_53\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__11729\,
            I => \N__11726\
        );

    \I__1730\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11723\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__11723\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_4\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__11720\,
            I => \N__11717\
        );

    \I__1727\ : InMux
    port map (
            O => \N__11717\,
            I => \N__11714\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__11714\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_5\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__11711\,
            I => \N__11708\
        );

    \I__1724\ : InMux
    port map (
            O => \N__11708\,
            I => \N__11705\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__11705\,
            I => \POWERLED.mult1_un47_sum_axb_4\
        );

    \I__1722\ : InMux
    port map (
            O => \N__11702\,
            I => \N__11698\
        );

    \I__1721\ : InMux
    port map (
            O => \N__11701\,
            I => \N__11695\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__11698\,
            I => \HDA_STRAP.N_5_0\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__11695\,
            I => \HDA_STRAP.N_5_0\
        );

    \I__1718\ : InMux
    port map (
            O => \N__11690\,
            I => \N__11684\
        );

    \I__1717\ : InMux
    port map (
            O => \N__11689\,
            I => \N__11684\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__11684\,
            I => \HDA_STRAP.curr_stateZ0Z_2\
        );

    \I__1715\ : IoInMux
    port map (
            O => \N__11681\,
            I => \N__11678\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__11678\,
            I => \N__11675\
        );

    \I__1713\ : IoSpan4Mux
    port map (
            O => \N__11675\,
            I => \N__11672\
        );

    \I__1712\ : Span4Mux_s0_h
    port map (
            O => \N__11672\,
            I => \N__11669\
        );

    \I__1711\ : Span4Mux_h
    port map (
            O => \N__11669\,
            I => \N__11666\
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__11666\,
            I => hda_sdo_atp
        );

    \I__1709\ : InMux
    port map (
            O => \N__11663\,
            I => \N__11660\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__11660\,
            I => \N__11657\
        );

    \I__1707\ : Odrv12
    port map (
            O => \N__11657\,
            I => \POWERLED.mult1_un82_sum_i\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__11654\,
            I => \N__11651\
        );

    \I__1705\ : InMux
    port map (
            O => \N__11651\,
            I => \N__11648\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__11648\,
            I => \POWERLED.un1_dutycycle_1_i_28\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__11645\,
            I => \POWERLED.un1_dutycycle_1_19_0_cascade_\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__11642\,
            I => \POWERLED.un1_countlto15_5_cascade_\
        );

    \I__1701\ : InMux
    port map (
            O => \N__11639\,
            I => \N__11636\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__11636\,
            I => \POWERLED.g0_0_4\
        );

    \I__1699\ : InMux
    port map (
            O => \N__11633\,
            I => \N__11630\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__11630\,
            I => \POWERLED.un1_countlt6\
        );

    \I__1697\ : InMux
    port map (
            O => \N__11627\,
            I => \N__11624\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__11624\,
            I => \POWERLED.g0_0_5\
        );

    \I__1695\ : CascadeMux
    port map (
            O => \N__11621\,
            I => \POWERLED.un1_countlto15_4_cascade_\
        );

    \I__1694\ : InMux
    port map (
            O => \N__11618\,
            I => \N__11615\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__11615\,
            I => \POWERLED.un1_countlto15_7\
        );

    \I__1692\ : InMux
    port map (
            O => \N__11612\,
            I => \N__11609\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__11609\,
            I => \N__11606\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__11606\,
            I => \POWERLED.count_RNIOVT24Z0Z_11\
        );

    \I__1689\ : InMux
    port map (
            O => \N__11603\,
            I => \N__11597\
        );

    \I__1688\ : InMux
    port map (
            O => \N__11602\,
            I => \N__11594\
        );

    \I__1687\ : InMux
    port map (
            O => \N__11601\,
            I => \N__11591\
        );

    \I__1686\ : InMux
    port map (
            O => \N__11600\,
            I => \N__11588\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__11597\,
            I => \N__11585\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__11594\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__11591\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__11588\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__1681\ : Odrv12
    port map (
            O => \N__11585\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__11576\,
            I => \POWERLED.count_RNIOVT24Z0Z_11_cascade_\
        );

    \I__1679\ : IoInMux
    port map (
            O => \N__11573\,
            I => \N__11570\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__11570\,
            I => \N__11566\
        );

    \I__1677\ : IoInMux
    port map (
            O => \N__11569\,
            I => \N__11563\
        );

    \I__1676\ : Span4Mux_s3_h
    port map (
            O => \N__11566\,
            I => \N__11560\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__11563\,
            I => \N__11557\
        );

    \I__1674\ : Odrv4
    port map (
            O => \N__11560\,
            I => v5s_enn
        );

    \I__1673\ : Odrv12
    port map (
            O => \N__11557\,
            I => v5s_enn
        );

    \I__1672\ : InMux
    port map (
            O => \N__11552\,
            I => \N__11549\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__11549\,
            I => \N__11546\
        );

    \I__1670\ : Span4Mux_v
    port map (
            O => \N__11546\,
            I => \N__11543\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__11543\,
            I => \POWERLED.mult1_un159_sum_i\
        );

    \I__1668\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11537\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__11537\,
            I => \N__11534\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__11534\,
            I => \POWERLED.mult1_un152_sum_i\
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__11531\,
            I => \POWERLED.un1_countlt6_0_cascade_\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__11528\,
            I => \POWERLED.g0_0_7_cascade_\
        );

    \I__1663\ : InMux
    port map (
            O => \N__11525\,
            I => \N__11522\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__11522\,
            I => \N__11519\
        );

    \I__1661\ : Span4Mux_s3_h
    port map (
            O => \N__11519\,
            I => \N__11516\
        );

    \I__1660\ : Odrv4
    port map (
            O => \N__11516\,
            I => \POWERLED.un1_count_0\
        );

    \I__1659\ : InMux
    port map (
            O => \N__11513\,
            I => \N__11509\
        );

    \I__1658\ : InMux
    port map (
            O => \N__11512\,
            I => \N__11506\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__11509\,
            I => \POWERLED.mult1_un47_sum_cry_6_s\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__11506\,
            I => \POWERLED.mult1_un47_sum_cry_6_s\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__11501\,
            I => \N__11496\
        );

    \I__1654\ : InMux
    port map (
            O => \N__11500\,
            I => \N__11488\
        );

    \I__1653\ : InMux
    port map (
            O => \N__11499\,
            I => \N__11488\
        );

    \I__1652\ : InMux
    port map (
            O => \N__11496\,
            I => \N__11488\
        );

    \I__1651\ : InMux
    port map (
            O => \N__11495\,
            I => \N__11485\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__11488\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__11485\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__11480\,
            I => \N__11477\
        );

    \I__1647\ : InMux
    port map (
            O => \N__11477\,
            I => \N__11474\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__11474\,
            I => \N__11471\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__11471\,
            I => \POWERLED.mult1_un54_sum_cry_6_THRU_CO\
        );

    \I__1644\ : InMux
    port map (
            O => \N__11468\,
            I => \POWERLED.mult1_un61_sum_cry_7\
        );

    \I__1643\ : InMux
    port map (
            O => \N__11465\,
            I => \N__11461\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__11464\,
            I => \N__11457\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__11461\,
            I => \N__11454\
        );

    \I__1640\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11449\
        );

    \I__1639\ : InMux
    port map (
            O => \N__11457\,
            I => \N__11449\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__11454\,
            I => \N__11442\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__11449\,
            I => \N__11442\
        );

    \I__1636\ : InMux
    port map (
            O => \N__11448\,
            I => \N__11439\
        );

    \I__1635\ : InMux
    port map (
            O => \N__11447\,
            I => \N__11436\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__11442\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__11439\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__11436\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__11429\,
            I => \N__11425\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__11428\,
            I => \N__11421\
        );

    \I__1629\ : InMux
    port map (
            O => \N__11425\,
            I => \N__11414\
        );

    \I__1628\ : InMux
    port map (
            O => \N__11424\,
            I => \N__11414\
        );

    \I__1627\ : InMux
    port map (
            O => \N__11421\,
            I => \N__11414\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__11414\,
            I => \N__11411\
        );

    \I__1625\ : Odrv4
    port map (
            O => \N__11411\,
            I => \POWERLED.mult1_un61_sum_i_0_8\
        );

    \I__1624\ : InMux
    port map (
            O => \N__11408\,
            I => \N__11405\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__11405\,
            I => \N__11402\
        );

    \I__1622\ : Span4Mux_h
    port map (
            O => \N__11402\,
            I => \N__11399\
        );

    \I__1621\ : Odrv4
    port map (
            O => \N__11399\,
            I => \POWERLED.mult1_un110_sum_i\
        );

    \I__1620\ : InMux
    port map (
            O => \N__11396\,
            I => \N__11393\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__11393\,
            I => \N__11390\
        );

    \I__1618\ : Span4Mux_s3_h
    port map (
            O => \N__11390\,
            I => \N__11387\
        );

    \I__1617\ : Sp12to4
    port map (
            O => \N__11387\,
            I => \N__11384\
        );

    \I__1616\ : Odrv12
    port map (
            O => \N__11384\,
            I => \POWERLED.mult1_un138_sum_i\
        );

    \I__1615\ : InMux
    port map (
            O => \N__11381\,
            I => \N__11378\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__11378\,
            I => \N__11375\
        );

    \I__1613\ : Span4Mux_h
    port map (
            O => \N__11375\,
            I => \N__11372\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__11372\,
            I => \POWERLED.mult1_un124_sum_i\
        );

    \I__1611\ : InMux
    port map (
            O => \N__11369\,
            I => \N__11366\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__11366\,
            I => \N__11363\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__11363\,
            I => \POWERLED.mult1_un117_sum_i\
        );

    \I__1608\ : InMux
    port map (
            O => \N__11360\,
            I => \N__11357\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__11357\,
            I => \N__11353\
        );

    \I__1606\ : InMux
    port map (
            O => \N__11356\,
            I => \N__11350\
        );

    \I__1605\ : Odrv4
    port map (
            O => \N__11353\,
            I => \POWERLED.mult1_un138_sum_cry_6_s\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__11350\,
            I => \POWERLED.mult1_un138_sum_cry_6_s\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__11345\,
            I => \N__11342\
        );

    \I__1602\ : InMux
    port map (
            O => \N__11342\,
            I => \N__11339\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__11339\,
            I => \N__11336\
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__11336\,
            I => \POWERLED.mult1_un145_sum_axb_7_l_fx\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__11333\,
            I => \N__11327\
        );

    \I__1598\ : InMux
    port map (
            O => \N__11332\,
            I => \N__11320\
        );

    \I__1597\ : InMux
    port map (
            O => \N__11331\,
            I => \N__11320\
        );

    \I__1596\ : InMux
    port map (
            O => \N__11330\,
            I => \N__11315\
        );

    \I__1595\ : InMux
    port map (
            O => \N__11327\,
            I => \N__11315\
        );

    \I__1594\ : InMux
    port map (
            O => \N__11326\,
            I => \N__11312\
        );

    \I__1593\ : InMux
    port map (
            O => \N__11325\,
            I => \N__11309\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__11320\,
            I => \N__11306\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__11315\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__11312\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__11309\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__1588\ : Odrv12
    port map (
            O => \N__11306\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__1587\ : InMux
    port map (
            O => \N__11297\,
            I => \N__11294\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__11294\,
            I => \N__11291\
        );

    \I__1585\ : Span4Mux_s3_h
    port map (
            O => \N__11291\,
            I => \N__11288\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__11288\,
            I => \POWERLED.un1_count_2_4\
        );

    \I__1583\ : InMux
    port map (
            O => \N__11285\,
            I => \N__11282\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__11282\,
            I => \N__11279\
        );

    \I__1581\ : Odrv12
    port map (
            O => \N__11279\,
            I => \POWERLED.mult1_un68_sum_i\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__11276\,
            I => \N__11273\
        );

    \I__1579\ : InMux
    port map (
            O => \N__11273\,
            I => \N__11270\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__11270\,
            I => \N__11267\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__11267\,
            I => \POWERLED.mult1_un61_sum_cry_3_s\
        );

    \I__1576\ : InMux
    port map (
            O => \N__11264\,
            I => \POWERLED.mult1_un61_sum_cry_2\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__11261\,
            I => \N__11258\
        );

    \I__1574\ : InMux
    port map (
            O => \N__11258\,
            I => \N__11255\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__11255\,
            I => \N__11252\
        );

    \I__1572\ : Span4Mux_h
    port map (
            O => \N__11252\,
            I => \N__11249\
        );

    \I__1571\ : Odrv4
    port map (
            O => \N__11249\,
            I => \POWERLED.mult1_un54_sum_cry_3_s\
        );

    \I__1570\ : InMux
    port map (
            O => \N__11246\,
            I => \N__11243\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__11243\,
            I => \N__11240\
        );

    \I__1568\ : Odrv4
    port map (
            O => \N__11240\,
            I => \POWERLED.mult1_un61_sum_cry_4_s\
        );

    \I__1567\ : InMux
    port map (
            O => \N__11237\,
            I => \POWERLED.mult1_un61_sum_cry_3\
        );

    \I__1566\ : InMux
    port map (
            O => \N__11234\,
            I => \N__11231\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__11231\,
            I => \N__11228\
        );

    \I__1564\ : Odrv12
    port map (
            O => \N__11228\,
            I => \POWERLED.mult1_un54_sum_cry_4_s\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__11225\,
            I => \N__11222\
        );

    \I__1562\ : InMux
    port map (
            O => \N__11222\,
            I => \N__11219\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__11219\,
            I => \N__11216\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__11216\,
            I => \POWERLED.mult1_un61_sum_cry_5_s\
        );

    \I__1559\ : InMux
    port map (
            O => \N__11213\,
            I => \POWERLED.mult1_un61_sum_cry_4\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__11210\,
            I => \N__11207\
        );

    \I__1557\ : InMux
    port map (
            O => \N__11207\,
            I => \N__11204\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__11204\,
            I => \N__11201\
        );

    \I__1555\ : Odrv4
    port map (
            O => \N__11201\,
            I => \POWERLED.mult1_un54_sum_cry_5_s\
        );

    \I__1554\ : InMux
    port map (
            O => \N__11198\,
            I => \N__11195\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__11195\,
            I => \N__11192\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__11192\,
            I => \POWERLED.mult1_un61_sum_cry_6_s\
        );

    \I__1551\ : InMux
    port map (
            O => \N__11189\,
            I => \POWERLED.mult1_un61_sum_cry_5\
        );

    \I__1550\ : InMux
    port map (
            O => \N__11186\,
            I => \N__11183\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__11183\,
            I => \N__11180\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__11180\,
            I => \POWERLED.mult1_un54_sum_cry_6_s\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__11177\,
            I => \N__11173\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__11176\,
            I => \N__11169\
        );

    \I__1545\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11162\
        );

    \I__1544\ : InMux
    port map (
            O => \N__11172\,
            I => \N__11162\
        );

    \I__1543\ : InMux
    port map (
            O => \N__11169\,
            I => \N__11162\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__11162\,
            I => \POWERLED.mult1_un54_sum_i_8\
        );

    \I__1541\ : InMux
    port map (
            O => \N__11159\,
            I => \N__11156\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__11156\,
            I => \N__11153\
        );

    \I__1539\ : Odrv4
    port map (
            O => \N__11153\,
            I => \POWERLED.mult1_un68_sum_axb_8\
        );

    \I__1538\ : InMux
    port map (
            O => \N__11150\,
            I => \POWERLED.mult1_un61_sum_cry_6\
        );

    \I__1537\ : InMux
    port map (
            O => \N__11147\,
            I => \POWERLED.mult1_un54_sum_cry_5\
        );

    \I__1536\ : InMux
    port map (
            O => \N__11144\,
            I => \POWERLED.mult1_un54_sum_cry_6\
        );

    \I__1535\ : InMux
    port map (
            O => \N__11141\,
            I => \POWERLED.mult1_un54_sum_cry_7\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__11138\,
            I => \N__11135\
        );

    \I__1533\ : InMux
    port map (
            O => \N__11135\,
            I => \N__11132\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__11132\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__1531\ : InMux
    port map (
            O => \N__11129\,
            I => \POWERLED.mult1_un47_sum_cry_2\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__11126\,
            I => \N__11123\
        );

    \I__1529\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11120\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__11120\,
            I => \POWERLED.mult1_un47_sum_cry_4_s\
        );

    \I__1527\ : InMux
    port map (
            O => \N__11117\,
            I => \POWERLED.mult1_un47_sum_cry_3\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__11114\,
            I => \N__11111\
        );

    \I__1525\ : InMux
    port map (
            O => \N__11111\,
            I => \N__11108\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__11108\,
            I => \POWERLED.mult1_un47_sum_cry_5_s\
        );

    \I__1523\ : InMux
    port map (
            O => \N__11105\,
            I => \POWERLED.mult1_un47_sum_cry_4\
        );

    \I__1522\ : InMux
    port map (
            O => \N__11102\,
            I => \POWERLED.mult1_un47_sum_cry_5\
        );

    \I__1521\ : InMux
    port map (
            O => \N__11099\,
            I => \N__11096\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__11096\,
            I => \POWERLED.mult1_un54_sum_cry_7_THRU_CO\
        );

    \I__1519\ : InMux
    port map (
            O => \N__11093\,
            I => \POWERLED.mult1_un47_sum_cry_6\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__11090\,
            I => \POWERLED.un1_count_2_cry_15_THRU_CO_cascade_\
        );

    \I__1517\ : CEMux
    port map (
            O => \N__11087\,
            I => \N__11084\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__11084\,
            I => \N__11081\
        );

    \I__1515\ : Span4Mux_v
    port map (
            O => \N__11081\,
            I => \N__11078\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__11078\,
            I => \POWERLED.pwm_out_RNOZ0\
        );

    \I__1513\ : InMux
    port map (
            O => \N__11075\,
            I => \N__11072\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__11072\,
            I => \N__11069\
        );

    \I__1511\ : Span4Mux_s3_v
    port map (
            O => \N__11069\,
            I => \N__11066\
        );

    \I__1510\ : Odrv4
    port map (
            O => \N__11066\,
            I => vpp_ok
        );

    \I__1509\ : IoInMux
    port map (
            O => \N__11063\,
            I => \N__11060\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__11060\,
            I => \N__11057\
        );

    \I__1507\ : Span4Mux_s1_v
    port map (
            O => \N__11057\,
            I => \N__11054\
        );

    \I__1506\ : Odrv4
    port map (
            O => \N__11054\,
            I => vddq_en
        );

    \I__1505\ : InMux
    port map (
            O => \N__11051\,
            I => \N__11048\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__11048\,
            I => \N__11045\
        );

    \I__1503\ : Span4Mux_v
    port map (
            O => \N__11045\,
            I => \N__11042\
        );

    \I__1502\ : Span4Mux_h
    port map (
            O => \N__11042\,
            I => \N__11039\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__11039\,
            I => gpio_fpga_soc_1
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__11036\,
            I => \HDA_STRAP.N_5_0_cascade_\
        );

    \I__1499\ : IoInMux
    port map (
            O => \N__11033\,
            I => \N__11030\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__11030\,
            I => \N__11026\
        );

    \I__1497\ : InMux
    port map (
            O => \N__11029\,
            I => \N__11022\
        );

    \I__1496\ : Span4Mux_s0_h
    port map (
            O => \N__11026\,
            I => \N__11018\
        );

    \I__1495\ : IoInMux
    port map (
            O => \N__11025\,
            I => \N__11015\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__11022\,
            I => \N__11012\
        );

    \I__1493\ : InMux
    port map (
            O => \N__11021\,
            I => \N__11009\
        );

    \I__1492\ : Sp12to4
    port map (
            O => \N__11018\,
            I => \N__11006\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__11015\,
            I => \N__11003\
        );

    \I__1490\ : Span4Mux_v
    port map (
            O => \N__11012\,
            I => \N__10998\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__11009\,
            I => \N__10998\
        );

    \I__1488\ : Span12Mux_v
    port map (
            O => \N__11006\,
            I => \N__10995\
        );

    \I__1487\ : Span4Mux_s0_h
    port map (
            O => \N__11003\,
            I => \N__10990\
        );

    \I__1486\ : Span4Mux_h
    port map (
            O => \N__10998\,
            I => \N__10990\
        );

    \I__1485\ : Odrv12
    port map (
            O => \N__10995\,
            I => pch_pwrok
        );

    \I__1484\ : Odrv4
    port map (
            O => \N__10990\,
            I => pch_pwrok
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__10985\,
            I => \N__10982\
        );

    \I__1482\ : InMux
    port map (
            O => \N__10982\,
            I => \N__10979\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__10979\,
            I => \HDA_STRAP.m14_ns_1\
        );

    \I__1480\ : InMux
    port map (
            O => \N__10976\,
            I => \POWERLED.mult1_un54_sum_cry_2\
        );

    \I__1479\ : InMux
    port map (
            O => \N__10973\,
            I => \POWERLED.mult1_un54_sum_cry_3\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10970\,
            I => \POWERLED.mult1_un54_sum_cry_4\
        );

    \I__1477\ : InMux
    port map (
            O => \N__10967\,
            I => \N__10964\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__10964\,
            I => \N__10961\
        );

    \I__1475\ : Odrv12
    port map (
            O => \N__10961\,
            I => \POWERLED.un1_count_2_9\
        );

    \I__1474\ : CascadeMux
    port map (
            O => \N__10958\,
            I => \N__10955\
        );

    \I__1473\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10952\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__10952\,
            I => \POWERLED.count_i_9\
        );

    \I__1471\ : InMux
    port map (
            O => \N__10949\,
            I => \N__10946\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__10946\,
            I => \POWERLED.un1_count_2_10\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__10943\,
            I => \N__10940\
        );

    \I__1468\ : InMux
    port map (
            O => \N__10940\,
            I => \N__10937\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__10937\,
            I => \POWERLED.count_i_10\
        );

    \I__1466\ : InMux
    port map (
            O => \N__10934\,
            I => \N__10931\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__10931\,
            I => \N__10928\
        );

    \I__1464\ : Odrv12
    port map (
            O => \N__10928\,
            I => \POWERLED.un1_count_2_11\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__10925\,
            I => \N__10922\
        );

    \I__1462\ : InMux
    port map (
            O => \N__10922\,
            I => \N__10919\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__10919\,
            I => \POWERLED.count_i_11\
        );

    \I__1460\ : InMux
    port map (
            O => \N__10916\,
            I => \N__10913\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__10913\,
            I => \N__10910\
        );

    \I__1458\ : Span4Mux_v
    port map (
            O => \N__10910\,
            I => \N__10907\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__10907\,
            I => \POWERLED.un1_count_2_12\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__10904\,
            I => \N__10901\
        );

    \I__1455\ : InMux
    port map (
            O => \N__10901\,
            I => \N__10898\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__10898\,
            I => \N__10895\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__10895\,
            I => \POWERLED.count_i_12\
        );

    \I__1452\ : InMux
    port map (
            O => \N__10892\,
            I => \N__10889\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__10889\,
            I => \N__10886\
        );

    \I__1450\ : Span12Mux_s4_v
    port map (
            O => \N__10886\,
            I => \N__10883\
        );

    \I__1449\ : Odrv12
    port map (
            O => \N__10883\,
            I => \POWERLED.un1_count_2_13\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__10880\,
            I => \N__10877\
        );

    \I__1447\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10874\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__10874\,
            I => \POWERLED.count_i_13\
        );

    \I__1445\ : InMux
    port map (
            O => \N__10871\,
            I => \N__10868\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__10868\,
            I => \N__10865\
        );

    \I__1443\ : Span4Mux_v
    port map (
            O => \N__10865\,
            I => \N__10862\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__10862\,
            I => \POWERLED.un1_count_2_14\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__10859\,
            I => \N__10856\
        );

    \I__1440\ : InMux
    port map (
            O => \N__10856\,
            I => \N__10853\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__10853\,
            I => \N__10850\
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__10850\,
            I => \POWERLED.count_i_14\
        );

    \I__1437\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10844\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__10844\,
            I => \N__10841\
        );

    \I__1435\ : Span4Mux_s3_v
    port map (
            O => \N__10841\,
            I => \N__10838\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__10838\,
            I => \POWERLED.un1_count_2_15\
        );

    \I__1433\ : CascadeMux
    port map (
            O => \N__10835\,
            I => \N__10832\
        );

    \I__1432\ : InMux
    port map (
            O => \N__10832\,
            I => \N__10829\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__10829\,
            I => \POWERLED.count_i_15\
        );

    \I__1430\ : InMux
    port map (
            O => \N__10826\,
            I => \bfn_2_15_0_\
        );

    \I__1429\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10820\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__10820\,
            I => \POWERLED.un1_count_2_cry_15_THRU_CO\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__10817\,
            I => \N__10814\
        );

    \I__1426\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10811\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__10811\,
            I => \POWERLED.un1_count_2_1\
        );

    \I__1424\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10805\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__10805\,
            I => \N__10802\
        );

    \I__1422\ : Odrv4
    port map (
            O => \N__10802\,
            I => \POWERLED.count_i_1\
        );

    \I__1421\ : InMux
    port map (
            O => \N__10799\,
            I => \N__10796\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__10796\,
            I => \POWERLED.un1_count_2_2\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__10793\,
            I => \N__10790\
        );

    \I__1418\ : InMux
    port map (
            O => \N__10790\,
            I => \N__10787\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__10787\,
            I => \POWERLED.count_i_2\
        );

    \I__1416\ : InMux
    port map (
            O => \N__10784\,
            I => \N__10781\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__10781\,
            I => \N__10778\
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__10778\,
            I => \POWERLED.un1_count_2_3\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__10775\,
            I => \N__10772\
        );

    \I__1412\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10769\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__10769\,
            I => \POWERLED.count_i_3\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__10766\,
            I => \N__10763\
        );

    \I__1409\ : InMux
    port map (
            O => \N__10763\,
            I => \N__10760\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__10760\,
            I => \N__10757\
        );

    \I__1407\ : Odrv4
    port map (
            O => \N__10757\,
            I => \POWERLED.count_i_4\
        );

    \I__1406\ : InMux
    port map (
            O => \N__10754\,
            I => \N__10751\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__10751\,
            I => \N__10748\
        );

    \I__1404\ : Odrv12
    port map (
            O => \N__10748\,
            I => \POWERLED.un1_count_2_5\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__10745\,
            I => \N__10742\
        );

    \I__1402\ : InMux
    port map (
            O => \N__10742\,
            I => \N__10739\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__10739\,
            I => \POWERLED.count_i_5\
        );

    \I__1400\ : InMux
    port map (
            O => \N__10736\,
            I => \N__10733\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__10733\,
            I => \N__10730\
        );

    \I__1398\ : Odrv12
    port map (
            O => \N__10730\,
            I => \POWERLED.un1_count_2_6\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__10727\,
            I => \N__10724\
        );

    \I__1396\ : InMux
    port map (
            O => \N__10724\,
            I => \N__10721\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__10721\,
            I => \N__10718\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__10718\,
            I => \POWERLED.count_i_6\
        );

    \I__1393\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10712\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__10712\,
            I => \N__10709\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__10709\,
            I => \POWERLED.un1_count_2_7\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__10706\,
            I => \N__10703\
        );

    \I__1389\ : InMux
    port map (
            O => \N__10703\,
            I => \N__10700\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__10700\,
            I => \N__10697\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__10697\,
            I => \POWERLED.count_i_7\
        );

    \I__1386\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10691\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__10691\,
            I => \N__10688\
        );

    \I__1384\ : Odrv12
    port map (
            O => \N__10688\,
            I => \POWERLED.un1_count_2_8\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__10685\,
            I => \N__10682\
        );

    \I__1382\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10679\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__10679\,
            I => \POWERLED.count_i_8\
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__10676\,
            I => \N__10673\
        );

    \I__1379\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10670\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__10670\,
            I => \POWERLED.mult1_un152_sum_cry_3_s\
        );

    \I__1377\ : InMux
    port map (
            O => \N__10667\,
            I => \POWERLED.mult1_un152_sum_cry_2\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__10664\,
            I => \N__10661\
        );

    \I__1375\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10658\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__10658\,
            I => \POWERLED.mult1_un145_sum_cry_3_s\
        );

    \I__1373\ : InMux
    port map (
            O => \N__10655\,
            I => \N__10652\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__10652\,
            I => \POWERLED.mult1_un152_sum_cry_4_s\
        );

    \I__1371\ : InMux
    port map (
            O => \N__10649\,
            I => \POWERLED.mult1_un152_sum_cry_3\
        );

    \I__1370\ : InMux
    port map (
            O => \N__10646\,
            I => \N__10643\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__10643\,
            I => \POWERLED.mult1_un145_sum_cry_4_s\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__10640\,
            I => \N__10637\
        );

    \I__1367\ : InMux
    port map (
            O => \N__10637\,
            I => \N__10634\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__10634\,
            I => \POWERLED.mult1_un152_sum_cry_5_s\
        );

    \I__1365\ : InMux
    port map (
            O => \N__10631\,
            I => \POWERLED.mult1_un152_sum_cry_4\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__10628\,
            I => \N__10623\
        );

    \I__1363\ : InMux
    port map (
            O => \N__10627\,
            I => \N__10619\
        );

    \I__1362\ : InMux
    port map (
            O => \N__10626\,
            I => \N__10614\
        );

    \I__1361\ : InMux
    port map (
            O => \N__10623\,
            I => \N__10614\
        );

    \I__1360\ : InMux
    port map (
            O => \N__10622\,
            I => \N__10611\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__10619\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__10614\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__10611\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__10604\,
            I => \N__10601\
        );

    \I__1355\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10598\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__10598\,
            I => \POWERLED.mult1_un145_sum_cry_5_s\
        );

    \I__1353\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10592\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__10592\,
            I => \POWERLED.mult1_un152_sum_cry_6_s\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10589\,
            I => \POWERLED.mult1_un152_sum_cry_5\
        );

    \I__1350\ : InMux
    port map (
            O => \N__10586\,
            I => \N__10583\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__10583\,
            I => \POWERLED.mult1_un145_sum_cry_6_s\
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__10580\,
            I => \N__10576\
        );

    \I__1347\ : CascadeMux
    port map (
            O => \N__10579\,
            I => \N__10572\
        );

    \I__1346\ : InMux
    port map (
            O => \N__10576\,
            I => \N__10565\
        );

    \I__1345\ : InMux
    port map (
            O => \N__10575\,
            I => \N__10565\
        );

    \I__1344\ : InMux
    port map (
            O => \N__10572\,
            I => \N__10565\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__10565\,
            I => \POWERLED.mult1_un145_sum_i_0_8\
        );

    \I__1342\ : InMux
    port map (
            O => \N__10562\,
            I => \N__10559\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__10559\,
            I => \POWERLED.mult1_un159_sum_axb_7\
        );

    \I__1340\ : InMux
    port map (
            O => \N__10556\,
            I => \POWERLED.mult1_un152_sum_cry_6\
        );

    \I__1339\ : InMux
    port map (
            O => \N__10553\,
            I => \N__10550\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__10550\,
            I => \POWERLED.mult1_un152_sum_axb_8\
        );

    \I__1337\ : InMux
    port map (
            O => \N__10547\,
            I => \POWERLED.mult1_un152_sum_cry_7\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__10544\,
            I => \N__10539\
        );

    \I__1335\ : InMux
    port map (
            O => \N__10543\,
            I => \N__10535\
        );

    \I__1334\ : InMux
    port map (
            O => \N__10542\,
            I => \N__10530\
        );

    \I__1333\ : InMux
    port map (
            O => \N__10539\,
            I => \N__10530\
        );

    \I__1332\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10527\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__10535\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__10530\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__10527\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__10520\,
            I => \POWERLED.mult1_un152_sum_s_8_cascade_\
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__10517\,
            I => \N__10513\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__10516\,
            I => \N__10509\
        );

    \I__1325\ : InMux
    port map (
            O => \N__10513\,
            I => \N__10502\
        );

    \I__1324\ : InMux
    port map (
            O => \N__10512\,
            I => \N__10502\
        );

    \I__1323\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10502\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__10502\,
            I => \POWERLED.mult1_un152_sum_i_0_8\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__10499\,
            I => \N__10496\
        );

    \I__1320\ : InMux
    port map (
            O => \N__10496\,
            I => \N__10493\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__10493\,
            I => \POWERLED.un1_count_2_0\
        );

    \I__1318\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10487\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__10487\,
            I => \POWERLED.count_i_0_0\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__10484\,
            I => \N__10481\
        );

    \I__1315\ : InMux
    port map (
            O => \N__10481\,
            I => \N__10478\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__10478\,
            I => \POWERLED.mult1_un138_sum_i_0_8\
        );

    \I__1313\ : InMux
    port map (
            O => \N__10475\,
            I => \POWERLED.mult1_un145_sum_cry_2\
        );

    \I__1312\ : InMux
    port map (
            O => \N__10472\,
            I => \N__10468\
        );

    \I__1311\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10465\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__10468\,
            I => \POWERLED.mult1_un138_sum_cry_3_s\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__10465\,
            I => \POWERLED.mult1_un138_sum_cry_3_s\
        );

    \I__1308\ : CascadeMux
    port map (
            O => \N__10460\,
            I => \N__10457\
        );

    \I__1307\ : InMux
    port map (
            O => \N__10457\,
            I => \N__10454\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__10454\,
            I => \POWERLED.mult1_un145_sum_axb_4_l_fx\
        );

    \I__1305\ : InMux
    port map (
            O => \N__10451\,
            I => \POWERLED.mult1_un145_sum_cry_3\
        );

    \I__1304\ : InMux
    port map (
            O => \N__10448\,
            I => \N__10445\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__10445\,
            I => \N__10442\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__10442\,
            I => \POWERLED.mult1_un138_sum_cry_4_s\
        );

    \I__1301\ : InMux
    port map (
            O => \N__10439\,
            I => \POWERLED.mult1_un145_sum_cry_4\
        );

    \I__1300\ : CascadeMux
    port map (
            O => \N__10436\,
            I => \N__10433\
        );

    \I__1299\ : InMux
    port map (
            O => \N__10433\,
            I => \N__10430\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__10430\,
            I => \POWERLED.mult1_un138_sum_cry_5_s\
        );

    \I__1297\ : InMux
    port map (
            O => \N__10427\,
            I => \POWERLED.mult1_un145_sum_cry_5\
        );

    \I__1296\ : InMux
    port map (
            O => \N__10424\,
            I => \POWERLED.mult1_un145_sum_cry_6\
        );

    \I__1295\ : InMux
    port map (
            O => \N__10421\,
            I => \N__10418\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__10418\,
            I => \POWERLED.mult1_un145_sum_axb_8\
        );

    \I__1293\ : InMux
    port map (
            O => \N__10415\,
            I => \POWERLED.mult1_un145_sum_cry_7\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__10412\,
            I => \POWERLED.mult1_un145_sum_s_8_cascade_\
        );

    \I__1291\ : InMux
    port map (
            O => \N__10409\,
            I => \N__10406\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__10406\,
            I => \N__10403\
        );

    \I__1289\ : Odrv4
    port map (
            O => \N__10403\,
            I => \POWERLED.mult1_un145_sum_i\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__10400\,
            I => \POWERLED.mult1_un117_sum_s_8_cascade_\
        );

    \I__1287\ : CascadeMux
    port map (
            O => \N__10397\,
            I => \N__10393\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__10396\,
            I => \N__10389\
        );

    \I__1285\ : InMux
    port map (
            O => \N__10393\,
            I => \N__10382\
        );

    \I__1284\ : InMux
    port map (
            O => \N__10392\,
            I => \N__10382\
        );

    \I__1283\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10382\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__10382\,
            I => \POWERLED.mult1_un117_sum_i_0_8\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__10379\,
            I => \N__10374\
        );

    \I__1280\ : InMux
    port map (
            O => \N__10378\,
            I => \N__10370\
        );

    \I__1279\ : InMux
    port map (
            O => \N__10377\,
            I => \N__10365\
        );

    \I__1278\ : InMux
    port map (
            O => \N__10374\,
            I => \N__10365\
        );

    \I__1277\ : InMux
    port map (
            O => \N__10373\,
            I => \N__10362\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__10370\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__10365\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__10362\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__10355\,
            I => \N__10350\
        );

    \I__1272\ : InMux
    port map (
            O => \N__10354\,
            I => \N__10346\
        );

    \I__1271\ : InMux
    port map (
            O => \N__10353\,
            I => \N__10341\
        );

    \I__1270\ : InMux
    port map (
            O => \N__10350\,
            I => \N__10341\
        );

    \I__1269\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10338\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__10346\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__10341\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__10338\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__1265\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10328\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__10328\,
            I => \N__10325\
        );

    \I__1263\ : Odrv4
    port map (
            O => \N__10325\,
            I => \POWERLED.mult1_un131_sum_i\
        );

    \I__1262\ : InMux
    port map (
            O => \N__10322\,
            I => \N__10318\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__10321\,
            I => \N__10314\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__10318\,
            I => \N__10310\
        );

    \I__1259\ : InMux
    port map (
            O => \N__10317\,
            I => \N__10305\
        );

    \I__1258\ : InMux
    port map (
            O => \N__10314\,
            I => \N__10305\
        );

    \I__1257\ : InMux
    port map (
            O => \N__10313\,
            I => \N__10302\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__10310\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__10305\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__10302\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1253\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10292\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__10292\,
            I => \N__10289\
        );

    \I__1251\ : Span4Mux_s1_h
    port map (
            O => \N__10289\,
            I => \N__10286\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__10286\,
            I => \POWERLED.mult1_un89_sum_i\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__10283\,
            I => \N__10280\
        );

    \I__1248\ : InMux
    port map (
            O => \N__10280\,
            I => \N__10277\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__10277\,
            I => \POWERLED.mult1_un117_sum_cry_3_s\
        );

    \I__1246\ : InMux
    port map (
            O => \N__10274\,
            I => \POWERLED.mult1_un117_sum_cry_2\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__10271\,
            I => \N__10268\
        );

    \I__1244\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10265\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__10265\,
            I => \POWERLED.mult1_un110_sum_cry_3_s\
        );

    \I__1242\ : InMux
    port map (
            O => \N__10262\,
            I => \N__10259\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__10259\,
            I => \POWERLED.mult1_un117_sum_cry_4_s\
        );

    \I__1240\ : InMux
    port map (
            O => \N__10256\,
            I => \POWERLED.mult1_un117_sum_cry_3\
        );

    \I__1239\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10250\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__10250\,
            I => \POWERLED.mult1_un110_sum_cry_4_s\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__10247\,
            I => \N__10244\
        );

    \I__1236\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10241\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__10241\,
            I => \POWERLED.mult1_un117_sum_cry_5_s\
        );

    \I__1234\ : InMux
    port map (
            O => \N__10238\,
            I => \POWERLED.mult1_un117_sum_cry_4\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__10235\,
            I => \N__10230\
        );

    \I__1232\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10226\
        );

    \I__1231\ : InMux
    port map (
            O => \N__10233\,
            I => \N__10221\
        );

    \I__1230\ : InMux
    port map (
            O => \N__10230\,
            I => \N__10221\
        );

    \I__1229\ : InMux
    port map (
            O => \N__10229\,
            I => \N__10218\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__10226\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__10221\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__10218\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__10211\,
            I => \N__10208\
        );

    \I__1224\ : InMux
    port map (
            O => \N__10208\,
            I => \N__10205\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__10205\,
            I => \POWERLED.mult1_un110_sum_cry_5_s\
        );

    \I__1222\ : InMux
    port map (
            O => \N__10202\,
            I => \N__10199\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__10199\,
            I => \POWERLED.mult1_un117_sum_cry_6_s\
        );

    \I__1220\ : InMux
    port map (
            O => \N__10196\,
            I => \POWERLED.mult1_un117_sum_cry_5\
        );

    \I__1219\ : InMux
    port map (
            O => \N__10193\,
            I => \N__10190\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__10190\,
            I => \POWERLED.mult1_un110_sum_cry_6_s\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__10187\,
            I => \N__10183\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__10186\,
            I => \N__10179\
        );

    \I__1215\ : InMux
    port map (
            O => \N__10183\,
            I => \N__10172\
        );

    \I__1214\ : InMux
    port map (
            O => \N__10182\,
            I => \N__10172\
        );

    \I__1213\ : InMux
    port map (
            O => \N__10179\,
            I => \N__10172\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__10172\,
            I => \POWERLED.mult1_un110_sum_i_0_8\
        );

    \I__1211\ : InMux
    port map (
            O => \N__10169\,
            I => \N__10166\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__10166\,
            I => \POWERLED.mult1_un124_sum_axb_8\
        );

    \I__1209\ : InMux
    port map (
            O => \N__10163\,
            I => \POWERLED.mult1_un117_sum_cry_6\
        );

    \I__1208\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10157\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__10157\,
            I => \POWERLED.mult1_un117_sum_axb_8\
        );

    \I__1206\ : InMux
    port map (
            O => \N__10154\,
            I => \POWERLED.mult1_un117_sum_cry_7\
        );

    \I__1205\ : InMux
    port map (
            O => \N__10151\,
            I => \POWERLED.mult1_un68_sum_cry_7\
        );

    \I__1204\ : CascadeMux
    port map (
            O => \N__10148\,
            I => \N__10144\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__10147\,
            I => \N__10140\
        );

    \I__1202\ : InMux
    port map (
            O => \N__10144\,
            I => \N__10133\
        );

    \I__1201\ : InMux
    port map (
            O => \N__10143\,
            I => \N__10133\
        );

    \I__1200\ : InMux
    port map (
            O => \N__10140\,
            I => \N__10133\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__10133\,
            I => \POWERLED.mult1_un68_sum_i_0_8\
        );

    \I__1198\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10126\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__10129\,
            I => \N__10122\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__10126\,
            I => \N__10118\
        );

    \I__1195\ : InMux
    port map (
            O => \N__10125\,
            I => \N__10113\
        );

    \I__1194\ : InMux
    port map (
            O => \N__10122\,
            I => \N__10113\
        );

    \I__1193\ : InMux
    port map (
            O => \N__10121\,
            I => \N__10110\
        );

    \I__1192\ : Odrv4
    port map (
            O => \N__10118\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__10113\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__10110\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__1189\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10099\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__10102\,
            I => \N__10095\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__10099\,
            I => \N__10091\
        );

    \I__1186\ : InMux
    port map (
            O => \N__10098\,
            I => \N__10086\
        );

    \I__1185\ : InMux
    port map (
            O => \N__10095\,
            I => \N__10086\
        );

    \I__1184\ : InMux
    port map (
            O => \N__10094\,
            I => \N__10083\
        );

    \I__1183\ : Odrv4
    port map (
            O => \N__10091\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__10086\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__10083\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__10076\,
            I => \N__10071\
        );

    \I__1179\ : InMux
    port map (
            O => \N__10075\,
            I => \N__10066\
        );

    \I__1178\ : InMux
    port map (
            O => \N__10074\,
            I => \N__10061\
        );

    \I__1177\ : InMux
    port map (
            O => \N__10071\,
            I => \N__10061\
        );

    \I__1176\ : InMux
    port map (
            O => \N__10070\,
            I => \N__10058\
        );

    \I__1175\ : InMux
    port map (
            O => \N__10069\,
            I => \N__10055\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__10066\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__10061\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__10058\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__10055\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__1170\ : InMux
    port map (
            O => \N__10046\,
            I => \N__10042\
        );

    \I__1169\ : CascadeMux
    port map (
            O => \N__10045\,
            I => \N__10038\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__10042\,
            I => \N__10034\
        );

    \I__1167\ : InMux
    port map (
            O => \N__10041\,
            I => \N__10029\
        );

    \I__1166\ : InMux
    port map (
            O => \N__10038\,
            I => \N__10029\
        );

    \I__1165\ : InMux
    port map (
            O => \N__10037\,
            I => \N__10026\
        );

    \I__1164\ : Odrv4
    port map (
            O => \N__10034\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__10029\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__10026\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__1161\ : InMux
    port map (
            O => \N__10019\,
            I => \N__10016\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__10016\,
            I => \POWERLED.mult1_un103_sum_i\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__10013\,
            I => \N__10008\
        );

    \I__1158\ : InMux
    port map (
            O => \N__10012\,
            I => \N__10004\
        );

    \I__1157\ : InMux
    port map (
            O => \N__10011\,
            I => \N__9999\
        );

    \I__1156\ : InMux
    port map (
            O => \N__10008\,
            I => \N__9999\
        );

    \I__1155\ : InMux
    port map (
            O => \N__10007\,
            I => \N__9996\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__10004\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__9999\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__9996\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1151\ : InMux
    port map (
            O => \N__9989\,
            I => \N__9986\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__9986\,
            I => \POWERLED.mult1_un82_sum_axb_8\
        );

    \I__1149\ : InMux
    port map (
            O => \N__9983\,
            I => \POWERLED.mult1_un75_sum_cry_6\
        );

    \I__1148\ : InMux
    port map (
            O => \N__9980\,
            I => \POWERLED.mult1_un75_sum_cry_7\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__9977\,
            I => \POWERLED.mult1_un75_sum_s_8_cascade_\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__9974\,
            I => \N__9970\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__9973\,
            I => \N__9966\
        );

    \I__1144\ : InMux
    port map (
            O => \N__9970\,
            I => \N__9959\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9969\,
            I => \N__9959\
        );

    \I__1142\ : InMux
    port map (
            O => \N__9966\,
            I => \N__9959\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__9959\,
            I => \POWERLED.mult1_un75_sum_i_0_8\
        );

    \I__1140\ : CascadeMux
    port map (
            O => \N__9956\,
            I => \N__9953\
        );

    \I__1139\ : InMux
    port map (
            O => \N__9953\,
            I => \N__9950\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__9950\,
            I => \POWERLED.mult1_un68_sum_cry_3_s\
        );

    \I__1137\ : InMux
    port map (
            O => \N__9947\,
            I => \POWERLED.mult1_un68_sum_cry_2\
        );

    \I__1136\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9941\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__9941\,
            I => \POWERLED.mult1_un68_sum_cry_4_s\
        );

    \I__1134\ : InMux
    port map (
            O => \N__9938\,
            I => \POWERLED.mult1_un68_sum_cry_3\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__9935\,
            I => \N__9932\
        );

    \I__1132\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9929\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__9929\,
            I => \POWERLED.mult1_un68_sum_cry_5_s\
        );

    \I__1130\ : InMux
    port map (
            O => \N__9926\,
            I => \POWERLED.mult1_un68_sum_cry_4\
        );

    \I__1129\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9920\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__9920\,
            I => \POWERLED.mult1_un68_sum_cry_6_s\
        );

    \I__1127\ : InMux
    port map (
            O => \N__9917\,
            I => \POWERLED.mult1_un68_sum_cry_5\
        );

    \I__1126\ : InMux
    port map (
            O => \N__9914\,
            I => \N__9911\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__9911\,
            I => \POWERLED.mult1_un75_sum_axb_8\
        );

    \I__1124\ : InMux
    port map (
            O => \N__9908\,
            I => \POWERLED.mult1_un68_sum_cry_6\
        );

    \I__1123\ : InMux
    port map (
            O => \N__9905\,
            I => \N__9902\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__9902\,
            I => \POWERLED.mult1_un89_sum_axb_8\
        );

    \I__1121\ : InMux
    port map (
            O => \N__9899\,
            I => \POWERLED.mult1_un82_sum_cry_6\
        );

    \I__1120\ : InMux
    port map (
            O => \N__9896\,
            I => \POWERLED.mult1_un82_sum_cry_7\
        );

    \I__1119\ : CascadeMux
    port map (
            O => \N__9893\,
            I => \POWERLED.mult1_un82_sum_s_8_cascade_\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__9890\,
            I => \N__9886\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__9889\,
            I => \N__9882\
        );

    \I__1116\ : InMux
    port map (
            O => \N__9886\,
            I => \N__9875\
        );

    \I__1115\ : InMux
    port map (
            O => \N__9885\,
            I => \N__9875\
        );

    \I__1114\ : InMux
    port map (
            O => \N__9882\,
            I => \N__9875\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__9875\,
            I => \POWERLED.mult1_un82_sum_i_0_8\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__9872\,
            I => \N__9869\
        );

    \I__1111\ : InMux
    port map (
            O => \N__9869\,
            I => \N__9866\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__9866\,
            I => \POWERLED.mult1_un75_sum_cry_3_s\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9863\,
            I => \POWERLED.mult1_un75_sum_cry_2\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9857\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__9857\,
            I => \POWERLED.mult1_un75_sum_cry_4_s\
        );

    \I__1106\ : InMux
    port map (
            O => \N__9854\,
            I => \POWERLED.mult1_un75_sum_cry_3\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__9851\,
            I => \N__9848\
        );

    \I__1104\ : InMux
    port map (
            O => \N__9848\,
            I => \N__9845\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__9845\,
            I => \POWERLED.mult1_un75_sum_cry_5_s\
        );

    \I__1102\ : InMux
    port map (
            O => \N__9842\,
            I => \POWERLED.mult1_un75_sum_cry_4\
        );

    \I__1101\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9836\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__9836\,
            I => \POWERLED.mult1_un75_sum_cry_6_s\
        );

    \I__1099\ : InMux
    port map (
            O => \N__9833\,
            I => \POWERLED.mult1_un75_sum_cry_5\
        );

    \I__1098\ : InMux
    port map (
            O => \N__9830\,
            I => \N__9826\
        );

    \I__1097\ : InMux
    port map (
            O => \N__9829\,
            I => \N__9823\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__9826\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__9823\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__1094\ : InMux
    port map (
            O => \N__9818\,
            I => \PCH_PWRGD.un1_count_1_cry_12\
        );

    \I__1093\ : InMux
    port map (
            O => \N__9815\,
            I => \N__9811\
        );

    \I__1092\ : InMux
    port map (
            O => \N__9814\,
            I => \N__9808\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__9811\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__9808\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__1089\ : InMux
    port map (
            O => \N__9803\,
            I => \PCH_PWRGD.un1_count_1_cry_13\
        );

    \I__1088\ : InMux
    port map (
            O => \N__9800\,
            I => \bfn_2_4_0_\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__9797\,
            I => \N__9793\
        );

    \I__1086\ : InMux
    port map (
            O => \N__9796\,
            I => \N__9790\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9787\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__9790\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__9787\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__1082\ : CEMux
    port map (
            O => \N__9782\,
            I => \N__9779\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__9779\,
            I => \N__9776\
        );

    \I__1080\ : Span4Mux_v
    port map (
            O => \N__9776\,
            I => \N__9773\
        );

    \I__1079\ : Odrv4
    port map (
            O => \N__9773\,
            I => \PCH_PWRGD.N_65_3\
        );

    \I__1078\ : SRMux
    port map (
            O => \N__9770\,
            I => \N__9765\
        );

    \I__1077\ : SRMux
    port map (
            O => \N__9769\,
            I => \N__9762\
        );

    \I__1076\ : SRMux
    port map (
            O => \N__9768\,
            I => \N__9759\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__9765\,
            I => \PCH_PWRGD.curr_state_RNI7N705Z0Z_0\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__9762\,
            I => \PCH_PWRGD.curr_state_RNI7N705Z0Z_0\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__9759\,
            I => \PCH_PWRGD.curr_state_RNI7N705Z0Z_0\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__9752\,
            I => \N__9749\
        );

    \I__1071\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9746\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__9746\,
            I => \POWERLED.mult1_un82_sum_cry_3_s\
        );

    \I__1069\ : InMux
    port map (
            O => \N__9743\,
            I => \POWERLED.mult1_un82_sum_cry_2\
        );

    \I__1068\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9737\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__9737\,
            I => \POWERLED.mult1_un82_sum_cry_4_s\
        );

    \I__1066\ : InMux
    port map (
            O => \N__9734\,
            I => \POWERLED.mult1_un82_sum_cry_3\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__9731\,
            I => \N__9728\
        );

    \I__1064\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9725\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__9725\,
            I => \POWERLED.mult1_un82_sum_cry_5_s\
        );

    \I__1062\ : InMux
    port map (
            O => \N__9722\,
            I => \POWERLED.mult1_un82_sum_cry_4\
        );

    \I__1061\ : InMux
    port map (
            O => \N__9719\,
            I => \N__9716\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__9716\,
            I => \POWERLED.mult1_un82_sum_cry_6_s\
        );

    \I__1059\ : InMux
    port map (
            O => \N__9713\,
            I => \POWERLED.mult1_un82_sum_cry_5\
        );

    \I__1058\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9706\
        );

    \I__1057\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9703\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__9706\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__9703\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__1054\ : InMux
    port map (
            O => \N__9698\,
            I => \PCH_PWRGD.un1_count_1_cry_4\
        );

    \I__1053\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9691\
        );

    \I__1052\ : InMux
    port map (
            O => \N__9694\,
            I => \N__9688\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__9691\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__9688\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__1049\ : InMux
    port map (
            O => \N__9683\,
            I => \PCH_PWRGD.un1_count_1_cry_5\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__9680\,
            I => \N__9676\
        );

    \I__1047\ : InMux
    port map (
            O => \N__9679\,
            I => \N__9673\
        );

    \I__1046\ : InMux
    port map (
            O => \N__9676\,
            I => \N__9670\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__9673\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__9670\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__1043\ : InMux
    port map (
            O => \N__9665\,
            I => \PCH_PWRGD.un1_count_1_cry_6\
        );

    \I__1042\ : InMux
    port map (
            O => \N__9662\,
            I => \N__9658\
        );

    \I__1041\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9655\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__9658\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__9655\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__1038\ : InMux
    port map (
            O => \N__9650\,
            I => \bfn_2_3_0_\
        );

    \I__1037\ : InMux
    port map (
            O => \N__9647\,
            I => \N__9643\
        );

    \I__1036\ : InMux
    port map (
            O => \N__9646\,
            I => \N__9640\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__9643\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__9640\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__1033\ : InMux
    port map (
            O => \N__9635\,
            I => \PCH_PWRGD.un1_count_1_cry_8\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__9632\,
            I => \N__9628\
        );

    \I__1031\ : InMux
    port map (
            O => \N__9631\,
            I => \N__9625\
        );

    \I__1030\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9622\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__9625\,
            I => \PCH_PWRGD.countZ0Z_10\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__9622\,
            I => \PCH_PWRGD.countZ0Z_10\
        );

    \I__1027\ : InMux
    port map (
            O => \N__9617\,
            I => \PCH_PWRGD.un1_count_1_cry_9\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__9614\,
            I => \N__9610\
        );

    \I__1025\ : InMux
    port map (
            O => \N__9613\,
            I => \N__9607\
        );

    \I__1024\ : InMux
    port map (
            O => \N__9610\,
            I => \N__9604\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__9607\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__9604\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__1021\ : InMux
    port map (
            O => \N__9599\,
            I => \PCH_PWRGD.un1_count_1_cry_10\
        );

    \I__1020\ : InMux
    port map (
            O => \N__9596\,
            I => \N__9592\
        );

    \I__1019\ : InMux
    port map (
            O => \N__9595\,
            I => \N__9589\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__9592\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__9589\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__1016\ : InMux
    port map (
            O => \N__9584\,
            I => \PCH_PWRGD.un1_count_1_cry_11\
        );

    \I__1015\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9578\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__9578\,
            I => \N__9575\
        );

    \I__1013\ : Odrv12
    port map (
            O => \N__9575\,
            I => \POWERLED.mult1_un96_sum_i\
        );

    \I__1012\ : InMux
    port map (
            O => \N__9572\,
            I => \N__9569\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__9569\,
            I => \N__9565\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__9568\,
            I => \N__9561\
        );

    \I__1009\ : Span12Mux_s4_v
    port map (
            O => \N__9565\,
            I => \N__9557\
        );

    \I__1008\ : InMux
    port map (
            O => \N__9564\,
            I => \N__9552\
        );

    \I__1007\ : InMux
    port map (
            O => \N__9561\,
            I => \N__9552\
        );

    \I__1006\ : InMux
    port map (
            O => \N__9560\,
            I => \N__9549\
        );

    \I__1005\ : Odrv12
    port map (
            O => \N__9557\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__9552\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__9549\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__1002\ : IoInMux
    port map (
            O => \N__9542\,
            I => \N__9539\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__9539\,
            I => \N__9536\
        );

    \I__1000\ : Odrv4
    port map (
            O => \N__9536\,
            I => pwrbtn_led
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__9533\,
            I => \N__9529\
        );

    \I__998\ : InMux
    port map (
            O => \N__9532\,
            I => \N__9526\
        );

    \I__997\ : InMux
    port map (
            O => \N__9529\,
            I => \N__9523\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__9526\,
            I => \N__9518\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__9523\,
            I => \N__9518\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__9518\,
            I => \PCH_PWRGD.un1_curr_state10_0\
        );

    \I__993\ : InMux
    port map (
            O => \N__9515\,
            I => \N__9511\
        );

    \I__992\ : InMux
    port map (
            O => \N__9514\,
            I => \N__9508\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__9511\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__9508\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__989\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9499\
        );

    \I__988\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9496\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__9499\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__9496\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__985\ : InMux
    port map (
            O => \N__9491\,
            I => \PCH_PWRGD.un1_count_1_cry_0\
        );

    \I__984\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9484\
        );

    \I__983\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9481\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__9484\,
            I => \PCH_PWRGD.countZ0Z_2\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__9481\,
            I => \PCH_PWRGD.countZ0Z_2\
        );

    \I__980\ : InMux
    port map (
            O => \N__9476\,
            I => \PCH_PWRGD.un1_count_1_cry_1\
        );

    \I__979\ : InMux
    port map (
            O => \N__9473\,
            I => \N__9469\
        );

    \I__978\ : InMux
    port map (
            O => \N__9472\,
            I => \N__9466\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__9469\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__9466\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__975\ : InMux
    port map (
            O => \N__9461\,
            I => \PCH_PWRGD.un1_count_1_cry_2\
        );

    \I__974\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9454\
        );

    \I__973\ : InMux
    port map (
            O => \N__9457\,
            I => \N__9451\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__9454\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__9451\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__970\ : InMux
    port map (
            O => \N__9446\,
            I => \PCH_PWRGD.un1_count_1_cry_3\
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__9443\,
            I => \N__9440\
        );

    \I__968\ : InMux
    port map (
            O => \N__9440\,
            I => \N__9437\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__9437\,
            I => \POWERLED.mult1_un159_sum_cry_2_s\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__9434\,
            I => \N__9431\
        );

    \I__965\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__9428\,
            I => \POWERLED.mult1_un159_sum_cry_3_s\
        );

    \I__963\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9422\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__9422\,
            I => \POWERLED.mult1_un159_sum_cry_4_s\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__9419\,
            I => \N__9415\
        );

    \I__960\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9410\
        );

    \I__959\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9403\
        );

    \I__958\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9403\
        );

    \I__957\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9403\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__9410\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__9403\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__954\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9395\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__9395\,
            I => \POWERLED.mult1_un159_sum_cry_5_s\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__9392\,
            I => \N__9388\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__9391\,
            I => \N__9384\
        );

    \I__950\ : InMux
    port map (
            O => \N__9388\,
            I => \N__9377\
        );

    \I__949\ : InMux
    port map (
            O => \N__9387\,
            I => \N__9377\
        );

    \I__948\ : InMux
    port map (
            O => \N__9384\,
            I => \N__9377\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__9377\,
            I => \G_407\
        );

    \I__946\ : InMux
    port map (
            O => \N__9374\,
            I => \N__9371\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__9371\,
            I => \POWERLED.mult1_un166_sum_axb_6\
        );

    \I__944\ : InMux
    port map (
            O => \N__9368\,
            I => \POWERLED.mult1_un166_sum_cry_5\
        );

    \I__943\ : InMux
    port map (
            O => \N__9365\,
            I => \POWERLED.mult1_un138_sum_cry_7\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__9362\,
            I => \POWERLED.mult1_un138_sum_s_8_cascade_\
        );

    \I__941\ : InMux
    port map (
            O => \N__9359\,
            I => \POWERLED.mult1_un159_sum_cry_1\
        );

    \I__940\ : InMux
    port map (
            O => \N__9356\,
            I => \POWERLED.mult1_un159_sum_cry_2\
        );

    \I__939\ : InMux
    port map (
            O => \N__9353\,
            I => \POWERLED.mult1_un159_sum_cry_3\
        );

    \I__938\ : InMux
    port map (
            O => \N__9350\,
            I => \POWERLED.mult1_un159_sum_cry_4\
        );

    \I__937\ : InMux
    port map (
            O => \N__9347\,
            I => \POWERLED.mult1_un159_sum_cry_5\
        );

    \I__936\ : InMux
    port map (
            O => \N__9344\,
            I => \POWERLED.mult1_un159_sum_cry_6\
        );

    \I__935\ : CascadeMux
    port map (
            O => \N__9341\,
            I => \POWERLED.mult1_un159_sum_s_7_cascade_\
        );

    \I__934\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9335\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__9335\,
            I => \POWERLED.mult1_un131_sum_axb_8\
        );

    \I__932\ : InMux
    port map (
            O => \N__9332\,
            I => \POWERLED.mult1_un131_sum_cry_7\
        );

    \I__931\ : CascadeMux
    port map (
            O => \N__9329\,
            I => \POWERLED.mult1_un131_sum_s_8_cascade_\
        );

    \I__930\ : InMux
    port map (
            O => \N__9326\,
            I => \POWERLED.mult1_un138_sum_cry_2\
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__9323\,
            I => \N__9320\
        );

    \I__928\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9317\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__9317\,
            I => \POWERLED.mult1_un131_sum_cry_3_s\
        );

    \I__926\ : InMux
    port map (
            O => \N__9314\,
            I => \POWERLED.mult1_un138_sum_cry_3\
        );

    \I__925\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9308\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__9308\,
            I => \POWERLED.mult1_un131_sum_cry_4_s\
        );

    \I__923\ : InMux
    port map (
            O => \N__9305\,
            I => \POWERLED.mult1_un138_sum_cry_4\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__9302\,
            I => \N__9299\
        );

    \I__921\ : InMux
    port map (
            O => \N__9299\,
            I => \N__9296\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__9296\,
            I => \POWERLED.mult1_un131_sum_cry_5_s\
        );

    \I__919\ : InMux
    port map (
            O => \N__9293\,
            I => \POWERLED.mult1_un138_sum_cry_5\
        );

    \I__918\ : InMux
    port map (
            O => \N__9290\,
            I => \N__9287\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__9287\,
            I => \POWERLED.mult1_un131_sum_cry_6_s\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__9284\,
            I => \N__9280\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__9283\,
            I => \N__9276\
        );

    \I__914\ : InMux
    port map (
            O => \N__9280\,
            I => \N__9269\
        );

    \I__913\ : InMux
    port map (
            O => \N__9279\,
            I => \N__9269\
        );

    \I__912\ : InMux
    port map (
            O => \N__9276\,
            I => \N__9269\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__9269\,
            I => \POWERLED.mult1_un131_sum_i_0_8\
        );

    \I__910\ : InMux
    port map (
            O => \N__9266\,
            I => \POWERLED.mult1_un138_sum_cry_6\
        );

    \I__909\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__9260\,
            I => \POWERLED.mult1_un138_sum_axb_8\
        );

    \I__907\ : InMux
    port map (
            O => \N__9257\,
            I => \POWERLED.mult1_un124_sum_cry_6\
        );

    \I__906\ : InMux
    port map (
            O => \N__9254\,
            I => \POWERLED.mult1_un124_sum_cry_7\
        );

    \I__905\ : CascadeMux
    port map (
            O => \N__9251\,
            I => \POWERLED.mult1_un124_sum_s_8_cascade_\
        );

    \I__904\ : InMux
    port map (
            O => \N__9248\,
            I => \POWERLED.mult1_un131_sum_cry_2\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__9245\,
            I => \N__9242\
        );

    \I__902\ : InMux
    port map (
            O => \N__9242\,
            I => \N__9239\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__9239\,
            I => \POWERLED.mult1_un124_sum_cry_3_s\
        );

    \I__900\ : InMux
    port map (
            O => \N__9236\,
            I => \POWERLED.mult1_un131_sum_cry_3\
        );

    \I__899\ : InMux
    port map (
            O => \N__9233\,
            I => \N__9230\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__9230\,
            I => \POWERLED.mult1_un124_sum_cry_4_s\
        );

    \I__897\ : InMux
    port map (
            O => \N__9227\,
            I => \POWERLED.mult1_un131_sum_cry_4\
        );

    \I__896\ : CascadeMux
    port map (
            O => \N__9224\,
            I => \N__9221\
        );

    \I__895\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9218\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__9218\,
            I => \POWERLED.mult1_un124_sum_cry_5_s\
        );

    \I__893\ : InMux
    port map (
            O => \N__9215\,
            I => \POWERLED.mult1_un131_sum_cry_5\
        );

    \I__892\ : InMux
    port map (
            O => \N__9212\,
            I => \N__9209\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__9209\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__9206\,
            I => \N__9202\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__9205\,
            I => \N__9198\
        );

    \I__888\ : InMux
    port map (
            O => \N__9202\,
            I => \N__9191\
        );

    \I__887\ : InMux
    port map (
            O => \N__9201\,
            I => \N__9191\
        );

    \I__886\ : InMux
    port map (
            O => \N__9198\,
            I => \N__9191\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__9191\,
            I => \POWERLED.mult1_un124_sum_i_0_8\
        );

    \I__884\ : InMux
    port map (
            O => \N__9188\,
            I => \POWERLED.mult1_un131_sum_cry_6\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__9185\,
            I => \N__9182\
        );

    \I__882\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9179\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__9179\,
            I => \POWERLED.mult1_un103_sum_cry_5_s\
        );

    \I__880\ : InMux
    port map (
            O => \N__9176\,
            I => \POWERLED.mult1_un110_sum_cry_5\
        );

    \I__879\ : InMux
    port map (
            O => \N__9173\,
            I => \N__9170\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__9170\,
            I => \POWERLED.mult1_un103_sum_cry_6_s\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__9167\,
            I => \N__9163\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__9166\,
            I => \N__9159\
        );

    \I__875\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9152\
        );

    \I__874\ : InMux
    port map (
            O => \N__9162\,
            I => \N__9152\
        );

    \I__873\ : InMux
    port map (
            O => \N__9159\,
            I => \N__9152\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__9152\,
            I => \POWERLED.mult1_un103_sum_i_0_8\
        );

    \I__871\ : InMux
    port map (
            O => \N__9149\,
            I => \POWERLED.mult1_un110_sum_cry_6\
        );

    \I__870\ : InMux
    port map (
            O => \N__9146\,
            I => \N__9143\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__9143\,
            I => \POWERLED.mult1_un110_sum_axb_8\
        );

    \I__868\ : InMux
    port map (
            O => \N__9140\,
            I => \POWERLED.mult1_un110_sum_cry_7\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__9137\,
            I => \POWERLED.mult1_un110_sum_s_8_cascade_\
        );

    \I__866\ : InMux
    port map (
            O => \N__9134\,
            I => \POWERLED.mult1_un124_sum_cry_2\
        );

    \I__865\ : InMux
    port map (
            O => \N__9131\,
            I => \POWERLED.mult1_un124_sum_cry_3\
        );

    \I__864\ : InMux
    port map (
            O => \N__9128\,
            I => \POWERLED.mult1_un124_sum_cry_4\
        );

    \I__863\ : InMux
    port map (
            O => \N__9125\,
            I => \POWERLED.mult1_un124_sum_cry_5\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__861\ : InMux
    port map (
            O => \N__9119\,
            I => \N__9116\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__9116\,
            I => \POWERLED.mult1_un96_sum_cry_5_s\
        );

    \I__859\ : InMux
    port map (
            O => \N__9113\,
            I => \POWERLED.mult1_un103_sum_cry_5\
        );

    \I__858\ : InMux
    port map (
            O => \N__9110\,
            I => \N__9107\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__9107\,
            I => \POWERLED.mult1_un96_sum_cry_6_s\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__9104\,
            I => \N__9100\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__9103\,
            I => \N__9096\
        );

    \I__854\ : InMux
    port map (
            O => \N__9100\,
            I => \N__9089\
        );

    \I__853\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9089\
        );

    \I__852\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9089\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__9089\,
            I => \POWERLED.mult1_un96_sum_i_0_8\
        );

    \I__850\ : InMux
    port map (
            O => \N__9086\,
            I => \POWERLED.mult1_un103_sum_cry_6\
        );

    \I__849\ : InMux
    port map (
            O => \N__9083\,
            I => \N__9080\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__9080\,
            I => \POWERLED.mult1_un103_sum_axb_8\
        );

    \I__847\ : InMux
    port map (
            O => \N__9077\,
            I => \POWERLED.mult1_un103_sum_cry_7\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__9074\,
            I => \POWERLED.mult1_un103_sum_s_8_cascade_\
        );

    \I__845\ : InMux
    port map (
            O => \N__9071\,
            I => \POWERLED.mult1_un110_sum_cry_2\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__9068\,
            I => \N__9065\
        );

    \I__843\ : InMux
    port map (
            O => \N__9065\,
            I => \N__9062\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__9062\,
            I => \POWERLED.mult1_un103_sum_cry_3_s\
        );

    \I__841\ : InMux
    port map (
            O => \N__9059\,
            I => \POWERLED.mult1_un110_sum_cry_3\
        );

    \I__840\ : InMux
    port map (
            O => \N__9056\,
            I => \N__9053\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__9053\,
            I => \POWERLED.mult1_un103_sum_cry_4_s\
        );

    \I__838\ : InMux
    port map (
            O => \N__9050\,
            I => \POWERLED.mult1_un110_sum_cry_4\
        );

    \I__837\ : InMux
    port map (
            O => \N__9047\,
            I => \N__9044\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__9044\,
            I => \POWERLED.mult1_un89_sum_cry_4_s\
        );

    \I__835\ : InMux
    port map (
            O => \N__9041\,
            I => \POWERLED.mult1_un96_sum_cry_4\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__833\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__9032\,
            I => \POWERLED.mult1_un89_sum_cry_5_s\
        );

    \I__831\ : InMux
    port map (
            O => \N__9029\,
            I => \POWERLED.mult1_un96_sum_cry_5\
        );

    \I__830\ : InMux
    port map (
            O => \N__9026\,
            I => \N__9023\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__9023\,
            I => \POWERLED.mult1_un89_sum_cry_6_s\
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__9020\,
            I => \N__9016\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__9019\,
            I => \N__9012\
        );

    \I__826\ : InMux
    port map (
            O => \N__9016\,
            I => \N__9005\
        );

    \I__825\ : InMux
    port map (
            O => \N__9015\,
            I => \N__9005\
        );

    \I__824\ : InMux
    port map (
            O => \N__9012\,
            I => \N__9005\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__9005\,
            I => \POWERLED.mult1_un89_sum_i_0_8\
        );

    \I__822\ : InMux
    port map (
            O => \N__9002\,
            I => \POWERLED.mult1_un96_sum_cry_6\
        );

    \I__821\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8996\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__8996\,
            I => \POWERLED.mult1_un96_sum_axb_8\
        );

    \I__819\ : InMux
    port map (
            O => \N__8993\,
            I => \POWERLED.mult1_un96_sum_cry_7\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__8990\,
            I => \POWERLED.mult1_un96_sum_s_8_cascade_\
        );

    \I__817\ : InMux
    port map (
            O => \N__8987\,
            I => \POWERLED.mult1_un103_sum_cry_2\
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__815\ : InMux
    port map (
            O => \N__8981\,
            I => \N__8978\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__8978\,
            I => \POWERLED.mult1_un96_sum_cry_3_s\
        );

    \I__813\ : InMux
    port map (
            O => \N__8975\,
            I => \POWERLED.mult1_un103_sum_cry_3\
        );

    \I__812\ : InMux
    port map (
            O => \N__8972\,
            I => \N__8969\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__8969\,
            I => \POWERLED.mult1_un96_sum_cry_4_s\
        );

    \I__810\ : InMux
    port map (
            O => \N__8966\,
            I => \POWERLED.mult1_un103_sum_cry_4\
        );

    \I__809\ : InMux
    port map (
            O => \N__8963\,
            I => \POWERLED.mult1_un89_sum_cry_3\
        );

    \I__808\ : InMux
    port map (
            O => \N__8960\,
            I => \POWERLED.mult1_un89_sum_cry_4\
        );

    \I__807\ : InMux
    port map (
            O => \N__8957\,
            I => \POWERLED.mult1_un89_sum_cry_5\
        );

    \I__806\ : InMux
    port map (
            O => \N__8954\,
            I => \POWERLED.mult1_un89_sum_cry_6\
        );

    \I__805\ : InMux
    port map (
            O => \N__8951\,
            I => \POWERLED.mult1_un89_sum_cry_7\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__8948\,
            I => \POWERLED.mult1_un89_sum_s_8_cascade_\
        );

    \I__803\ : InMux
    port map (
            O => \N__8945\,
            I => \POWERLED.mult1_un96_sum_cry_2\
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__801\ : InMux
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__8936\,
            I => \POWERLED.mult1_un89_sum_cry_3_s\
        );

    \I__799\ : InMux
    port map (
            O => \N__8933\,
            I => \POWERLED.mult1_un96_sum_cry_3\
        );

    \I__798\ : CascadeMux
    port map (
            O => \N__8930\,
            I => \PCH_PWRGD.curr_state_RNI7N705Z0Z_0_cascade_\
        );

    \I__797\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8924\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__8924\,
            I => \PCH_PWRGD.un4_count_8\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__8921\,
            I => \PCH_PWRGD.N_3_i_cascade_\
        );

    \I__794\ : InMux
    port map (
            O => \N__8918\,
            I => \N__8912\
        );

    \I__793\ : InMux
    port map (
            O => \N__8917\,
            I => \N__8912\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__8912\,
            I => \N__8909\
        );

    \I__791\ : Span4Mux_v
    port map (
            O => \N__8909\,
            I => \N__8906\
        );

    \I__790\ : Span4Mux_v
    port map (
            O => \N__8906\,
            I => \N__8903\
        );

    \I__789\ : Odrv4
    port map (
            O => \N__8903\,
            I => vr_ready_vccin
        );

    \I__788\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8887\
        );

    \I__787\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8887\
        );

    \I__786\ : InMux
    port map (
            O => \N__8898\,
            I => \N__8887\
        );

    \I__785\ : InMux
    port map (
            O => \N__8897\,
            I => \N__8887\
        );

    \I__784\ : InMux
    port map (
            O => \N__8896\,
            I => \N__8884\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__8887\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__8884\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__781\ : InMux
    port map (
            O => \N__8879\,
            I => \N__8873\
        );

    \I__780\ : InMux
    port map (
            O => \N__8878\,
            I => \N__8873\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__8873\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__778\ : CascadeMux
    port map (
            O => \N__8870\,
            I => \N__8866\
        );

    \I__777\ : InMux
    port map (
            O => \N__8869\,
            I => \N__8862\
        );

    \I__776\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8859\
        );

    \I__775\ : InMux
    port map (
            O => \N__8865\,
            I => \N__8856\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__8862\,
            I => \N__8853\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__8859\,
            I => \PCH_PWRGD.N_3_i\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__8856\,
            I => \PCH_PWRGD.N_3_i\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__8853\,
            I => \PCH_PWRGD.N_3_i\
        );

    \I__770\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8839\
        );

    \I__769\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8830\
        );

    \I__768\ : InMux
    port map (
            O => \N__8844\,
            I => \N__8830\
        );

    \I__767\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8830\
        );

    \I__766\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8830\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__8839\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__8830\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__763\ : InMux
    port map (
            O => \N__8825\,
            I => \POWERLED.mult1_un89_sum_cry_2\
        );

    \I__762\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__8819\,
            I => \PCH_PWRGD.un4_count_11\
        );

    \I__760\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8813\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__8813\,
            I => \PCH_PWRGD.un4_count_9\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__8810\,
            I => \PCH_PWRGD.un4_count_10_cascade_\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__8807\,
            I => \PCH_PWRGD.N_1_i_cascade_\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__8804\,
            I => \PCH_PWRGD.un1_curr_state_0_sqmuxa_0_cascade_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.dutycycle_cry_6\,
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_7_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.dutycycle_cry_14\,
            carryinitout => \bfn_7_9_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_5_0_\
        );

    \IN_MUX_bfv_2_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_5_0_\
        );

    \IN_MUX_bfv_2_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_6_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_4_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_7_0_\
        );

    \IN_MUX_bfv_4_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_5_0_\
        );

    \IN_MUX_bfv_4_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_6_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_8_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_1_cry_8\,
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_5_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO\,
            carryinitout => \bfn_5_16_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.un4_counter_7\,
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_9_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_1_0_\
        );

    \IN_MUX_bfv_9_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_8\,
            carryinitout => \bfn_9_2_0_\
        );

    \IN_MUX_bfv_9_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_16\,
            carryinitout => \bfn_9_3_0_\
        );

    \IN_MUX_bfv_9_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_24\,
            carryinitout => \bfn_9_4_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_7\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_2_cry_7\,
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_2_cry_15\,
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_1_cry_7\,
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_1_cry_15\,
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_off_1_cry_7\,
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_clk_1_cry_7\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_2_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_2_0_\
        );

    \IN_MUX_bfv_2_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_2_3_0_\
        );

    \IN_MUX_bfv_2_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_2_4_0_\
        );

    \IN_MUX_bfv_6_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_1_0_\
        );

    \IN_MUX_bfv_6_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un1_count_1_cry_7\,
            carryinitout => \bfn_6_2_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un1_count_1_cry_15\,
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALL_SYS_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_8_7_0_\
        );

    \COUNTER.tmp_RNIRH3P_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__17737\,
            GLOBALBUFFEROUTPUT => \N_65_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIESHJ_1_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9694\,
            in1 => \N__9487\,
            in2 => \N__9632\,
            in3 => \N__9502\,
            lcout => \PCH_PWRGD.un4_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI7J2B_3_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9709\,
            in1 => \N__9457\,
            in2 => \N__9680\,
            in3 => \N__9472\,
            lcout => \PCH_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIN5IJ_0_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9646\,
            in1 => \N__9514\,
            in2 => \N__9614\,
            in3 => \N__9661\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un4_count_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8822\,
            in1 => \N__8816\,
            in2 => \N__8810\,
            in3 => \N__8927\,
            lcout => \PCH_PWRGD.N_1_i\,
            ltout => \PCH_PWRGD.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIC5474_0_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011011111"
        )
    port map (
            in0 => \N__8846\,
            in1 => \N__8896\,
            in2 => \N__8807\,
            in3 => \N__8869\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un1_curr_state_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI7N705_0_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8804\,
            in3 => \N__20059\,
            lcout => \PCH_PWRGD.curr_state_RNI7N705Z0Z_0\,
            ltout => \PCH_PWRGD.curr_state_RNI7N705Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_RNO_0_15_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__20060\,
            in1 => \_gnd_net_\,
            in2 => \N__8930\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.N_65_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_RNIFR521_15_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9814\,
            in1 => \N__9829\,
            in2 => \N__9797\,
            in3 => \N__9595\,
            lcout => \PCH_PWRGD.un4_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_sys_pwrok_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__19283\,
            in1 => \N__8918\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.N_3_i\,
            ltout => \PCH_PWRGD.N_3_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_0_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__8898\,
            in1 => \N__8878\,
            in2 => \N__8921\,
            in3 => \N__8845\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20560\,
            ce => \N__19787\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.pch_pwrok_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8900\,
            in1 => \N__8844\,
            in2 => \_gnd_net_\,
            in3 => \N__8865\,
            lcout => pch_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20560\,
            ce => \N__19787\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIHKNI1_0_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__8842\,
            in1 => \N__8897\,
            in2 => \N__19286\,
            in3 => \N__8917\,
            lcout => \PCH_PWRGD.un1_curr_state10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_1_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101010000"
        )
    port map (
            in0 => \N__8899\,
            in1 => \N__8879\,
            in2 => \N__8870\,
            in3 => \N__8843\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20560\,
            ce => \N__19787\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12848\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_5_0_\,
            carryout => \POWERLED.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11663\,
            in2 => \N__9889\,
            in3 => \N__8825\,
            lcout => \POWERLED.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_2\,
            carryout => \POWERLED.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9885\,
            in2 => \N__9752\,
            in3 => \N__8963\,
            lcout => \POWERLED.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_3\,
            carryout => \POWERLED.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9740\,
            in2 => \N__10102\,
            in3 => \N__8960\,
            lcout => \POWERLED.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_4\,
            carryout => \POWERLED.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10098\,
            in2 => \N__9731\,
            in3 => \N__8957\,
            lcout => \POWERLED.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_5\,
            carryout => \POWERLED.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10121\,
            in1 => \N__9719\,
            in2 => \N__9890\,
            in3 => \N__8954\,
            lcout => \POWERLED.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_6\,
            carryout => \POWERLED.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9905\,
            in2 => \_gnd_net_\,
            in3 => \N__8951\,
            lcout => \POWERLED.mult1_un89_sum_s_8\,
            ltout => \POWERLED.mult1_un89_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8948\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12874\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \POWERLED.mult1_un96_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10295\,
            in2 => \N__9019\,
            in3 => \N__8945\,
            lcout => \POWERLED.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_2\,
            carryout => \POWERLED.mult1_un96_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9015\,
            in2 => \N__8942\,
            in3 => \N__8933\,
            lcout => \POWERLED.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_3\,
            carryout => \POWERLED.mult1_un96_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9047\,
            in2 => \N__10129\,
            in3 => \N__9041\,
            lcout => \POWERLED.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_4\,
            carryout => \POWERLED.mult1_un96_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10125\,
            in2 => \N__9038\,
            in3 => \N__9029\,
            lcout => \POWERLED.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_5\,
            carryout => \POWERLED.mult1_un96_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9560\,
            in1 => \N__9026\,
            in2 => \N__9020\,
            in3 => \N__9002\,
            lcout => \POWERLED.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_6\,
            carryout => \POWERLED.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8999\,
            in2 => \_gnd_net_\,
            in3 => \N__8993\,
            lcout => \POWERLED.mult1_un96_sum_s_8\,
            ltout => \POWERLED.mult1_un96_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8990\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12916\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => \POWERLED.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9581\,
            in2 => \N__9103\,
            in3 => \N__8987\,
            lcout => \POWERLED.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_2\,
            carryout => \POWERLED.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9099\,
            in2 => \N__8984\,
            in3 => \N__8975\,
            lcout => \POWERLED.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_3\,
            carryout => \POWERLED.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8972\,
            in2 => \N__9568\,
            in3 => \N__8966\,
            lcout => \POWERLED.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_4\,
            carryout => \POWERLED.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9564\,
            in2 => \N__9122\,
            in3 => \N__9113\,
            lcout => \POWERLED.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_5\,
            carryout => \POWERLED.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10007\,
            in1 => \N__9110\,
            in2 => \N__9104\,
            in3 => \N__9086\,
            lcout => \POWERLED.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_6\,
            carryout => \POWERLED.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9083\,
            in2 => \_gnd_net_\,
            in3 => \N__9077\,
            lcout => \POWERLED.mult1_un103_sum_s_8\,
            ltout => \POWERLED.mult1_un103_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9074\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12950\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_8_0_\,
            carryout => \POWERLED.mult1_un110_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10019\,
            in2 => \N__9166\,
            in3 => \N__9071\,
            lcout => \POWERLED.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_2\,
            carryout => \POWERLED.mult1_un110_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9162\,
            in2 => \N__9068\,
            in3 => \N__9059\,
            lcout => \POWERLED.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_3\,
            carryout => \POWERLED.mult1_un110_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9056\,
            in2 => \N__10013\,
            in3 => \N__9050\,
            lcout => \POWERLED.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_4\,
            carryout => \POWERLED.mult1_un110_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10011\,
            in2 => \N__9185\,
            in3 => \N__9176\,
            lcout => \POWERLED.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_5\,
            carryout => \POWERLED.mult1_un110_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10229\,
            in1 => \N__9173\,
            in2 => \N__9167\,
            in3 => \N__9149\,
            lcout => \POWERLED.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_6\,
            carryout => \POWERLED.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9146\,
            in2 => \_gnd_net_\,
            in3 => \N__9140\,
            lcout => \POWERLED.mult1_un110_sum_s_8\,
            ltout => \POWERLED.mult1_un110_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9137\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13007\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \POWERLED.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11369\,
            in2 => \N__10396\,
            in3 => \N__9134\,
            lcout => \POWERLED.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_2\,
            carryout => \POWERLED.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10392\,
            in2 => \N__10283\,
            in3 => \N__9131\,
            lcout => \POWERLED.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_3\,
            carryout => \POWERLED.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10262\,
            in2 => \N__10321\,
            in3 => \N__9128\,
            lcout => \POWERLED.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_4\,
            carryout => \POWERLED.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10317\,
            in2 => \N__10247\,
            in3 => \N__9125\,
            lcout => \POWERLED.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_5\,
            carryout => \POWERLED.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10373\,
            in1 => \N__10202\,
            in2 => \N__10397\,
            in3 => \N__9257\,
            lcout => \POWERLED.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_6\,
            carryout => \POWERLED.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10169\,
            in2 => \_gnd_net_\,
            in3 => \N__9254\,
            lcout => \POWERLED.mult1_un124_sum_s_8\,
            ltout => \POWERLED.mult1_un124_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9251\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12682\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \POWERLED.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11381\,
            in2 => \N__9205\,
            in3 => \N__9248\,
            lcout => \POWERLED.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_2\,
            carryout => \POWERLED.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9201\,
            in2 => \N__9245\,
            in3 => \N__9236\,
            lcout => \POWERLED.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_3\,
            carryout => \POWERLED.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9233\,
            in2 => \N__10379\,
            in3 => \N__9227\,
            lcout => \POWERLED.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_4\,
            carryout => \POWERLED.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10377\,
            in2 => \N__9224\,
            in3 => \N__9215\,
            lcout => \POWERLED.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_5\,
            carryout => \POWERLED.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10349\,
            in1 => \N__9212\,
            in2 => \N__9206\,
            in3 => \N__9188\,
            lcout => \POWERLED.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_6\,
            carryout => \POWERLED.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9338\,
            in2 => \_gnd_net_\,
            in3 => \N__9332\,
            lcout => \POWERLED.mult1_un131_sum_s_8\,
            ltout => \POWERLED.mult1_un131_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9329\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12730\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \POWERLED.mult1_un138_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10331\,
            in2 => \N__9283\,
            in3 => \N__9326\,
            lcout => \POWERLED.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_2\,
            carryout => \POWERLED.mult1_un138_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9279\,
            in2 => \N__9323\,
            in3 => \N__9314\,
            lcout => \POWERLED.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_3\,
            carryout => \POWERLED.mult1_un138_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9311\,
            in2 => \N__10355\,
            in3 => \N__9305\,
            lcout => \POWERLED.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_4\,
            carryout => \POWERLED.mult1_un138_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10353\,
            in2 => \N__9302\,
            in3 => \N__9293\,
            lcout => \POWERLED.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_5\,
            carryout => \POWERLED.mult1_un138_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11326\,
            in1 => \N__9290\,
            in2 => \N__9284\,
            in3 => \N__9266\,
            lcout => \POWERLED.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_6\,
            carryout => \POWERLED.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9263\,
            in2 => \_gnd_net_\,
            in3 => \N__9365\,
            lcout => \POWERLED.mult1_un138_sum_s_8\,
            ltout => \POWERLED.mult1_un138_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9362\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14129\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \POWERLED.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11540\,
            in2 => \N__10516\,
            in3 => \N__9359\,
            lcout => \POWERLED.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_1\,
            carryout => \POWERLED.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10512\,
            in2 => \N__10676\,
            in3 => \N__9356\,
            lcout => \POWERLED.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_2\,
            carryout => \POWERLED.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10655\,
            in2 => \N__10544\,
            in3 => \N__9353\,
            lcout => \POWERLED.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_3\,
            carryout => \POWERLED.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10542\,
            in2 => \N__10640\,
            in3 => \N__9350\,
            lcout => \POWERLED.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_4\,
            carryout => \POWERLED.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9418\,
            in1 => \N__10595\,
            in2 => \N__10517\,
            in3 => \N__9347\,
            lcout => \POWERLED.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_5\,
            carryout => \POWERLED.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10562\,
            in2 => \_gnd_net_\,
            in3 => \N__9344\,
            lcout => \POWERLED.mult1_un159_sum_s_7\,
            ltout => \POWERLED.mult1_un159_sum_s_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9341\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14209\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \POWERLED.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11552\,
            in2 => \N__9391\,
            in3 => \N__9413\,
            lcout => \G_407\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_0\,
            carryout => \POWERLED.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9387\,
            in2 => \N__9443\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_1\,
            carryout => \POWERLED.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9414\,
            in2 => \N__9434\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_2\,
            carryout => \POWERLED.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9425\,
            in2 => \N__9419\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_3\,
            carryout => \POWERLED.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9398\,
            in2 => \N__9392\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_4\,
            carryout => \POWERLED.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9374\,
            in2 => \_gnd_net_\,
            in3 => \N__9368\,
            lcout => \POWERLED.un1_count_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10543\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12878\,
            lcout => \POWERLED.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9572\,
            lcout => \POWERLED.un1_count_2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11602\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => pwrbtn_led,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20628\,
            ce => \N__11087\,
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_0_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__11601\,
            in1 => \N__11612\,
            in2 => \_gnd_net_\,
            in3 => \N__10823\,
            lcout => \POWERLED.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20629\,
            ce => \N__19812\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20074\,
            in1 => \N__9515\,
            in2 => \N__9533\,
            in3 => \N__9532\,
            lcout => \PCH_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_2_0_\,
            carryout => \PCH_PWRGD.un1_count_1_cry_0\,
            clk => \N__20466\,
            ce => 'H',
            sr => \N__9769\
        );

    \PCH_PWRGD.count_1_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20067\,
            in1 => \N__9503\,
            in2 => \_gnd_net_\,
            in3 => \N__9491\,
            lcout => \PCH_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_0\,
            carryout => \PCH_PWRGD.un1_count_1_cry_1\,
            clk => \N__20466\,
            ce => 'H',
            sr => \N__9769\
        );

    \PCH_PWRGD.count_2_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20075\,
            in1 => \N__9488\,
            in2 => \_gnd_net_\,
            in3 => \N__9476\,
            lcout => \PCH_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_1\,
            carryout => \PCH_PWRGD.un1_count_1_cry_2\,
            clk => \N__20466\,
            ce => 'H',
            sr => \N__9769\
        );

    \PCH_PWRGD.count_3_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20068\,
            in1 => \N__9473\,
            in2 => \_gnd_net_\,
            in3 => \N__9461\,
            lcout => \PCH_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_2\,
            carryout => \PCH_PWRGD.un1_count_1_cry_3\,
            clk => \N__20466\,
            ce => 'H',
            sr => \N__9769\
        );

    \PCH_PWRGD.count_4_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20076\,
            in1 => \N__9458\,
            in2 => \_gnd_net_\,
            in3 => \N__9446\,
            lcout => \PCH_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_3\,
            carryout => \PCH_PWRGD.un1_count_1_cry_4\,
            clk => \N__20466\,
            ce => 'H',
            sr => \N__9769\
        );

    \PCH_PWRGD.count_5_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20069\,
            in1 => \N__9710\,
            in2 => \_gnd_net_\,
            in3 => \N__9698\,
            lcout => \PCH_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_4\,
            carryout => \PCH_PWRGD.un1_count_1_cry_5\,
            clk => \N__20466\,
            ce => 'H',
            sr => \N__9769\
        );

    \PCH_PWRGD.count_6_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20077\,
            in1 => \N__9695\,
            in2 => \_gnd_net_\,
            in3 => \N__9683\,
            lcout => \PCH_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_5\,
            carryout => \PCH_PWRGD.un1_count_1_cry_6\,
            clk => \N__20466\,
            ce => 'H',
            sr => \N__9769\
        );

    \PCH_PWRGD.count_7_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20070\,
            in1 => \N__9679\,
            in2 => \_gnd_net_\,
            in3 => \N__9665\,
            lcout => \PCH_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_6\,
            carryout => \PCH_PWRGD.un1_count_1_cry_7\,
            clk => \N__20466\,
            ce => 'H',
            sr => \N__9769\
        );

    \PCH_PWRGD.count_8_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20117\,
            in1 => \N__9662\,
            in2 => \_gnd_net_\,
            in3 => \N__9650\,
            lcout => \PCH_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_3_0_\,
            carryout => \PCH_PWRGD.un1_count_1_cry_8\,
            clk => \N__20532\,
            ce => 'H',
            sr => \N__9768\
        );

    \PCH_PWRGD.count_9_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20102\,
            in1 => \N__9647\,
            in2 => \_gnd_net_\,
            in3 => \N__9635\,
            lcout => \PCH_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_8\,
            carryout => \PCH_PWRGD.un1_count_1_cry_9\,
            clk => \N__20532\,
            ce => 'H',
            sr => \N__9768\
        );

    \PCH_PWRGD.count_10_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20114\,
            in1 => \N__9631\,
            in2 => \_gnd_net_\,
            in3 => \N__9617\,
            lcout => \PCH_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_9\,
            carryout => \PCH_PWRGD.un1_count_1_cry_10\,
            clk => \N__20532\,
            ce => 'H',
            sr => \N__9768\
        );

    \PCH_PWRGD.count_11_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20100\,
            in1 => \N__9613\,
            in2 => \_gnd_net_\,
            in3 => \N__9599\,
            lcout => \PCH_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_10\,
            carryout => \PCH_PWRGD.un1_count_1_cry_11\,
            clk => \N__20532\,
            ce => 'H',
            sr => \N__9768\
        );

    \PCH_PWRGD.count_12_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20115\,
            in1 => \N__9596\,
            in2 => \_gnd_net_\,
            in3 => \N__9584\,
            lcout => \PCH_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_11\,
            carryout => \PCH_PWRGD.un1_count_1_cry_12\,
            clk => \N__20532\,
            ce => 'H',
            sr => \N__9768\
        );

    \PCH_PWRGD.count_13_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20101\,
            in1 => \N__9830\,
            in2 => \_gnd_net_\,
            in3 => \N__9818\,
            lcout => \PCH_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_12\,
            carryout => \PCH_PWRGD.un1_count_1_cry_13\,
            clk => \N__20532\,
            ce => 'H',
            sr => \N__9768\
        );

    \PCH_PWRGD.count_14_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20116\,
            in1 => \N__9815\,
            in2 => \_gnd_net_\,
            in3 => \N__9803\,
            lcout => \PCH_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_13\,
            carryout => \PCH_PWRGD.un1_count_1_cry_14\,
            clk => \N__20532\,
            ce => 'H',
            sr => \N__9768\
        );

    \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18395\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_14\,
            carryout => \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_15_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9796\,
            in2 => \_gnd_net_\,
            in3 => \N__9800\,
            lcout => \PCH_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20542\,
            ce => \N__9782\,
            sr => \N__9770\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12818\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_5_0_\,
            carryout => \POWERLED.mult1_un82_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11753\,
            in2 => \N__9973\,
            in3 => \N__9743\,
            lcout => \POWERLED.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_2\,
            carryout => \POWERLED.mult1_un82_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9969\,
            in2 => \N__9872\,
            in3 => \N__9734\,
            lcout => \POWERLED.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_3\,
            carryout => \POWERLED.mult1_un82_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9860\,
            in2 => \N__10045\,
            in3 => \N__9722\,
            lcout => \POWERLED.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_4\,
            carryout => \POWERLED.mult1_un82_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10041\,
            in2 => \N__9851\,
            in3 => \N__9713\,
            lcout => \POWERLED.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_5\,
            carryout => \POWERLED.mult1_un82_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10094\,
            in1 => \N__9839\,
            in2 => \N__9974\,
            in3 => \N__9899\,
            lcout => \POWERLED.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_6\,
            carryout => \POWERLED.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9989\,
            in2 => \_gnd_net_\,
            in3 => \N__9896\,
            lcout => \POWERLED.mult1_un82_sum_s_8\,
            ltout => \POWERLED.mult1_un82_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9893\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12794\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_6_0_\,
            carryout => \POWERLED.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11285\,
            in2 => \N__10147\,
            in3 => \N__9863\,
            lcout => \POWERLED.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_2\,
            carryout => \POWERLED.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10143\,
            in2 => \N__9956\,
            in3 => \N__9854\,
            lcout => \POWERLED.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_3\,
            carryout => \POWERLED.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9944\,
            in2 => \N__10076\,
            in3 => \N__9842\,
            lcout => \POWERLED.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_4\,
            carryout => \POWERLED.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10074\,
            in2 => \N__9935\,
            in3 => \N__9833\,
            lcout => \POWERLED.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_5\,
            carryout => \POWERLED.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10037\,
            in1 => \N__9923\,
            in2 => \N__10148\,
            in3 => \N__9983\,
            lcout => \POWERLED.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_6\,
            carryout => \POWERLED.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9914\,
            in2 => \_gnd_net_\,
            in3 => \N__9980\,
            lcout => \POWERLED.mult1_un75_sum_s_8\,
            ltout => \POWERLED.mult1_un75_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9977\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13184\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => \POWERLED.mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11768\,
            in2 => \N__11428\,
            in3 => \N__9947\,
            lcout => \POWERLED.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_2\,
            carryout => \POWERLED.mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11424\,
            in2 => \N__11276\,
            in3 => \N__9938\,
            lcout => \POWERLED.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_3\,
            carryout => \POWERLED.mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11246\,
            in2 => \N__11464\,
            in3 => \N__9926\,
            lcout => \POWERLED.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_4\,
            carryout => \POWERLED.mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11460\,
            in2 => \N__11225\,
            in3 => \N__9917\,
            lcout => \POWERLED.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_5\,
            carryout => \POWERLED.mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10070\,
            in1 => \N__11198\,
            in2 => \N__11429\,
            in3 => \N__9908\,
            lcout => \POWERLED.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_6\,
            carryout => \POWERLED.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11159\,
            in2 => \_gnd_net_\,
            in3 => \N__10151\,
            lcout => \POWERLED.mult1_un68_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10069\,
            lcout => \POWERLED.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10234\,
            lcout => \POWERLED.un1_count_2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10130\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10103\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10075\,
            lcout => \POWERLED.un1_count_2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10046\,
            lcout => \POWERLED.un1_count_2_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12917\,
            lcout => \POWERLED.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10012\,
            lcout => \POWERLED.un1_count_2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12847\,
            lcout => \POWERLED.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12979\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => \POWERLED.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11408\,
            in2 => \N__10186\,
            in3 => \N__10274\,
            lcout => \POWERLED.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_2\,
            carryout => \POWERLED.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10182\,
            in2 => \N__10271\,
            in3 => \N__10256\,
            lcout => \POWERLED.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_3\,
            carryout => \POWERLED.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10253\,
            in2 => \N__10235\,
            in3 => \N__10238\,
            lcout => \POWERLED.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_4\,
            carryout => \POWERLED.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10233\,
            in2 => \N__10211\,
            in3 => \N__10196\,
            lcout => \POWERLED.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_5\,
            carryout => \POWERLED.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10313\,
            in1 => \N__10193\,
            in2 => \N__10187\,
            in3 => \N__10163\,
            lcout => \POWERLED.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_6\,
            carryout => \POWERLED.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10160\,
            in2 => \_gnd_net_\,
            in3 => \N__10154\,
            lcout => \POWERLED.mult1_un117_sum_s_8\,
            ltout => \POWERLED.mult1_un117_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10400\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10378\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10354\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_4_l_fx_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__10472\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11325\,
            lcout => \POWERLED.mult1_un145_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10627\,
            lcout => \POWERLED.un1_count_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12683\,
            lcout => \POWERLED.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12758\,
            lcout => \POWERLED.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10322\,
            lcout => \POWERLED.un1_count_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11465\,
            lcout => \POWERLED.un1_count_2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12757\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \POWERLED.mult1_un145_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11396\,
            in2 => \N__10484\,
            in3 => \N__10475\,
            lcout => \POWERLED.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_2\,
            carryout => \POWERLED.mult1_un145_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10471\,
            in2 => \N__10460\,
            in3 => \N__10451\,
            lcout => \POWERLED.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_3\,
            carryout => \POWERLED.mult1_un145_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10448\,
            in2 => \N__11333\,
            in3 => \N__10439\,
            lcout => \POWERLED.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_4\,
            carryout => \POWERLED.mult1_un145_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11330\,
            in2 => \N__10436\,
            in3 => \N__10427\,
            lcout => \POWERLED.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_5\,
            carryout => \POWERLED.mult1_un145_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10622\,
            in1 => \N__11356\,
            in2 => \N__11345\,
            in3 => \N__10424\,
            lcout => \POWERLED.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_6\,
            carryout => \POWERLED.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10421\,
            in2 => \_gnd_net_\,
            in3 => \N__10415\,
            lcout => \POWERLED.mult1_un145_sum_s_8\,
            ltout => \POWERLED.mult1_un145_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10412\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14752\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \POWERLED.mult1_un152_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10409\,
            in2 => \N__10579\,
            in3 => \N__10667\,
            lcout => \POWERLED.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_2\,
            carryout => \POWERLED.mult1_un152_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10575\,
            in2 => \N__10664\,
            in3 => \N__10649\,
            lcout => \POWERLED.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_3\,
            carryout => \POWERLED.mult1_un152_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10646\,
            in2 => \N__10628\,
            in3 => \N__10631\,
            lcout => \POWERLED.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_4\,
            carryout => \POWERLED.mult1_un152_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10626\,
            in2 => \N__10604\,
            in3 => \N__10589\,
            lcout => \POWERLED.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_5\,
            carryout => \POWERLED.mult1_un152_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10538\,
            in1 => \N__10586\,
            in2 => \N__10580\,
            in3 => \N__10556\,
            lcout => \POWERLED.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_6\,
            carryout => \POWERLED.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10553\,
            in2 => \_gnd_net_\,
            in3 => \N__10547\,
            lcout => \POWERLED.mult1_un152_sum_s_8\,
            ltout => \POWERLED.mult1_un152_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10520\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_0_c_inv_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10490\,
            in2 => \N__10499\,
            in3 => \N__12041\,
            lcout => \POWERLED.count_i_0_0\,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \POWERLED.un1_count_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_1_c_inv_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10808\,
            in2 => \N__10817\,
            in3 => \N__12017\,
            lcout => \POWERLED.count_i_1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_0\,
            carryout => \POWERLED.un1_count_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_2_c_inv_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11990\,
            in1 => \N__10799\,
            in2 => \N__10793\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_i_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_1\,
            carryout => \POWERLED.un1_count_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_3_c_inv_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10784\,
            in2 => \N__10775\,
            in3 => \N__11960\,
            lcout => \POWERLED.count_i_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_2\,
            carryout => \POWERLED.un1_count_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_4_c_inv_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11297\,
            in2 => \N__10766\,
            in3 => \N__12476\,
            lcout => \POWERLED.count_i_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_3\,
            carryout => \POWERLED.un1_count_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_5_c_inv_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10754\,
            in2 => \N__10745\,
            in3 => \N__12446\,
            lcout => \POWERLED.count_i_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_4\,
            carryout => \POWERLED.un1_count_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_6_c_inv_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10736\,
            in2 => \N__10727\,
            in3 => \N__12416\,
            lcout => \POWERLED.count_i_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_5\,
            carryout => \POWERLED.un1_count_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_7_c_inv_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10715\,
            in2 => \N__10706\,
            in3 => \N__12385\,
            lcout => \POWERLED.count_i_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_6\,
            carryout => \POWERLED.un1_count_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_8_c_inv_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10694\,
            in2 => \N__10685\,
            in3 => \N__12353\,
            lcout => \POWERLED.count_i_8\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \POWERLED.un1_count_2_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_9_c_inv_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10967\,
            in2 => \N__10958\,
            in3 => \N__12326\,
            lcout => \POWERLED.count_i_9\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_8\,
            carryout => \POWERLED.un1_count_2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_10_c_inv_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12290\,
            in1 => \N__10949\,
            in2 => \N__10943\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_i_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_9\,
            carryout => \POWERLED.un1_count_2_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_11_c_inv_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10934\,
            in2 => \N__10925\,
            in3 => \N__12260\,
            lcout => \POWERLED.count_i_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_10\,
            carryout => \POWERLED.un1_count_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_12_c_inv_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10916\,
            in2 => \N__10904\,
            in3 => \N__12227\,
            lcout => \POWERLED.count_i_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_11\,
            carryout => \POWERLED.un1_count_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_13_c_inv_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10892\,
            in2 => \N__10880\,
            in3 => \N__12626\,
            lcout => \POWERLED.count_i_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_12\,
            carryout => \POWERLED.un1_count_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_14_c_inv_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10871\,
            in2 => \N__10859\,
            in3 => \N__12596\,
            lcout => \POWERLED.count_i_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_13\,
            carryout => \POWERLED.un1_count_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_15_c_inv_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10847\,
            in2 => \N__10835\,
            in3 => \N__12560\,
            lcout => \POWERLED.count_i_15\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_14\,
            carryout => \POWERLED.un1_count_2_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10826\,
            lcout => \POWERLED.un1_count_2_cry_15_THRU_CO\,
            ltout => \POWERLED.un1_count_2_cry_15_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__11600\,
            in1 => \N__11525\,
            in2 => \N__11090\,
            in3 => \N__17738\,
            lcout => \POWERLED.pwm_out_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_vddq_en_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11075\,
            in2 => \_gnd_net_\,
            in3 => \N__15659\,
            lcout => vddq_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNI1S0J_0_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11021\,
            in2 => \_gnd_net_\,
            in3 => \N__15777\,
            lcout => \HDA_STRAP.N_5_0\,
            ltout => \HDA_STRAP.N_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_0_0_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101010101"
        )
    port map (
            in0 => \N__15778\,
            in1 => \N__11051\,
            in2 => \N__11036\,
            in3 => \N__15867\,
            lcout => \HDA_STRAP.m14_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_0_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010100011"
        )
    port map (
            in0 => \N__11029\,
            in1 => \N__15735\,
            in2 => \N__10985\,
            in3 => \N__15914\,
            lcout => \HDA_STRAP.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20428\,
            ce => \N__19740\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13139\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_5_0_\,
            carryout => \POWERLED.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11654\,
            in3 => \N__10976\,
            lcout => \POWERLED.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_2\,
            carryout => \POWERLED.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11138\,
            in3 => \N__10973\,
            lcout => \POWERLED.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_3\,
            carryout => \POWERLED.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18387\,
            in2 => \N__11126\,
            in3 => \N__10970\,
            lcout => \POWERLED.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_4\,
            carryout => \POWERLED.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18388\,
            in2 => \N__11114\,
            in3 => \N__11147\,
            lcout => \POWERLED.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_5\,
            carryout => \POWERLED.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11512\,
            in2 => \_gnd_net_\,
            in3 => \N__11144\,
            lcout => \POWERLED.mult1_un54_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_6\,
            carryout => \POWERLED.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11141\,
            lcout => \POWERLED.mult1_un54_sum_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13118\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_6_0_\,
            carryout => \POWERLED.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11777\,
            in3 => \N__11129\,
            lcout => \POWERLED.mult1_un47_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_2\,
            carryout => \POWERLED.mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11711\,
            in3 => \N__11117\,
            lcout => \POWERLED.mult1_un47_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_3\,
            carryout => \POWERLED.mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18376\,
            in2 => \N__11729\,
            in3 => \N__11105\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_4\,
            carryout => \POWERLED.mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18377\,
            in2 => \N__11720\,
            in3 => \N__11102\,
            lcout => \POWERLED.mult1_un47_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_5\,
            carryout => \POWERLED.mult1_un47_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11099\,
            in2 => \_gnd_net_\,
            in3 => \N__11093\,
            lcout => \POWERLED.mult1_un54_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13183\,
            lcout => \POWERLED.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11495\,
            lcout => \POWERLED.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13160\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_7_0_\,
            carryout => \POWERLED.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11759\,
            in2 => \N__11176\,
            in3 => \N__11264\,
            lcout => \POWERLED.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_2\,
            carryout => \POWERLED.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11172\,
            in2 => \N__11261\,
            in3 => \N__11237\,
            lcout => \POWERLED.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_3\,
            carryout => \POWERLED.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11234\,
            in2 => \N__11501\,
            in3 => \N__11213\,
            lcout => \POWERLED.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_4\,
            carryout => \POWERLED.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11499\,
            in2 => \N__11210\,
            in3 => \N__11189\,
            lcout => \POWERLED.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_5\,
            carryout => \POWERLED.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11448\,
            in1 => \N__11186\,
            in2 => \N__11177\,
            in3 => \N__11150\,
            lcout => \POWERLED.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_6\,
            carryout => \POWERLED.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11513\,
            in1 => \N__11500\,
            in2 => \N__11480\,
            in3 => \N__11468\,
            lcout => \POWERLED.mult1_un61_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11447\,
            lcout => \POWERLED.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12949\,
            lcout => \POWERLED.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12731\,
            lcout => \POWERLED.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13006\,
            lcout => \POWERLED.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12983\,
            lcout => \POWERLED.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIV4PD6_1_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__13706\,
            in1 => \N__15302\,
            in2 => \_gnd_net_\,
            in3 => \N__13529\,
            lcout => \POWERLED.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_7_l_fx_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__11360\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11331\,
            lcout => \POWERLED.mult1_un145_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11332\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_EN_i_i_i_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15019\,
            lcout => v5s_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14127\,
            lcout => \POWERLED.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14753\,
            lcout => \POWERLED.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_1_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__12015\,
            in1 => \N__12040\,
            in2 => \_gnd_net_\,
            in3 => \N__20123\,
            lcout => \POWERLED.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20615\,
            ce => 'H',
            sr => \N__12524\
        );

    \POWERLED.count_0_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12039\,
            in2 => \_gnd_net_\,
            in3 => \N__20122\,
            lcout => \POWERLED.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20615\,
            ce => 'H',
            sr => \N__12524\
        );

    \POWERLED.pwm_out_RNO_4_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12468\,
            in1 => \N__11952\,
            in2 => \_gnd_net_\,
            in3 => \N__11982\,
            lcout => OPEN,
            ltout => \POWERLED.un1_countlt6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_2_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__12441\,
            in1 => \N__11627\,
            in2 => \N__11531\,
            in3 => \N__12411\,
            lcout => OPEN,
            ltout => \POWERLED.g0_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_0_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__12282\,
            in1 => \N__12384\,
            in2 => \N__11528\,
            in3 => \N__11639\,
            lcout => \POWERLED.un1_count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNID4E61_7_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12320\,
            in1 => \N__12347\,
            in2 => \N__12386\,
            in3 => \N__12281\,
            lcout => OPEN,
            ltout => \POWERLED.un1_countlto15_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI6IPJ2_5_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001110000"
        )
    port map (
            in0 => \N__12410\,
            in1 => \N__12440\,
            in2 => \N__11642\,
            in3 => \N__11633\,
            lcout => \POWERLED.un1_countlto15_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_1_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12222\,
            in1 => \N__12254\,
            in2 => \_gnd_net_\,
            in3 => \N__12348\,
            lcout => \POWERLED.g0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNICO6R_2_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12467\,
            in1 => \N__11951\,
            in2 => \_gnd_net_\,
            in3 => \N__11981\,
            lcout => \POWERLED.un1_countlt6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_3_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12621\,
            in1 => \N__12591\,
            in2 => \N__12325\,
            in3 => \N__12551\,
            lcout => \POWERLED.g0_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_esr_RNIBHMO_15_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12552\,
            in1 => \N__12590\,
            in2 => \_gnd_net_\,
            in3 => \N__12620\,
            lcout => OPEN,
            ltout => \POWERLED.un1_countlto15_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIOVT24_11_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__12221\,
            in1 => \N__12255\,
            in2 => \N__11621\,
            in3 => \N__11618\,
            lcout => \POWERLED.count_RNIOVT24Z0Z_11\,
            ltout => \POWERLED.count_RNIOVT24Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNI75RB5_0_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11603\,
            in2 => \N__11576\,
            in3 => \N__20063\,
            lcout => \POWERLED.curr_state_RNI75RB5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_esr_RNO_0_15_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__12514\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20066\,
            lcout => \POWERLED.N_65_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_0_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__15807\,
            in1 => \N__15737\,
            in2 => \N__15901\,
            in3 => \N__12488\,
            lcout => \HDA_STRAP.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20443\,
            ce => \N__19784\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_1_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100011111000"
        )
    port map (
            in0 => \N__15736\,
            in1 => \N__15808\,
            in2 => \N__15900\,
            in3 => \N__11702\,
            lcout => \HDA_STRAP.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20443\,
            ce => \N__19784\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_11_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__15787\,
            in1 => \N__15734\,
            in2 => \N__15899\,
            in3 => \N__12635\,
            lcout => \HDA_STRAP.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20467\,
            ce => \N__19763\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_2_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000001100"
        )
    port map (
            in0 => \N__11701\,
            in1 => \N__11689\,
            in2 => \N__14036\,
            in3 => \N__15872\,
            lcout => \HDA_STRAP.curr_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20467\,
            ce => \N__19763\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.HDA_SDO_FPGA_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__15788\,
            in1 => \N__15868\,
            in2 => \_gnd_net_\,
            in3 => \N__11690\,
            lcout => hda_sdo_atp,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20467\,
            ce => \N__19763\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIFHLJ_0_0_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14604\,
            in2 => \N__14110\,
            in3 => \N__14177\,
            lcout => \POWERLED.un1_dutycycle_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI16B71_5_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__12697\,
            in1 => \N__14530\,
            in2 => \N__14751\,
            in3 => \N__14088\,
            lcout => \POWERLED.dutycycle_RNI16B71Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12811\,
            lcout => \POWERLED.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13114\,
            lcout => \POWERLED.un1_dutycycle_1_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNIMOAE_5_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16081\,
            in2 => \_gnd_net_\,
            in3 => \N__13041\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_1_19_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIEJ021_4_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__14605\,
            in1 => \N__14398\,
            in2 => \N__11645\,
            in3 => \N__14666\,
            lcout => \POWERLED.dutycycle_RNIEJ021Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12793\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIFHLJ_0_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14606\,
            in2 => \N__14111\,
            in3 => \N__14178\,
            lcout => \POWERLED.dutycycle_RNIFHLJZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16769\,
            in1 => \N__11744\,
            in2 => \_gnd_net_\,
            in3 => \N__14051\,
            lcout => \POWERLED.dutycycleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20471\,
            ce => \N__19773\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_0_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11743\,
            in1 => \N__16770\,
            in2 => \_gnd_net_\,
            in3 => \N__14144\,
            lcout => \POWERLED.dutycycleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20471\,
            ce => \N__19773\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNIVCSK_5_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14736\,
            in2 => \N__14112\,
            in3 => \N__13042\,
            lcout => \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_5_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__13430\,
            in1 => \N__16771\,
            in2 => \N__13593\,
            in3 => \N__14486\,
            lcout => \POWERLED.dutycycle_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20471\,
            ce => \N__19773\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13069\,
            in2 => \N__13097\,
            in3 => \N__13051\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__13052\,
            in1 => \_gnd_net_\,
            in2 => \N__13073\,
            in3 => \N__13095\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13096\,
            in3 => \N__13068\,
            lcout => \POWERLED.mult1_un47_sum_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13088\,
            lcout => \POWERLED.un1_dutycycle_1_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13156\,
            lcout => \POWERLED.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13135\,
            lcout => \POWERLED.mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI4I7Q_0_5_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__14123\,
            in1 => \N__14196\,
            in2 => \N__14532\,
            in3 => \N__14444\,
            lcout => \POWERLED.N_234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_5_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__16773\,
            in1 => \N__13421\,
            in2 => \N__13594\,
            in3 => \N__14485\,
            lcout => \POWERLED.dutycycleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20564\,
            ce => \N__19798\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6NI81_5_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__13021\,
            in1 => \N__16242\,
            in2 => \N__14531\,
            in3 => \N__14443\,
            lcout => \POWERLED.dutycycle_RNI6NI81Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_6_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__16774\,
            in1 => \N__13422\,
            in2 => \N__13595\,
            in3 => \N__14416\,
            lcout => \POWERLED.dutycycleZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20564\,
            ce => \N__19798\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_6_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101010"
        )
    port map (
            in0 => \N__14417\,
            in1 => \N__13586\,
            in2 => \N__13429\,
            in3 => \N__16775\,
            lcout => \POWERLED.dutycycle_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20564\,
            ce => \N__19798\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJNBA1_6_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__13198\,
            in1 => \N__14442\,
            in2 => \N__16292\,
            in3 => \N__14385\,
            lcout => \POWERLED.dutycycle_RNIJNBA1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNILMLM_6_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16288\,
            in2 => \N__14397\,
            in3 => \N__13218\,
            lcout => \POWERLED.dutycycle_fast_RNILMLMZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_0_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12062\,
            in1 => \N__11842\,
            in2 => \N__13457\,
            in3 => \N__13456\,
            lcout => \POWERLED.count_offZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \POWERLED.un1_count_off_1_cry_0\,
            clk => \N__20585\,
            ce => \N__19797\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_1_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12116\,
            in1 => \N__11869\,
            in2 => \_gnd_net_\,
            in3 => \N__11801\,
            lcout => \POWERLED.count_offZ0Z_1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_0\,
            carryout => \POWERLED.un1_count_off_1_cry_1\,
            clk => \N__20585\,
            ce => \N__19797\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_2_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12063\,
            in1 => \N__13325\,
            in2 => \_gnd_net_\,
            in3 => \N__11798\,
            lcout => \POWERLED.count_offZ0Z_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_1\,
            carryout => \POWERLED.un1_count_off_1_cry_2\,
            clk => \N__20585\,
            ce => \N__19797\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_3_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12117\,
            in1 => \N__13367\,
            in2 => \_gnd_net_\,
            in3 => \N__11795\,
            lcout => \POWERLED.count_offZ0Z_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_2\,
            carryout => \POWERLED.un1_count_off_1_cry_3\,
            clk => \N__20585\,
            ce => \N__19797\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_4_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12119\,
            in1 => \N__13339\,
            in2 => \_gnd_net_\,
            in3 => \N__11792\,
            lcout => \POWERLED.count_offZ0Z_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_3\,
            carryout => \POWERLED.un1_count_off_1_cry_4\,
            clk => \N__20585\,
            ce => \N__19797\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_5_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12065\,
            in1 => \N__12148\,
            in2 => \_gnd_net_\,
            in3 => \N__11789\,
            lcout => \POWERLED.count_offZ0Z_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_4\,
            carryout => \POWERLED.un1_count_off_1_cry_5\,
            clk => \N__20585\,
            ce => \N__19797\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_6_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12064\,
            in1 => \N__12178\,
            in2 => \_gnd_net_\,
            in3 => \N__11786\,
            lcout => \POWERLED.count_offZ0Z_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_5\,
            carryout => \POWERLED.un1_count_off_1_cry_6\,
            clk => \N__20585\,
            ce => \N__19797\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_7_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12118\,
            in1 => \N__13354\,
            in2 => \_gnd_net_\,
            in3 => \N__11783\,
            lcout => \POWERLED.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_6\,
            carryout => \POWERLED.un1_count_off_1_cry_7\,
            clk => \N__20585\,
            ce => \N__19797\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_8_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12111\,
            in1 => \N__12193\,
            in2 => \_gnd_net_\,
            in3 => \N__11780\,
            lcout => \POWERLED.count_offZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => \POWERLED.un1_count_off_1_cry_8\,
            clk => \N__20604\,
            ce => \N__19807\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_9_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12114\,
            in1 => \N__12163\,
            in2 => \_gnd_net_\,
            in3 => \N__11930\,
            lcout => \POWERLED.count_offZ0Z_9\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_8\,
            carryout => \POWERLED.un1_count_off_1_cry_9\,
            clk => \N__20604\,
            ce => \N__19807\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_10_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12108\,
            in1 => \N__11813\,
            in2 => \_gnd_net_\,
            in3 => \N__11927\,
            lcout => \POWERLED.count_offZ0Z_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_9\,
            carryout => \POWERLED.un1_count_off_1_cry_10\,
            clk => \N__20604\,
            ce => \N__19807\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_11_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12112\,
            in1 => \N__11855\,
            in2 => \_gnd_net_\,
            in3 => \N__11924\,
            lcout => \POWERLED.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_10\,
            carryout => \POWERLED.un1_count_off_1_cry_11\,
            clk => \N__20604\,
            ce => \N__19807\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_12_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12109\,
            in1 => \N__11909\,
            in2 => \_gnd_net_\,
            in3 => \N__11921\,
            lcout => \POWERLED.count_offZ0Z_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_11\,
            carryout => \POWERLED.un1_count_off_1_cry_12\,
            clk => \N__20604\,
            ce => \N__19807\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_13_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12113\,
            in1 => \N__11897\,
            in2 => \_gnd_net_\,
            in3 => \N__11918\,
            lcout => \POWERLED.count_offZ0Z_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_12\,
            carryout => \POWERLED.un1_count_off_1_cry_13\,
            clk => \N__20604\,
            ce => \N__19807\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_14_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12110\,
            in1 => \N__11827\,
            in2 => \_gnd_net_\,
            in3 => \N__11915\,
            lcout => \POWERLED.count_offZ0Z_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_13\,
            carryout => \POWERLED.un1_count_off_1_cry_14\,
            clk => \N__20604\,
            ce => \N__19807\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_15_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12115\,
            in1 => \N__11884\,
            in2 => \_gnd_net_\,
            in3 => \N__11912\,
            lcout => \POWERLED.count_offZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20604\,
            ce => \N__19807\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIAJ6S_15_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11908\,
            in1 => \N__11896\,
            in2 => \N__11885\,
            in3 => \N__11870\,
            lcout => \POWERLED.func_state_ns_0_a2_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI4D6S_10_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11854\,
            in1 => \N__11843\,
            in2 => \N__11828\,
            in3 => \N__11812\,
            lcout => \POWERLED.func_state_ns_0_a2_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI8GP11_5_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__12194\,
            in1 => \N__12179\,
            in2 => \N__12164\,
            in3 => \N__12149\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_ns_0_a2_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIIKVR3_10_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12134\,
            in1 => \N__12128\,
            in2 => \N__12122\,
            in3 => \N__13313\,
            lcout => \POWERLED.count_off_RNIIKVR3Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIHPO9A_0_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__13698\,
            in1 => \N__14901\,
            in2 => \_gnd_net_\,
            in3 => \N__13521\,
            lcout => \POWERLED.count_off_0_sqmuxa\,
            ltout => \POWERLED.count_off_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI9LL3G_1_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__14933\,
            in1 => \_gnd_net_\,
            in2 => \N__12068\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_85_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__13712\,
            in1 => \N__13528\,
            in2 => \N__13643\,
            in3 => \N__14906\,
            lcout => \POWERLED.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20605\,
            ce => \N__19808\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_1_cry_1_c_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12038\,
            in2 => \N__12016\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \POWERLED.un1_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_2_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20124\,
            in1 => \N__11986\,
            in2 => \_gnd_net_\,
            in3 => \N__11963\,
            lcout => \POWERLED.countZ0Z_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_1\,
            carryout => \POWERLED.un1_count_1_cry_2\,
            clk => \N__20596\,
            ce => 'H',
            sr => \N__12519\
        );

    \POWERLED.count_3_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20107\,
            in1 => \N__11956\,
            in2 => \_gnd_net_\,
            in3 => \N__11933\,
            lcout => \POWERLED.countZ0Z_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_2\,
            carryout => \POWERLED.un1_count_1_cry_3\,
            clk => \N__20596\,
            ce => 'H',
            sr => \N__12519\
        );

    \POWERLED.count_4_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20125\,
            in1 => \N__12472\,
            in2 => \_gnd_net_\,
            in3 => \N__12449\,
            lcout => \POWERLED.countZ0Z_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_3\,
            carryout => \POWERLED.un1_count_1_cry_4\,
            clk => \N__20596\,
            ce => 'H',
            sr => \N__12519\
        );

    \POWERLED.count_5_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20108\,
            in1 => \N__12442\,
            in2 => \_gnd_net_\,
            in3 => \N__12419\,
            lcout => \POWERLED.countZ0Z_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_4\,
            carryout => \POWERLED.un1_count_1_cry_5\,
            clk => \N__20596\,
            ce => 'H',
            sr => \N__12519\
        );

    \POWERLED.count_6_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20126\,
            in1 => \N__12412\,
            in2 => \_gnd_net_\,
            in3 => \N__12389\,
            lcout => \POWERLED.countZ0Z_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_5\,
            carryout => \POWERLED.un1_count_1_cry_6\,
            clk => \N__20596\,
            ce => 'H',
            sr => \N__12519\
        );

    \POWERLED.count_7_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20109\,
            in1 => \N__12377\,
            in2 => \_gnd_net_\,
            in3 => \N__12356\,
            lcout => \POWERLED.countZ0Z_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_6\,
            carryout => \POWERLED.un1_count_1_cry_7\,
            clk => \N__20596\,
            ce => 'H',
            sr => \N__12519\
        );

    \POWERLED.count_8_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20127\,
            in1 => \N__12352\,
            in2 => \_gnd_net_\,
            in3 => \N__12329\,
            lcout => \POWERLED.countZ0Z_8\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_7\,
            carryout => \POWERLED.un1_count_1_cry_8\,
            clk => \N__20596\,
            ce => 'H',
            sr => \N__12519\
        );

    \POWERLED.count_9_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20141\,
            in1 => \N__12321\,
            in2 => \_gnd_net_\,
            in3 => \N__12293\,
            lcout => \POWERLED.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \POWERLED.un1_count_1_cry_9\,
            clk => \N__20630\,
            ce => 'H',
            sr => \N__12515\
        );

    \POWERLED.count_10_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20150\,
            in1 => \N__12286\,
            in2 => \_gnd_net_\,
            in3 => \N__12263\,
            lcout => \POWERLED.countZ0Z_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_9\,
            carryout => \POWERLED.un1_count_1_cry_10\,
            clk => \N__20630\,
            ce => 'H',
            sr => \N__12515\
        );

    \POWERLED.count_11_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20139\,
            in1 => \N__12256\,
            in2 => \_gnd_net_\,
            in3 => \N__12230\,
            lcout => \POWERLED.countZ0Z_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_10\,
            carryout => \POWERLED.un1_count_1_cry_11\,
            clk => \N__20630\,
            ce => 'H',
            sr => \N__12515\
        );

    \POWERLED.count_12_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20151\,
            in1 => \N__12223\,
            in2 => \_gnd_net_\,
            in3 => \N__12197\,
            lcout => \POWERLED.countZ0Z_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_11\,
            carryout => \POWERLED.un1_count_1_cry_12\,
            clk => \N__20630\,
            ce => 'H',
            sr => \N__12515\
        );

    \POWERLED.count_13_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20140\,
            in1 => \N__12622\,
            in2 => \_gnd_net_\,
            in3 => \N__12599\,
            lcout => \POWERLED.countZ0Z_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_12\,
            carryout => \POWERLED.un1_count_1_cry_13\,
            clk => \N__20630\,
            ce => 'H',
            sr => \N__12515\
        );

    \POWERLED.count_14_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20152\,
            in1 => \N__12592\,
            in2 => \_gnd_net_\,
            in3 => \N__12566\,
            lcout => \POWERLED.countZ0Z_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_13\,
            carryout => \POWERLED.un1_count_1_cry_14\,
            clk => \N__20630\,
            ce => 'H',
            sr => \N__12515\
        );

    \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18301\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_14\,
            carryout => \POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__18318\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryout => \POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_esr_15_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12556\,
            in2 => \_gnd_net_\,
            in3 => \N__12563\,
            lcout => \POWERLED.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20635\,
            ce => \N__12533\,
            sr => \N__12520\
        );

    \HDA_STRAP.count_RNO_0_0_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13874\,
            in2 => \N__13928\,
            in3 => \N__13927\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_6_1_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_1_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13901\,
            in2 => \_gnd_net_\,
            in3 => \N__12482\,
            lcout => \HDA_STRAP.countZ0Z_1\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_0\,
            carryout => \HDA_STRAP.un1_count_1_cry_1\,
            clk => \N__20205\,
            ce => \N__19712\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_2_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13913\,
            in2 => \_gnd_net_\,
            in3 => \N__12479\,
            lcout => \HDA_STRAP.countZ0Z_2\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_1\,
            carryout => \HDA_STRAP.un1_count_1_cry_2\,
            clk => \N__20205\,
            ce => \N__19712\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_3_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13888\,
            in2 => \_gnd_net_\,
            in3 => \N__12659\,
            lcout => \HDA_STRAP.countZ0Z_3\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_2\,
            carryout => \HDA_STRAP.un1_count_1_cry_3\,
            clk => \N__20205\,
            ce => \N__19712\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_4_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13766\,
            in2 => \_gnd_net_\,
            in3 => \N__12656\,
            lcout => \HDA_STRAP.countZ0Z_4\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_3\,
            carryout => \HDA_STRAP.un1_count_1_cry_4\,
            clk => \N__20205\,
            ce => \N__19712\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_5_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13793\,
            in2 => \_gnd_net_\,
            in3 => \N__12653\,
            lcout => \HDA_STRAP.countZ0Z_5\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_4\,
            carryout => \HDA_STRAP.un1_count_1_cry_5\,
            clk => \N__20205\,
            ce => \N__19712\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_6_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15686\,
            in2 => \_gnd_net_\,
            in3 => \N__12650\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_5\,
            carryout => \HDA_STRAP.un1_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_7_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13805\,
            in2 => \_gnd_net_\,
            in3 => \N__12647\,
            lcout => \HDA_STRAP.countZ0Z_7\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_6\,
            carryout => \HDA_STRAP.un1_count_1_cry_7\,
            clk => \N__20205\,
            ce => \N__19712\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_8_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13958\,
            in2 => \_gnd_net_\,
            in3 => \N__12644\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_6_2_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_9_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13780\,
            in2 => \_gnd_net_\,
            in3 => \N__12641\,
            lcout => \HDA_STRAP.countZ0Z_9\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_8\,
            carryout => \HDA_STRAP.un1_count_1_cry_9\,
            clk => \N__20370\,
            ce => \N__19741\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_10_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14011\,
            in2 => \_gnd_net_\,
            in3 => \N__12638\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_9\,
            carryout => \HDA_STRAP.un1_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_11_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13753\,
            in2 => \_gnd_net_\,
            in3 => \N__12629\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_10\,
            carryout => \HDA_STRAP.un1_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_12_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13832\,
            in2 => \_gnd_net_\,
            in3 => \N__12776\,
            lcout => \HDA_STRAP.countZ0Z_12\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_11\,
            carryout => \HDA_STRAP.un1_count_1_cry_12\,
            clk => \N__20370\,
            ce => \N__19741\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_13_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13817\,
            in2 => \_gnd_net_\,
            in3 => \N__12773\,
            lcout => \HDA_STRAP.countZ0Z_13\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_12\,
            carryout => \HDA_STRAP.un1_count_1_cry_13\,
            clk => \N__20370\,
            ce => \N__19741\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_14_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13859\,
            in2 => \_gnd_net_\,
            in3 => \N__12770\,
            lcout => \HDA_STRAP.countZ0Z_14\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_13\,
            carryout => \HDA_STRAP.un1_count_1_cry_14\,
            clk => \N__20370\,
            ce => \N__19741\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_15_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13846\,
            in2 => \_gnd_net_\,
            in3 => \N__12767\,
            lcout => \HDA_STRAP.countZ0Z_15\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_14\,
            carryout => \HDA_STRAP.un1_count_1_cry_15\,
            clk => \N__20370\,
            ce => \N__19741\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_16_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13994\,
            in2 => \_gnd_net_\,
            in3 => \N__12764\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNO_0_17_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13976\,
            in2 => \_gnd_net_\,
            in3 => \N__12761\,
            lcout => \HDA_STRAP.count_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIVL3D_0_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14658\,
            in2 => \N__14194\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_dutycycle_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_6_5_0_\,
            carryout => \POWERLED.un1_dutycycle_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12740\,
            in3 => \N__12707\,
            lcout => \POWERLED.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_0\,
            carryout => \POWERLED.un1_dutycycle_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12704\,
            in2 => \N__12698\,
            in3 => \N__12662\,
            lcout => \POWERLED.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_1\,
            carryout => \POWERLED.un1_dutycycle_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14261\,
            in2 => \N__14278\,
            in3 => \N__12986\,
            lcout => \POWERLED.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_2\,
            carryout => \POWERLED.un1_dutycycle_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14225\,
            in2 => \N__14243\,
            in3 => \N__12962\,
            lcout => \POWERLED.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_3\,
            carryout => \POWERLED.un1_dutycycle_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14219\,
            in2 => \N__12959\,
            in3 => \N__12929\,
            lcout => \POWERLED.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_4\,
            carryout => \POWERLED.un1_dutycycle_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12926\,
            in2 => \N__13025\,
            in3 => \N__12893\,
            lcout => \POWERLED.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_5\,
            carryout => \POWERLED.un1_dutycycle_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12890\,
            in2 => \N__13202\,
            in3 => \N__12851\,
            lcout => \POWERLED.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_6\,
            carryout => \POWERLED.un1_dutycycle_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13250\,
            in2 => \N__13235\,
            in3 => \N__12821\,
            lcout => \POWERLED.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => \POWERLED.un1_dutycycle_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13271\,
            in2 => \N__14315\,
            in3 => \N__12797\,
            lcout => \POWERLED.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_8\,
            carryout => \POWERLED.un1_dutycycle_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13289\,
            in2 => \N__13301\,
            in3 => \N__12779\,
            lcout => \POWERLED.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_9\,
            carryout => \POWERLED.un1_dutycycle_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13376\,
            in2 => \N__16493\,
            in3 => \N__13163\,
            lcout => \POWERLED.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_10\,
            carryout => \POWERLED.un1_dutycycle_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13385\,
            in2 => \N__13400\,
            in3 => \N__13142\,
            lcout => \POWERLED.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_11\,
            carryout => \POWERLED.un1_dutycycle_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13481\,
            in2 => \N__13946\,
            in3 => \N__13121\,
            lcout => \POWERLED.mult1_un54_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_12\,
            carryout => \POWERLED.un1_dutycycle_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13277\,
            in2 => \N__13937\,
            in3 => \N__13100\,
            lcout => \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_13\,
            carryout => \POWERLED.un1_dutycycle_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13283\,
            in2 => \N__13493\,
            in3 => \N__13076\,
            lcout => \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_14\,
            carryout => \POWERLED.un1_dutycycle_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16128\,
            in2 => \N__13265\,
            in3 => \N__13058\,
            lcout => \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71\,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => \POWERLED.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.CO2_THRU_LUT4_0_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13055\,
            lcout => \POWERLED.CO2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNI8MSK_5_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__16066\,
            in1 => \N__14601\,
            in2 => \_gnd_net_\,
            in3 => \N__13043\,
            lcout => \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIE4FL_9_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__16388\,
            in1 => \N__16237\,
            in2 => \_gnd_net_\,
            in3 => \N__16068\,
            lcout => \POWERLED.dutycycle_RNIE4FLZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI53MG_14_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16339\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16460\,
            lcout => \POWERLED.dutycycle_RNI53MGZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNI2GSK_6_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14644\,
            in2 => \N__13223\,
            in3 => \N__14722\,
            lcout => \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI84C11_14_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101101111000"
        )
    port map (
            in0 => \N__16458\,
            in1 => \N__16389\,
            in2 => \N__16345\,
            in3 => \N__16459\,
            lcout => \POWERLED.dutycycle_RNI84C11Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIB1FL_8_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__14393\,
            in1 => \N__16185\,
            in2 => \_gnd_net_\,
            in3 => \N__16067\,
            lcout => \POWERLED.dutycycle_RNIB1FLZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI75MG_15_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__16117\,
            in1 => \_gnd_net_\,
            in2 => \N__16344\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI75MGZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIM0TE_8_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16065\,
            in2 => \_gnd_net_\,
            in3 => \N__16167\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_1_34_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIUUB41_6_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000101111000"
        )
    port map (
            in0 => \N__16281\,
            in1 => \N__14445\,
            in2 => \N__13256\,
            in3 => \N__14373\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_1_axb_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJL1R1_6_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13253\,
            in3 => \N__13246\,
            lcout => \POWERLED.dutycycle_RNIJL1R1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNIBPSK_6_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__16231\,
            in1 => \N__14523\,
            in2 => \_gnd_net_\,
            in3 => \N__13222\,
            lcout => \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2V0P_10_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__16173\,
            in1 => \N__16330\,
            in2 => \_gnd_net_\,
            in3 => \N__16283\,
            lcout => \POWERLED.dutycycle_RNI2V0PZ0Z_10\,
            ltout => \POWERLED.dutycycle_RNI2V0PZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI712I1_15_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__16116\,
            in1 => \N__16172\,
            in2 => \N__13388\,
            in3 => \N__16394\,
            lcout => \POWERLED.dutycycle_RNI712I1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQ09G1_10_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__16489\,
            in1 => \N__16329\,
            in2 => \N__16184\,
            in3 => \N__16282\,
            lcout => \POWERLED.dutycycle_RNIQ09G1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_0_2_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111011101110"
        )
    port map (
            in0 => \N__15359\,
            in1 => \N__15098\,
            in2 => \N__16590\,
            in3 => \N__15298\,
            lcout => \POWERLED.dutycycle_lm_0_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIS3P11_2_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__13366\,
            in1 => \N__13355\,
            in2 => \N__13340\,
            in3 => \N__13324\,
            lcout => \POWERLED.func_state_ns_0_a2_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI1DHM_6_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__18055\,
            in1 => \N__18007\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_368_0_i_i_a6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI1VLG_10_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16284\,
            in2 => \_gnd_net_\,
            in3 => \N__16448\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_1_44_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIF3561_9_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \N__16082\,
            in1 => \N__16236\,
            in2 => \N__13304\,
            in3 => \N__16393\,
            lcout => \POWERLED.dutycycle_RNIF3561Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIC8C11_15_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001101101100"
        )
    port map (
            in0 => \N__16334\,
            in1 => \N__16118\,
            in2 => \N__16466\,
            in3 => \N__16335\,
            lcout => \POWERLED.dutycycle_RNIC8C11Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI73C11_15_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \N__16465\,
            in1 => \N__16168\,
            in2 => \N__16402\,
            in3 => \N__16115\,
            lcout => \POWERLED.dutycycle_RNI73C11Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIBR4E9_6_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16676\,
            in1 => \N__13606\,
            in2 => \N__13469\,
            in3 => \N__16630\,
            lcout => \POWERLED.N_177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIAA8L4_0_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101110"
        )
    port map (
            in0 => \N__13548\,
            in1 => \N__15220\,
            in2 => \N__14306\,
            in3 => \N__16000\,
            lcout => \POWERLED.N_200_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIS0FM9_7_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__13701\,
            in1 => \N__16631\,
            in2 => \N__13442\,
            in3 => \N__18019\,
            lcout => OPEN,
            ltout => \POWERLED.N_207_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI5LMRL_1_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__14762\,
            in1 => \N__16814\,
            in2 => \N__13460\,
            in3 => \N__14926\,
            lcout => \POWERLED.N_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIG4MR5_1_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__15300\,
            in1 => \N__16652\,
            in2 => \_gnd_net_\,
            in3 => \N__15147\,
            lcout => \POWERLED.N_149\,
            ltout => \POWERLED.N_149_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIJ13KB_7_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__18018\,
            in1 => \N__15651\,
            in2 => \N__13433\,
            in3 => \N__15419\,
            lcout => \POWERLED.un2_slp_s3n_2_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5J285_5_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__13702\,
            in1 => \N__16001\,
            in2 => \N__15446\,
            in3 => \N__13549\,
            lcout => \POWERLED.N_214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI0AN05_0_0_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__15996\,
            in1 => \N__13683\,
            in2 => \N__15223\,
            in3 => \N__14304\,
            lcout => \POWERLED.N_248\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_2_0_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__15282\,
            in1 => \N__13556\,
            in2 => \N__13700\,
            in3 => \N__15999\,
            lcout => \POWERLED.N_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI1UHM1_0_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000100"
        )
    port map (
            in0 => \N__16581\,
            in1 => \N__15093\,
            in2 => \N__15224\,
            in3 => \N__15636\,
            lcout => \POWERLED.N_213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3T7Q4_5_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__15635\,
            in1 => \N__13555\,
            in2 => \N__15445\,
            in3 => \N__15997\,
            lcout => OPEN,
            ltout => \POWERLED.N_218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNITEUV5_5_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__15350\,
            in1 => \_gnd_net_\,
            in2 => \N__13532\,
            in3 => \N__15010\,
            lcout => \POWERLED.count_clk_1_sqmuxa_5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI9HME_1_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15212\,
            in2 => \_gnd_net_\,
            in3 => \N__15258\,
            lcout => \POWERLED.N_88\,
            ltout => \POWERLED.N_88_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIIA93A_0_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111001100"
        )
    port map (
            in0 => \N__15137\,
            in1 => \N__13517\,
            in2 => \N__13496\,
            in3 => \N__15011\,
            lcout => \POWERLED.count_clk_1_sqmuxa_5_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI0AN05_0_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__14305\,
            in1 => \N__15216\,
            in2 => \N__13699\,
            in3 => \N__15998\,
            lcout => \POWERLED.N_250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_1_sqmuxa_5_0_a2_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__15002\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15355\,
            lcout => \POWERLED.N_228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_1_0_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__15356\,
            in1 => \N__15211\,
            in2 => \N__15161\,
            in3 => \N__15003\,
            lcout => \POWERLED.N_179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_3_1_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15091\,
            in1 => \N__15104\,
            in2 => \N__16591\,
            in3 => \N__15645\,
            lcout => OPEN,
            ltout => \POWERLED.N_208_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_1_1_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__13655\,
            in1 => \N__16583\,
            in2 => \N__13715\,
            in3 => \N__14897\,
            lcout => \POWERLED.func_state_ns_i_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_ns_0_i_0_0_a2_0_0_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__15092\,
            in1 => \N__15357\,
            in2 => \_gnd_net_\,
            in3 => \N__20708\,
            lcout => \POWERLED.N_222\,
            ltout => \POWERLED.N_222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_2_1_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15294\,
            in1 => \N__15210\,
            in2 => \N__13658\,
            in3 => \N__15148\,
            lcout => OPEN,
            ltout => \POWERLED.N_211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_0_1_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13654\,
            in2 => \N__13646\,
            in3 => \N__15374\,
            lcout => \POWERLED.func_state_ns_i_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_0_0_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__15646\,
            in1 => \N__15090\,
            in2 => \N__14902\,
            in3 => \N__16582\,
            lcout => \POWERLED.N_178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13634\,
            in1 => \N__13628\,
            in2 => \N__13622\,
            in3 => \N__13610\,
            lcout => \POWERLED.func_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20534\,
            ce => \N__19806\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_1_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100100010"
        )
    port map (
            in0 => \N__15512\,
            in1 => \N__15584\,
            in2 => \N__18881\,
            in3 => \N__15542\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20593\,
            ce => \N__19811\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_0_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15541\,
            in2 => \_gnd_net_\,
            in3 => \N__15583\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20593\,
            ce => \N__19811\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIH91A_0_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15879\,
            in2 => \_gnd_net_\,
            in3 => \N__15809\,
            lcout => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIQC821_0_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13912\,
            in1 => \N__13900\,
            in2 => \N__13889\,
            in3 => \N__13873\,
            lcout => \HDA_STRAP.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIDLB61_6_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__13858\,
            in1 => \N__13957\,
            in2 => \N__13847\,
            in3 => \N__15679\,
            lcout => OPEN,
            ltout => \HDA_STRAP.un4_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIUKIR1_12_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__13831\,
            in1 => \_gnd_net_\,
            in2 => \N__13820\,
            in3 => \N__13816\,
            lcout => \HDA_STRAP.un4_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNID0921_4_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13804\,
            in1 => \N__13792\,
            in2 => \N__13781\,
            in3 => \N__13765\,
            lcout => \HDA_STRAP.un4_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI63EA1_17_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13993\,
            in1 => \N__13754\,
            in2 => \N__14015\,
            in3 => \N__13975\,
            lcout => OPEN,
            ltout => \HDA_STRAP.un4_count_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIB5IA5_0_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13739\,
            in1 => \N__13733\,
            in2 => \N__13727\,
            in3 => \N__13724\,
            lcout => \HDA_STRAP.count_RNIB5IA5Z0Z_0\,
            ltout => \HDA_STRAP.count_RNIB5IA5Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_0_2_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__15902\,
            in1 => \_gnd_net_\,
            in2 => \N__13718\,
            in3 => \N__15810\,
            lcout => \HDA_STRAP.curr_state_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_10_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011110000"
        )
    port map (
            in0 => \N__15811\,
            in1 => \N__15904\,
            in2 => \N__14024\,
            in3 => \N__15723\,
            lcout => \HDA_STRAP.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20341\,
            ce => \N__19762\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_16_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__15722\,
            in1 => \N__14000\,
            in2 => \N__15915\,
            in3 => \N__15814\,
            lcout => \HDA_STRAP.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20341\,
            ce => \N__19762\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_17_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__15812\,
            in1 => \N__13982\,
            in2 => \N__15916\,
            in3 => \N__15724\,
            lcout => \HDA_STRAP.countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20341\,
            ce => \N__19762\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_8_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__15813\,
            in1 => \N__13964\,
            in2 => \N__15917\,
            in3 => \N__15725\,
            lcout => \HDA_STRAP.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20341\,
            ce => \N__19762\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI8M7Q_2_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__14726\,
            in1 => \N__14602\,
            in2 => \N__14665\,
            in3 => \N__14394\,
            lcout => \POWERLED.un2_slp_s3n_2_0_o2_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI31MG_0_12_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16467\,
            in2 => \_gnd_net_\,
            in3 => \N__16398\,
            lcout => \POWERLED.dutycycle_RNI31MG_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI31MG_12_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__16468\,
            in1 => \_gnd_net_\,
            in2 => \N__16403\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI31MGZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIO2TE_9_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16243\,
            in2 => \_gnd_net_\,
            in3 => \N__16397\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_1_39_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI34C41_8_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__16186\,
            in1 => \N__14395\,
            in2 => \N__14318\,
            in3 => \N__16080\,
            lcout => \POWERLED.dutycycle_RNI34C41Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI4I7Q_5_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__14119\,
            in1 => \N__14195\,
            in2 => \N__14543\,
            in3 => \N__14455\,
            lcout => \POWERLED.N_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIK4I81_6_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__14645\,
            in1 => \N__14279\,
            in2 => \N__14740\,
            in3 => \N__14454\,
            lcout => \POWERLED.dutycycle_RNIK4I81Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_2_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__14675\,
            in1 => \N__16761\,
            in2 => \N__14255\,
            in3 => \N__20716\,
            lcout => \POWERLED.dutycycleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20384\,
            ce => \N__19749\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQAI81_4_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__14239\,
            in1 => \N__14585\,
            in2 => \N__14399\,
            in3 => \N__14646\,
            lcout => \POWERLED.dutycycle_RNIQAI81Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOQLJ_4_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__14586\,
            in1 => \N__14392\,
            in2 => \_gnd_net_\,
            in3 => \N__14647\,
            lcout => \POWERLED.dutycycle_RNIOQLJZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15388\,
            in2 => \N__15392\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \POWERLED.dutycycle_cry_c_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_0_0_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14836\,
            in2 => \N__14213\,
            in3 => \N__14132\,
            lcout => \POWERLED.dutycycle_s_0\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_c_0_THRU_CO\,
            carryout => \POWERLED.dutycycle_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_0_1_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14128\,
            in2 => \N__14853\,
            in3 => \N__14039\,
            lcout => \POWERLED.dutycycle_s_1\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_0\,
            carryout => \POWERLED.dutycycle_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_1_2_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14840\,
            in2 => \N__14741\,
            in3 => \N__14669\,
            lcout => \POWERLED.dutycycle_s_2\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_1\,
            carryout => \POWERLED.dutycycle_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_3_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__16772\,
            in1 => \N__14654\,
            in2 => \N__14854\,
            in3 => \N__14609\,
            lcout => \POWERLED.dutycycleZ0Z_3\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_2\,
            carryout => \POWERLED.dutycycle_cry_3\,
            clk => \N__20450\,
            ce => \N__19786\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_4_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__16760\,
            in1 => \N__14844\,
            in2 => \N__14603\,
            in3 => \N__14546\,
            lcout => \POWERLED.dutycycleZ0Z_4\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_3\,
            carryout => \POWERLED.dutycycle_cry_4\,
            clk => \N__20450\,
            ce => \N__19786\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_cry_c_RNIV95M9_4_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14542\,
            in2 => \N__14855\,
            in3 => \N__14462\,
            lcout => \POWERLED.dutycycle_s_5\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_4\,
            carryout => \POWERLED.dutycycle_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_cry_c_RNI1C5M9_5_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14848\,
            in2 => \N__14459\,
            in3 => \N__14402\,
            lcout => \POWERLED.dutycycle_s_6\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_5\,
            carryout => \POWERLED.dutycycle_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_7_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__16758\,
            in1 => \N__14820\,
            in2 => \N__14396\,
            in3 => \N__14327\,
            lcout => \POWERLED.dutycycleZ0Z_7\,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => \POWERLED.dutycycle_cry_7\,
            clk => \N__20473\,
            ce => \N__19774\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_8_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__16738\,
            in1 => \N__16073\,
            in2 => \N__14849\,
            in3 => \N__14324\,
            lcout => \POWERLED.dutycycleZ0Z_8\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_7\,
            carryout => \POWERLED.dutycycle_cry_8\,
            clk => \N__20473\,
            ce => \N__19774\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_9_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__16759\,
            in1 => \N__14824\,
            in2 => \N__16244\,
            in3 => \N__14321\,
            lcout => \POWERLED.dutycycleZ0Z_9\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_8\,
            carryout => \POWERLED.dutycycle_cry_9\,
            clk => \N__20473\,
            ce => \N__19774\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_10_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__16735\,
            in1 => \N__16287\,
            in2 => \N__14850\,
            in3 => \N__14870\,
            lcout => \POWERLED.dutycycleZ0Z_10\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_9\,
            carryout => \POWERLED.dutycycle_cry_10\,
            clk => \N__20473\,
            ce => \N__19774\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_11_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__16756\,
            in1 => \N__14828\,
            in2 => \N__16187\,
            in3 => \N__14867\,
            lcout => \POWERLED.dutycycleZ0Z_11\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_10\,
            carryout => \POWERLED.dutycycle_cry_11\,
            clk => \N__20473\,
            ce => \N__19774\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_12_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__16736\,
            in1 => \N__16396\,
            in2 => \N__14851\,
            in3 => \N__14864\,
            lcout => \POWERLED.dutycycleZ0Z_12\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_11\,
            carryout => \POWERLED.dutycycle_cry_12\,
            clk => \N__20473\,
            ce => \N__19774\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_13_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__16757\,
            in1 => \N__14832\,
            in2 => \N__16469\,
            in3 => \N__14861\,
            lcout => \POWERLED.dutycycleZ0Z_13\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_12\,
            carryout => \POWERLED.dutycycle_cry_13\,
            clk => \N__20473\,
            ce => \N__19774\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_14_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__16737\,
            in1 => \N__16343\,
            in2 => \N__14852\,
            in3 => \N__14858\,
            lcout => \POWERLED.dutycycleZ0Z_14\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_13\,
            carryout => \POWERLED.dutycycle_cry_14\,
            clk => \N__20473\,
            ce => \N__19774\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_15_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__16739\,
            in1 => \N__14804\,
            in2 => \N__16130\,
            in3 => \N__14768\,
            lcout => \POWERLED.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20451\,
            ce => \N__19785\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI33DK1_1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__15299\,
            in1 => \N__15222\,
            in2 => \N__15097\,
            in3 => \N__15648\,
            lcout => \POWERLED.N_246\,
            ltout => \POWERLED.N_246_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIS9OC3_1_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14765\,
            in3 => \N__16645\,
            lcout => \POWERLED.N_203_4\,
            ltout => \POWERLED.N_203_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI09QT9_1_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__16607\,
            in1 => \N__16825\,
            in2 => \N__14756\,
            in3 => \N__15162\,
            lcout => OPEN,
            ltout => \POWERLED.N_203_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNITU0DB_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__15650\,
            in1 => \N__15086\,
            in2 => \N__14960\,
            in3 => \N__16556\,
            lcout => \POWERLED.count_clk_139_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI2M0Q4_6_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__18056\,
            in1 => \N__15649\,
            in2 => \N__16672\,
            in3 => \N__16623\,
            lcout => \POWERLED.N_251\,
            ltout => \POWERLED.N_251_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI01TCL_7_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__18020\,
            in1 => \N__14912\,
            in2 => \N__14957\,
            in3 => \N__14954\,
            lcout => OPEN,
            ltout => \POWERLED.un2_slp_s3n_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIOH1J11_7_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14948\,
            in2 => \N__14942\,
            in3 => \N__20056\,
            lcout => \POWERLED.count_clk_RNIOH1J11Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIORSP5_1_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15163\,
            in1 => \N__16557\,
            in2 => \_gnd_net_\,
            in3 => \N__14939\,
            lcout => \POWERLED.N_205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIA8VP_7_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18016\,
            in2 => \_gnd_net_\,
            in3 => \N__15372\,
            lcout => OPEN,
            ltout => \POWERLED.un2_slp_s3n_2_0_a6_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIAIGJ4_7_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111010"
        )
    port map (
            in0 => \N__15012\,
            in1 => \N__15643\,
            in2 => \N__14915\,
            in3 => \N__16629\,
            lcout => \POWERLED.un2_slp_s3n_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI7LE01_7_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__15083\,
            in1 => \N__18017\,
            in2 => \_gnd_net_\,
            in3 => \N__15221\,
            lcout => \POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNINTA34_1_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15301\,
            in2 => \_gnd_net_\,
            in3 => \N__15157\,
            lcout => \POWERLED.N_127\,
            ltout => \POWERLED.N_127_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIUIEUK_1_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__15644\,
            in1 => \N__15461\,
            in2 => \N__15455\,
            in3 => \N__15452\,
            lcout => \POWERLED.count_clk_1_sqmuxa_5_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIH2SJ1_1_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100011001"
        )
    port map (
            in0 => \N__15351\,
            in1 => \N__15085\,
            in2 => \N__16577\,
            in3 => \N__15438\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_3_sqmuxa_1_i_0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI6KL57_0_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110100"
        )
    port map (
            in0 => \N__15084\,
            in1 => \N__15373\,
            in2 => \N__15422\,
            in3 => \N__15418\,
            lcout => \POWERLED.N_366_1\,
            ltout => \POWERLED.N_366_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI446AD_7_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110011"
        )
    port map (
            in0 => \N__15407\,
            in1 => \N__20704\,
            in2 => \N__15401\,
            in3 => \N__15398\,
            lcout => \POWERLED.dutycycle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI9HME_0_1_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15289\,
            in2 => \_gnd_net_\,
            in3 => \N__15208\,
            lcout => \POWERLED.N_243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.N_55_i_i_o6_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__15358\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20702\,
            lcout => \N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_4_1_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15293\,
            in1 => \N__15209\,
            in2 => \_gnd_net_\,
            in3 => \N__15164\,
            lcout => \POWERLED.N_148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_EN_i_i_0_a2_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20703\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15057\,
            lcout => vccst_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNIJKKQ_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__15647\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15554\,
            lcout => vpp_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__15582\,
            in1 => \N__15508\,
            in2 => \_gnd_net_\,
            in3 => \N__15540\,
            lcout => \VPP_VDDQ.G_127_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNIDNTT1_0_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__15507\,
            in1 => \N__15538\,
            in2 => \_gnd_net_\,
            in3 => \N__15581\,
            lcout => \VPP_VDDQ.N_108_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__19555\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15652\,
            lcout => \VPP_VDDQ.N_238\,
            ltout => \VPP_VDDQ.N_238_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNINMKE1_1_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15566\,
            in3 => \N__15537\,
            lcout => \VPP_VDDQ.N_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100010101010"
        )
    port map (
            in0 => \N__15553\,
            in1 => \N__15509\,
            in2 => \N__15482\,
            in3 => \N__20083\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__20084\,
            in1 => \_gnd_net_\,
            in2 => \N__15563\,
            in3 => \N__15560\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20547\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNI8I855_0_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15510\,
            in1 => \N__15539\,
            in2 => \_gnd_net_\,
            in3 => \N__18877\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.N_154_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNIGR9S7_0_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__15511\,
            in1 => \N__15475\,
            in2 => \N__15464\,
            in3 => \N__20062\,
            lcout => \VPP_VDDQ.curr_state_RNIGR9S7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNO_0_15_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16923\,
            in2 => \_gnd_net_\,
            in3 => \N__20078\,
            lcout => \VPP_VDDQ.N_65_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_6_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19444\,
            in1 => \_gnd_net_\,
            in2 => \N__17027\,
            in3 => \N__17009\,
            lcout => \COUNTER.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20206\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_5_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__17050\,
            in1 => \N__17036\,
            in2 => \_gnd_net_\,
            in3 => \N__19443\,
            lcout => \COUNTER.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20206\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19445\,
            in1 => \N__16909\,
            in2 => \_gnd_net_\,
            in3 => \N__17591\,
            lcout => \COUNTER.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20206\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_RNO_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__17022\,
            in1 => \N__17049\,
            in2 => \N__17000\,
            in3 => \N__16908\,
            lcout => \COUNTER.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_6_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010101010"
        )
    port map (
            in0 => \N__15929\,
            in1 => \N__15903\,
            in2 => \N__15818\,
            in3 => \N__15721\,
            lcout => \HDA_STRAP.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20377\,
            ce => \N__19742\,
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20118\,
            in1 => \N__17345\,
            in2 => \N__19384\,
            in3 => \N__19385\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_5_0_\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_0\,
            clk => \N__20533\,
            ce => 'H',
            sr => \N__17891\
        );

    \ALL_SYS_PWRGD.count_1_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20103\,
            in1 => \N__17384\,
            in2 => \_gnd_net_\,
            in3 => \N__15668\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_0\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_1\,
            clk => \N__20533\,
            ce => 'H',
            sr => \N__17891\
        );

    \ALL_SYS_PWRGD.count_2_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20119\,
            in1 => \N__17231\,
            in2 => \_gnd_net_\,
            in3 => \N__15665\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_1\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_2\,
            clk => \N__20533\,
            ce => 'H',
            sr => \N__17891\
        );

    \ALL_SYS_PWRGD.count_3_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20104\,
            in1 => \N__17258\,
            in2 => \_gnd_net_\,
            in3 => \N__15662\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_2\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_3\,
            clk => \N__20533\,
            ce => 'H',
            sr => \N__17891\
        );

    \ALL_SYS_PWRGD.count_4_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20120\,
            in1 => \N__17462\,
            in2 => \_gnd_net_\,
            in3 => \N__15956\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_3\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_4\,
            clk => \N__20533\,
            ce => 'H',
            sr => \N__17891\
        );

    \ALL_SYS_PWRGD.count_5_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20105\,
            in1 => \N__17270\,
            in2 => \_gnd_net_\,
            in3 => \N__15953\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_4\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_5\,
            clk => \N__20533\,
            ce => 'H',
            sr => \N__17891\
        );

    \ALL_SYS_PWRGD.count_6_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20121\,
            in1 => \N__17476\,
            in2 => \_gnd_net_\,
            in3 => \N__15950\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_5\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_6\,
            clk => \N__20533\,
            ce => 'H',
            sr => \N__17891\
        );

    \ALL_SYS_PWRGD.count_7_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20106\,
            in1 => \N__17501\,
            in2 => \_gnd_net_\,
            in3 => \N__15947\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_6\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_7\,
            clk => \N__20533\,
            ce => 'H',
            sr => \N__17891\
        );

    \ALL_SYS_PWRGD.count_8_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20082\,
            in1 => \N__17489\,
            in2 => \_gnd_net_\,
            in3 => \N__15944\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_8\,
            clk => \N__20472\,
            ce => 'H',
            sr => \N__17890\
        );

    \ALL_SYS_PWRGD.count_9_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20073\,
            in1 => \N__17372\,
            in2 => \_gnd_net_\,
            in3 => \N__15941\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_8\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_9\,
            clk => \N__20472\,
            ce => 'H',
            sr => \N__17890\
        );

    \ALL_SYS_PWRGD.count_10_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20079\,
            in1 => \N__17359\,
            in2 => \_gnd_net_\,
            in3 => \N__15938\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_9\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_10\,
            clk => \N__20472\,
            ce => 'H',
            sr => \N__17890\
        );

    \ALL_SYS_PWRGD.count_11_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20071\,
            in1 => \N__17245\,
            in2 => \_gnd_net_\,
            in3 => \N__15935\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_10\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_11\,
            clk => \N__20472\,
            ce => 'H',
            sr => \N__17890\
        );

    \ALL_SYS_PWRGD.count_12_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20080\,
            in1 => \N__17411\,
            in2 => \_gnd_net_\,
            in3 => \N__15932\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_11\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_12\,
            clk => \N__20472\,
            ce => 'H',
            sr => \N__17890\
        );

    \ALL_SYS_PWRGD.count_13_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20072\,
            in1 => \N__17425\,
            in2 => \_gnd_net_\,
            in3 => \N__16502\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_12\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_13\,
            clk => \N__20472\,
            ce => 'H',
            sr => \N__17890\
        );

    \ALL_SYS_PWRGD.count_14_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20081\,
            in1 => \N__17450\,
            in2 => \_gnd_net_\,
            in3 => \N__16499\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_13\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_14\,
            clk => \N__20472\,
            ce => 'H',
            sr => \N__17890\
        );

    \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18375\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_14\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_esr_15_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17438\,
            in2 => \_gnd_net_\,
            in3 => \N__16496\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20557\,
            ce => \N__17858\,
            sr => \N__17883\
        );

    \POWERLED.dutycycle_RNIO18N_9_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__16235\,
            in1 => \N__16452\,
            in2 => \_gnd_net_\,
            in3 => \N__16285\,
            lcout => \POWERLED.dutycycle_RNIO18NZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI51C11_10_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16461\,
            in1 => \N__16395\,
            in2 => \N__16346\,
            in3 => \N__16286\,
            lcout => \POWERLED.un2_slp_s3n_2_0_o2_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIH6QT_15_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16238\,
            in1 => \N__16180\,
            in2 => \N__16129\,
            in3 => \N__16072\,
            lcout => OPEN,
            ltout => \POWERLED.un2_slp_s3n_2_0_o2_3_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIUTDP2_2_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16022\,
            in2 => \N__16016\,
            in3 => \N__16013\,
            lcout => \POWERLED.N_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIROMF7_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16784\,
            in2 => \_gnd_net_\,
            in3 => \N__20715\,
            lcout => \POWERLED.un1_dutycycle_4_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIPG2D1_2_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18097\,
            in1 => \N__18115\,
            in2 => \N__17648\,
            in3 => \N__17950\,
            lcout => \POWERLED.N_177_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIP4HM_2_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18114\,
            in2 => \_gnd_net_\,
            in3 => \N__17643\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_0_sqmuxa_5_0_o2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIP6BO1_4_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__17949\,
            in1 => \N__18044\,
            in2 => \N__16655\,
            in3 => \N__18096\,
            lcout => \POWERLED.N_141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIKKV71_12_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18442\,
            in1 => \N__17680\,
            in2 => \N__18428\,
            in3 => \N__16598\,
            lcout => \POWERLED.N_136\,
            ltout => \POWERLED.N_136_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIHJP92_1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__17930\,
            in1 => \N__18077\,
            in2 => \N__16634\,
            in3 => \N__17666\,
            lcout => \POWERLED.N_146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIUL2D1_1_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__17667\,
            in1 => \N__17931\,
            in2 => \N__18006\,
            in3 => \N__18078\,
            lcout => \POWERLED.count_clk_0_sqmuxa_5_0_a6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_esr_RNO_0_15_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18233\,
            in2 => \_gnd_net_\,
            in3 => \N__20061\,
            lcout => \POWERLED.N_65_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_esr_RNIVU6L_15_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18409\,
            in1 => \N__18457\,
            in2 => \N__18281\,
            in3 => \N__17911\,
            lcout => \POWERLED.count_clk_0_sqmuxa_5_0_o2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI3G101_5_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17990\,
            in1 => \N__16537\,
            in2 => \_gnd_net_\,
            in3 => \N__18079\,
            lcout => OPEN,
            ltout => \POWERLED.count_off_1_sqmuxa_i_a6_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNILEIU2_1_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__17932\,
            in1 => \N__17668\,
            in2 => \N__16829\,
            in3 => \N__16826\,
            lcout => \POWERLED.count_off_1_sqmuxa_i_a6_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_0_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20142\,
            in1 => \N__18167\,
            in2 => \N__18491\,
            in3 => \N__18490\,
            lcout => \RSMRST_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_0\,
            clk => \N__20636\,
            ce => 'H',
            sr => \N__18530\
        );

    \RSMRST_PWRGD.count_1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20132\,
            in1 => \N__18551\,
            in2 => \_gnd_net_\,
            in3 => \N__16805\,
            lcout => \RSMRST_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_0\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_1\,
            clk => \N__20636\,
            ce => 'H',
            sr => \N__18530\
        );

    \RSMRST_PWRGD.count_2_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20143\,
            in1 => \N__18578\,
            in2 => \_gnd_net_\,
            in3 => \N__16802\,
            lcout => \RSMRST_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_1\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_2\,
            clk => \N__20636\,
            ce => 'H',
            sr => \N__18530\
        );

    \RSMRST_PWRGD.count_3_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20133\,
            in1 => \N__18608\,
            in2 => \_gnd_net_\,
            in3 => \N__16799\,
            lcout => \RSMRST_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_2\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_3\,
            clk => \N__20636\,
            ce => 'H',
            sr => \N__18530\
        );

    \RSMRST_PWRGD.count_4_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20144\,
            in1 => \N__18590\,
            in2 => \_gnd_net_\,
            in3 => \N__16796\,
            lcout => \RSMRST_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_3\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_4\,
            clk => \N__20636\,
            ce => 'H',
            sr => \N__18530\
        );

    \RSMRST_PWRGD.count_5_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20134\,
            in1 => \N__18565\,
            in2 => \_gnd_net_\,
            in3 => \N__16793\,
            lcout => \RSMRST_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_4\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_5\,
            clk => \N__20636\,
            ce => 'H',
            sr => \N__18530\
        );

    \RSMRST_PWRGD.count_6_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20145\,
            in1 => \N__18179\,
            in2 => \_gnd_net_\,
            in3 => \N__16790\,
            lcout => \RSMRST_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_5\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_6\,
            clk => \N__20636\,
            ce => 'H',
            sr => \N__18530\
        );

    \RSMRST_PWRGD.count_7_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20135\,
            in1 => \N__18623\,
            in2 => \_gnd_net_\,
            in3 => \N__16787\,
            lcout => \RSMRST_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_6\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_7\,
            clk => \N__20636\,
            ce => 'H',
            sr => \N__18530\
        );

    \RSMRST_PWRGD.count_8_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20149\,
            in1 => \N__18155\,
            in2 => \_gnd_net_\,
            in3 => \N__16853\,
            lcout => \RSMRST_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_8\,
            clk => \N__20631\,
            ce => 'H',
            sr => \N__18529\
        );

    \RSMRST_PWRGD.count_9_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20138\,
            in1 => \N__18142\,
            in2 => \_gnd_net_\,
            in3 => \N__16850\,
            lcout => \RSMRST_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_8\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_9\,
            clk => \N__20631\,
            ce => 'H',
            sr => \N__18529\
        );

    \RSMRST_PWRGD.count_10_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20146\,
            in1 => \N__18206\,
            in2 => \_gnd_net_\,
            in3 => \N__16847\,
            lcout => \RSMRST_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_9\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_10\,
            clk => \N__20631\,
            ce => 'H',
            sr => \N__18529\
        );

    \RSMRST_PWRGD.count_11_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20136\,
            in1 => \N__18218\,
            in2 => \_gnd_net_\,
            in3 => \N__16844\,
            lcout => \RSMRST_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_10\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_11\,
            clk => \N__20631\,
            ce => 'H',
            sr => \N__18529\
        );

    \RSMRST_PWRGD.count_12_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20147\,
            in1 => \N__18128\,
            in2 => \_gnd_net_\,
            in3 => \N__16841\,
            lcout => \RSMRST_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_11\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_12\,
            clk => \N__20631\,
            ce => 'H',
            sr => \N__18529\
        );

    \RSMRST_PWRGD.count_13_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20137\,
            in1 => \N__18193\,
            in2 => \_gnd_net_\,
            in3 => \N__16838\,
            lcout => \RSMRST_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_12\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_13\,
            clk => \N__20631\,
            ce => 'H',
            sr => \N__18529\
        );

    \RSMRST_PWRGD.count_14_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20148\,
            in1 => \N__18635\,
            in2 => \_gnd_net_\,
            in3 => \N__16835\,
            lcout => \RSMRST_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_13\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14\,
            clk => \N__20631\,
            ce => 'H',
            sr => \N__18529\
        );

    \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18337\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_14\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_15_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18647\,
            in2 => \_gnd_net_\,
            in3 => \N__16832\,
            lcout => \RSMRST_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20637\,
            ce => \N__18497\,
            sr => \N__18522\
        );

    \VPP_VDDQ.count_0_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20128\,
            in1 => \N__18914\,
            in2 => \N__16894\,
            in3 => \N__16895\,
            lcout => \VPP_VDDQ.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_0\,
            clk => \N__20600\,
            ce => 'H',
            sr => \N__16942\
        );

    \VPP_VDDQ.count_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20110\,
            in1 => \N__18968\,
            in2 => \_gnd_net_\,
            in3 => \N__16877\,
            lcout => \VPP_VDDQ.countZ0Z_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_0\,
            carryout => \VPP_VDDQ.un1_count_1_cry_1\,
            clk => \N__20600\,
            ce => 'H',
            sr => \N__16942\
        );

    \VPP_VDDQ.count_2_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20129\,
            in1 => \N__18995\,
            in2 => \_gnd_net_\,
            in3 => \N__16874\,
            lcout => \VPP_VDDQ.countZ0Z_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_1_cry_2\,
            clk => \N__20600\,
            ce => 'H',
            sr => \N__16942\
        );

    \VPP_VDDQ.count_3_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20111\,
            in1 => \N__19070\,
            in2 => \_gnd_net_\,
            in3 => \N__16871\,
            lcout => \VPP_VDDQ.countZ0Z_3\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_1_cry_3\,
            clk => \N__20600\,
            ce => 'H',
            sr => \N__16942\
        );

    \VPP_VDDQ.count_4_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20130\,
            in1 => \N__19097\,
            in2 => \_gnd_net_\,
            in3 => \N__16868\,
            lcout => \VPP_VDDQ.countZ0Z_4\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_1_cry_4\,
            clk => \N__20600\,
            ce => 'H',
            sr => \N__16942\
        );

    \VPP_VDDQ.count_5_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20112\,
            in1 => \N__18470\,
            in2 => \_gnd_net_\,
            in3 => \N__16865\,
            lcout => \VPP_VDDQ.countZ0Z_5\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_1_cry_5\,
            clk => \N__20600\,
            ce => 'H',
            sr => \N__16942\
        );

    \VPP_VDDQ.count_6_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20131\,
            in1 => \N__19007\,
            in2 => \_gnd_net_\,
            in3 => \N__16862\,
            lcout => \VPP_VDDQ.countZ0Z_6\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_1_cry_6\,
            clk => \N__20600\,
            ce => 'H',
            sr => \N__16942\
        );

    \VPP_VDDQ.count_7_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20113\,
            in1 => \N__19084\,
            in2 => \_gnd_net_\,
            in3 => \N__16859\,
            lcout => \VPP_VDDQ.countZ0Z_7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_1_cry_7\,
            clk => \N__20600\,
            ce => 'H',
            sr => \N__16942\
        );

    \VPP_VDDQ.count_8_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20159\,
            in1 => \N__18941\,
            in2 => \_gnd_net_\,
            in3 => \N__16856\,
            lcout => \VPP_VDDQ.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_8\,
            clk => \N__20641\,
            ce => 'H',
            sr => \N__16930\
        );

    \VPP_VDDQ.count_9_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20155\,
            in1 => \N__18955\,
            in2 => \_gnd_net_\,
            in3 => \N__16976\,
            lcout => \VPP_VDDQ.countZ0Z_9\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_8\,
            carryout => \VPP_VDDQ.un1_count_1_cry_9\,
            clk => \N__20641\,
            ce => 'H',
            sr => \N__16930\
        );

    \VPP_VDDQ.count_10_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20156\,
            in1 => \N__18982\,
            in2 => \_gnd_net_\,
            in3 => \N__16973\,
            lcout => \VPP_VDDQ.countZ0Z_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_1_cry_10\,
            clk => \N__20641\,
            ce => 'H',
            sr => \N__16930\
        );

    \VPP_VDDQ.count_11_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20153\,
            in1 => \N__18928\,
            in2 => \_gnd_net_\,
            in3 => \N__16970\,
            lcout => \VPP_VDDQ.countZ0Z_11\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_1_cry_11\,
            clk => \N__20641\,
            ce => 'H',
            sr => \N__16930\
        );

    \VPP_VDDQ.count_12_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20157\,
            in1 => \N__19019\,
            in2 => \_gnd_net_\,
            in3 => \N__16967\,
            lcout => \VPP_VDDQ.countZ0Z_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_1_cry_12\,
            clk => \N__20641\,
            ce => 'H',
            sr => \N__16930\
        );

    \VPP_VDDQ.count_13_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20154\,
            in1 => \N__19033\,
            in2 => \_gnd_net_\,
            in3 => \N__16964\,
            lcout => \VPP_VDDQ.countZ0Z_13\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_1_cry_13\,
            clk => \N__20641\,
            ce => 'H',
            sr => \N__16930\
        );

    \VPP_VDDQ.count_14_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20158\,
            in1 => \N__19058\,
            in2 => \_gnd_net_\,
            in3 => \N__16961\,
            lcout => \VPP_VDDQ.countZ0Z_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14\,
            clk => \N__20641\,
            ce => 'H',
            sr => \N__16930\
        );

    \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18336\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_14\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_15_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19046\,
            in2 => \_gnd_net_\,
            in3 => \N__16958\,
            lcout => \VPP_VDDQ.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20642\,
            ce => \N__16955\,
            sr => \N__16946\
        );

    \COUNTER.counter_1_cry_1_c_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16910\,
            in2 => \N__17590\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_1_0_\,
            carryout => \COUNTER.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17552\,
            in2 => \_gnd_net_\,
            in3 => \N__17060\,
            lcout => \COUNTER.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_1\,
            carryout => \COUNTER.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17522\,
            in2 => \_gnd_net_\,
            in3 => \N__17057\,
            lcout => \COUNTER.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_2\,
            carryout => \COUNTER.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17612\,
            in2 => \_gnd_net_\,
            in3 => \N__17054\,
            lcout => \COUNTER.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_3\,
            carryout => \COUNTER.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17051\,
            in2 => \_gnd_net_\,
            in3 => \N__17030\,
            lcout => \COUNTER.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_4\,
            carryout => \COUNTER.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17026\,
            in2 => \_gnd_net_\,
            in3 => \N__17003\,
            lcout => \COUNTER.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_5\,
            carryout => \COUNTER.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_7_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16999\,
            in2 => \_gnd_net_\,
            in3 => \N__16985\,
            lcout => \COUNTER.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_6\,
            carryout => \COUNTER.counter_1_cry_7\,
            clk => \N__20407\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_8_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18670\,
            in2 => \_gnd_net_\,
            in3 => \N__16982\,
            lcout => \COUNTER.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_7\,
            carryout => \COUNTER.counter_1_cry_8\,
            clk => \N__20407\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_9_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18709\,
            in2 => \_gnd_net_\,
            in3 => \N__16979\,
            lcout => \COUNTER.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_2_0_\,
            carryout => \COUNTER.counter_1_cry_9\,
            clk => \N__20465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_10_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18727\,
            in2 => \_gnd_net_\,
            in3 => \N__17087\,
            lcout => \COUNTER.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_9\,
            carryout => \COUNTER.counter_1_cry_10\,
            clk => \N__20465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_11_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18688\,
            in2 => \_gnd_net_\,
            in3 => \N__17084\,
            lcout => \COUNTER.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_10\,
            carryout => \COUNTER.counter_1_cry_11\,
            clk => \N__20465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_12_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18811\,
            in2 => \_gnd_net_\,
            in3 => \N__17081\,
            lcout => \COUNTER.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_11\,
            carryout => \COUNTER.counter_1_cry_12\,
            clk => \N__20465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_13_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18844\,
            in2 => \_gnd_net_\,
            in3 => \N__17078\,
            lcout => \COUNTER.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_12\,
            carryout => \COUNTER.counter_1_cry_13\,
            clk => \N__20465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_14_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18859\,
            in2 => \_gnd_net_\,
            in3 => \N__17075\,
            lcout => \COUNTER.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_13\,
            carryout => \COUNTER.counter_1_cry_14\,
            clk => \N__20465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_15_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18826\,
            in2 => \_gnd_net_\,
            in3 => \N__17072\,
            lcout => \COUNTER.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_14\,
            carryout => \COUNTER.counter_1_cry_15\,
            clk => \N__20465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_16_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18745\,
            in2 => \_gnd_net_\,
            in3 => \N__17069\,
            lcout => \COUNTER.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_15\,
            carryout => \COUNTER.counter_1_cry_16\,
            clk => \N__20465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_17_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18781\,
            in2 => \_gnd_net_\,
            in3 => \N__17066\,
            lcout => \COUNTER.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_9_3_0_\,
            carryout => \COUNTER.counter_1_cry_17\,
            clk => \N__20408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_18_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18796\,
            in2 => \_gnd_net_\,
            in3 => \N__17063\,
            lcout => \COUNTER.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_17\,
            carryout => \COUNTER.counter_1_cry_18\,
            clk => \N__20408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_19_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18766\,
            in2 => \_gnd_net_\,
            in3 => \N__17114\,
            lcout => \COUNTER.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_18\,
            carryout => \COUNTER.counter_1_cry_19\,
            clk => \N__20408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_20_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17282\,
            in2 => \_gnd_net_\,
            in3 => \N__17111\,
            lcout => \COUNTER.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_19\,
            carryout => \COUNTER.counter_1_cry_20\,
            clk => \N__20408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_21_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17309\,
            in2 => \_gnd_net_\,
            in3 => \N__17108\,
            lcout => \COUNTER.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_20\,
            carryout => \COUNTER.counter_1_cry_21\,
            clk => \N__20408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_22_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17321\,
            in2 => \_gnd_net_\,
            in3 => \N__17105\,
            lcout => \COUNTER.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_21\,
            carryout => \COUNTER.counter_1_cry_22\,
            clk => \N__20408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_23_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17296\,
            in2 => \_gnd_net_\,
            in3 => \N__17102\,
            lcout => \COUNTER.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_22\,
            carryout => \COUNTER.counter_1_cry_23\,
            clk => \N__20408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_24_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17179\,
            in2 => \_gnd_net_\,
            in3 => \N__17099\,
            lcout => \COUNTER.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_23\,
            carryout => \COUNTER.counter_1_cry_24\,
            clk => \N__20408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_25_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17207\,
            in2 => \_gnd_net_\,
            in3 => \N__17096\,
            lcout => \COUNTER.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_9_4_0_\,
            carryout => \COUNTER.counter_1_cry_25\,
            clk => \N__20491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_26_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17219\,
            in2 => \_gnd_net_\,
            in3 => \N__17093\,
            lcout => \COUNTER.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_25\,
            carryout => \COUNTER.counter_1_cry_26\,
            clk => \N__20491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_27_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17194\,
            in2 => \_gnd_net_\,
            in3 => \N__17090\,
            lcout => \COUNTER.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_26\,
            carryout => \COUNTER.counter_1_cry_27\,
            clk => \N__20491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_28_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17153\,
            in2 => \_gnd_net_\,
            in3 => \N__17333\,
            lcout => \COUNTER.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_27\,
            carryout => \COUNTER.counter_1_cry_28\,
            clk => \N__20491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_29_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17140\,
            in2 => \_gnd_net_\,
            in3 => \N__17330\,
            lcout => \COUNTER.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_28\,
            carryout => \COUNTER.counter_1_cry_29\,
            clk => \N__20491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_30_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17165\,
            in2 => \_gnd_net_\,
            in3 => \N__17327\,
            lcout => \COUNTER.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_29\,
            carryout => \COUNTER.counter_1_cry_30\,
            clk => \N__20491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_31_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17126\,
            in2 => \_gnd_net_\,
            in3 => \N__17324\,
            lcout => \COUNTER.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_RNO_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17320\,
            in1 => \N__17308\,
            in2 => \N__17297\,
            in3 => \N__17281\,
            lcout => \COUNTER.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_RNI027U_11_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17269\,
            in1 => \N__17257\,
            in2 => \N__17246\,
            in3 => \N__17230\,
            lcout => \ALL_SYS_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_0_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__19435\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17577\,
            lcout => \COUNTER.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_RNO_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17218\,
            in1 => \N__17206\,
            in2 => \N__17195\,
            in3 => \N__17180\,
            lcout => \COUNTER.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNO_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17164\,
            in1 => \N__17152\,
            in2 => \N__17141\,
            in3 => \N__17125\,
            lcout => \COUNTER.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_4_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__17624\,
            in1 => \N__17607\,
            in2 => \_gnd_net_\,
            in3 => \N__19434\,
            lcout => \COUNTER.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_RNO_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17514\,
            in1 => \N__17544\,
            in2 => \N__17611\,
            in3 => \N__17576\,
            lcout => \COUNTER.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_2_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__17545\,
            in1 => \N__17561\,
            in2 => \_gnd_net_\,
            in3 => \N__19432\,
            lcout => \COUNTER.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_3_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19433\,
            in1 => \_gnd_net_\,
            in2 => \N__17521\,
            in3 => \N__17531\,
            lcout => \COUNTER.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17500\,
            in1 => \N__17488\,
            in2 => \N__17477\,
            in3 => \N__17461\,
            lcout => \ALL_SYS_PWRGD.un4_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17449\,
            in1 => \N__17437\,
            in2 => \N__17426\,
            in3 => \N__17410\,
            lcout => OPEN,
            ltout => \ALL_SYS_PWRGD.un4_count_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17399\,
            in1 => \N__17897\,
            in2 => \N__17393\,
            in3 => \N__17390\,
            lcout => \ALL_SYS_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_RNIV07U_10_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__17383\,
            in1 => \N__17371\,
            in2 => \N__17360\,
            in3 => \N__17344\,
            lcout => \ALL_SYS_PWRGD.un4_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_RNIKNST6_0_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19337\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20057\,
            lcout => \ALL_SYS_PWRGD.curr_state_RNIKNST6Z0Z_0\,
            ltout => \ALL_SYS_PWRGD.curr_state_RNIKNST6Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__20058\,
            in1 => \_gnd_net_\,
            in2 => \N__17861\,
            in3 => \_gnd_net_\,
            lcout => \ALL_SYS_PWRGD.N_65_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17841\,
            in1 => \N__17819\,
            in2 => \N__17804\,
            in3 => \N__17776\,
            lcout => rsmrst_pwrgd_signal,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__19431\,
            in1 => \_gnd_net_\,
            in2 => \N__17750\,
            in3 => \_gnd_net_\,
            lcout => \COUNTER.tmp_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_RNIRH3P_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17746\,
            in2 => \_gnd_net_\,
            in3 => \N__19430\,
            lcout => \tmp_RNIRH3P\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20092\,
            in1 => \N__17681\,
            in2 => \N__17702\,
            in3 => \N__17701\,
            lcout => \POWERLED.count_clkZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \POWERLED.un1_count_clk_1_cry_0\,
            clk => \N__20558\,
            ce => 'H',
            sr => \N__18251\
        );

    \POWERLED.count_clk_1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20085\,
            in1 => \N__17669\,
            in2 => \_gnd_net_\,
            in3 => \N__17651\,
            lcout => \POWERLED.count_clkZ0Z_1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_0\,
            carryout => \POWERLED.un1_count_clk_1_cry_1\,
            clk => \N__20558\,
            ce => 'H',
            sr => \N__18251\
        );

    \POWERLED.count_clk_2_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20093\,
            in1 => \N__17647\,
            in2 => \_gnd_net_\,
            in3 => \N__17627\,
            lcout => \POWERLED.count_clkZ0Z_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_1\,
            carryout => \POWERLED.un1_count_clk_1_cry_2\,
            clk => \N__20558\,
            ce => 'H',
            sr => \N__18251\
        );

    \POWERLED.count_clk_3_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20086\,
            in1 => \N__18116\,
            in2 => \_gnd_net_\,
            in3 => \N__18101\,
            lcout => \POWERLED.count_clkZ0Z_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_2\,
            carryout => \POWERLED.un1_count_clk_1_cry_3\,
            clk => \N__20558\,
            ce => 'H',
            sr => \N__18251\
        );

    \POWERLED.count_clk_4_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20094\,
            in1 => \N__18098\,
            in2 => \_gnd_net_\,
            in3 => \N__18083\,
            lcout => \POWERLED.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_3\,
            carryout => \POWERLED.un1_count_clk_1_cry_4\,
            clk => \N__20558\,
            ce => 'H',
            sr => \N__18251\
        );

    \POWERLED.count_clk_5_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20087\,
            in1 => \N__18080\,
            in2 => \_gnd_net_\,
            in3 => \N__18059\,
            lcout => \POWERLED.count_clkZ0Z_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_4\,
            carryout => \POWERLED.un1_count_clk_1_cry_5\,
            clk => \N__20558\,
            ce => 'H',
            sr => \N__18251\
        );

    \POWERLED.count_clk_6_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20095\,
            in1 => \N__18051\,
            in2 => \_gnd_net_\,
            in3 => \N__18023\,
            lcout => \POWERLED.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_5\,
            carryout => \POWERLED.un1_count_clk_1_cry_6\,
            clk => \N__20558\,
            ce => 'H',
            sr => \N__18251\
        );

    \POWERLED.count_clk_7_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20088\,
            in1 => \N__18000\,
            in2 => \_gnd_net_\,
            in3 => \N__17954\,
            lcout => \POWERLED.count_clkZ0Z_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_6\,
            carryout => \POWERLED.un1_count_clk_1_cry_7\,
            clk => \N__20558\,
            ce => 'H',
            sr => \N__18251\
        );

    \POWERLED.count_clk_8_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20099\,
            in1 => \N__17951\,
            in2 => \_gnd_net_\,
            in3 => \N__17936\,
            lcout => \POWERLED.count_clkZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \POWERLED.un1_count_clk_1_cry_8\,
            clk => \N__20543\,
            ce => 'H',
            sr => \N__18243\
        );

    \POWERLED.count_clk_9_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20091\,
            in1 => \N__17933\,
            in2 => \_gnd_net_\,
            in3 => \N__17915\,
            lcout => \POWERLED.count_clkZ0Z_9\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_8\,
            carryout => \POWERLED.un1_count_clk_1_cry_9\,
            clk => \N__20543\,
            ce => 'H',
            sr => \N__18243\
        );

    \POWERLED.count_clk_10_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20096\,
            in1 => \N__17912\,
            in2 => \_gnd_net_\,
            in3 => \N__17900\,
            lcout => \POWERLED.count_clkZ0Z_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_9\,
            carryout => \POWERLED.un1_count_clk_1_cry_10\,
            clk => \N__20543\,
            ce => 'H',
            sr => \N__18243\
        );

    \POWERLED.count_clk_11_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20089\,
            in1 => \N__18458\,
            in2 => \_gnd_net_\,
            in3 => \N__18446\,
            lcout => \POWERLED.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_10\,
            carryout => \POWERLED.un1_count_clk_1_cry_11\,
            clk => \N__20543\,
            ce => 'H',
            sr => \N__18243\
        );

    \POWERLED.count_clk_12_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20097\,
            in1 => \N__18443\,
            in2 => \_gnd_net_\,
            in3 => \N__18431\,
            lcout => \POWERLED.count_clkZ0Z_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_11\,
            carryout => \POWERLED.un1_count_clk_1_cry_12\,
            clk => \N__20543\,
            ce => 'H',
            sr => \N__18243\
        );

    \POWERLED.count_clk_13_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20090\,
            in1 => \N__18427\,
            in2 => \_gnd_net_\,
            in3 => \N__18413\,
            lcout => \POWERLED.count_clkZ0Z_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_12\,
            carryout => \POWERLED.un1_count_clk_1_cry_13\,
            clk => \N__20543\,
            ce => 'H',
            sr => \N__18243\
        );

    \POWERLED.count_clk_14_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20098\,
            in1 => \N__18410\,
            in2 => \_gnd_net_\,
            in3 => \N__18398\,
            lcout => \POWERLED.count_clkZ0Z_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_13\,
            carryout => \POWERLED.un1_count_clk_1_cry_14\,
            clk => \N__20543\,
            ce => 'H',
            sr => \N__18243\
        );

    \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18356\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_14\,
            carryout => \POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_esr_15_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18280\,
            in2 => \_gnd_net_\,
            in3 => \N__18284\,
            lcout => \POWERLED.count_clkZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20559\,
            ce => \N__18266\,
            sr => \N__18250\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_11_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18217\,
            in1 => \N__18205\,
            in2 => \N__18194\,
            in3 => \N__18178\,
            lcout => \RSMRST_PWRGD.m4_i_i_a2_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_9_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__18166\,
            in1 => \N__18154\,
            in2 => \N__18143\,
            in3 => \N__18127\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.m4_i_i_a2_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18656\,
            in1 => \N__18539\,
            in2 => \N__18650\,
            in3 => \N__18596\,
            lcout => \RSMRST_PWRGD.N_241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_7_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18646\,
            in2 => \_gnd_net_\,
            in3 => \N__18634\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.m4_i_i_a2_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_12_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18622\,
            in1 => \N__19229\,
            in2 => \N__18611\,
            in3 => \N__18607\,
            lcout => \RSMRST_PWRGD.m4_i_i_a2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_10_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18589\,
            in1 => \N__18577\,
            in2 => \N__18566\,
            in3 => \N__18550\,
            lcout => \RSMRST_PWRGD.m4_i_i_a2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__19524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19227\,
            lcout => \RSMRST_PWRGD.N_240\,
            ltout => \RSMRST_PWRGD.N_240_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNIJULM7_0_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__19186\,
            in1 => \N__20747\,
            in2 => \N__18533\,
            in3 => \N__20064\,
            lcout => \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0\,
            ltout => \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__20065\,
            in1 => \_gnd_net_\,
            in2 => \N__18500\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.N_65_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__19525\,
            in1 => \N__20746\,
            in2 => \_gnd_net_\,
            in3 => \N__19226\,
            lcout => \RSMRST_PWRGD.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIVJP51_3_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18469\,
            in1 => \N__19096\,
            in2 => \N__19085\,
            in3 => \N__19069\,
            lcout => \VPP_VDDQ.un6_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNI7CQO_15_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19057\,
            in1 => \N__19045\,
            in2 => \N__19034\,
            in3 => \N__19018\,
            lcout => \VPP_VDDQ.un6_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI63141_10_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19006\,
            in1 => \N__18994\,
            in2 => \N__18983\,
            in3 => \N__18967\,
            lcout => \VPP_VDDQ.un6_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFC141_11_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__18956\,
            in1 => \N__18940\,
            in2 => \N__18929\,
            in3 => \N__18913\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un6_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNIRFM64_15_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18902\,
            in1 => \N__18896\,
            in2 => \N__18890\,
            in3 => \N__18887\,
            lcout => \VPP_VDDQ.count_esr_RNIRFM64Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_RNO_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18860\,
            in1 => \N__18845\,
            in2 => \N__18830\,
            in3 => \N__18812\,
            lcout => \COUNTER.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_RNO_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18797\,
            in1 => \N__18782\,
            in2 => \N__18767\,
            in3 => \N__18749\,
            lcout => \COUNTER.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_RNO_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18731\,
            in1 => \N__18713\,
            in2 => \N__18695\,
            in3 => \N__18674\,
            lcout => \COUNTER.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19175\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => \COUNTER.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19166\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_0\,
            carryout => \COUNTER.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19154\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_1\,
            carryout => \COUNTER.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19145\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_2\,
            carryout => \COUNTER.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19136\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_3\,
            carryout => \COUNTER.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19127\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_4\,
            carryout => \COUNTER.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19115\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_5\,
            carryout => \COUNTER.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19106\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_6\,
            carryout => \COUNTER.un4_counter_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_THRU_LUT4_0_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19448\,
            lcout => \COUNTER.un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__19304\,
            in1 => \N__19470\,
            in2 => \_gnd_net_\,
            in3 => \N__19325\,
            lcout => OPEN,
            ltout => \ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_0_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__19328\,
            in1 => \N__19360\,
            in2 => \N__19388\,
            in3 => \N__19307\,
            lcout => \ALL_SYS_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20538\,
            ce => \N__19802\,
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_RNIUU4I2_0_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__19303\,
            in1 => \N__19471\,
            in2 => \_gnd_net_\,
            in3 => \N__19324\,
            lcout => \ALL_SYS_PWRGD.un1_curr_state10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_1_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101000100"
        )
    port map (
            in0 => \N__19327\,
            in1 => \N__19466\,
            in2 => \N__19361\,
            in3 => \N__19306\,
            lcout => \ALL_SYS_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20538\,
            ce => \N__19802\,
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_RNIP5P46_0_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__19302\,
            in1 => \N__19323\,
            in2 => \N__19472\,
            in3 => \N__19356\,
            lcout => \ALL_SYS_PWRGD.N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__19326\,
            in1 => \N__19465\,
            in2 => \_gnd_net_\,
            in3 => \N__19305\,
            lcout => vccst_pwrgd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20538\,
            ce => \N__19802\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_1_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__20743\,
            in1 => \N__19532\,
            in2 => \N__19228\,
            in3 => \N__19195\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20594\,
            ce => \N__19810\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_0_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20744\,
            in1 => \N__20764\,
            in2 => \_gnd_net_\,
            in3 => \N__19196\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20594\,
            ce => \N__19810\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20768\,
            in2 => \_gnd_net_\,
            in3 => \N__20745\,
            lcout => rsmrstn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20595\,
            ce => \N__19809\,
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_1_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19562\,
            in2 => \_gnd_net_\,
            in3 => \N__19538\,
            lcout => OPEN,
            ltout => \ALL_SYS_PWRGD.m4_0_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19523\,
            in1 => \N__19499\,
            in2 => \N__19487\,
            in3 => \N__19484\,
            lcout => \ALL_SYS_PWRGD.N_245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
