-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 13 2022 22:25:48

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : in std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : in std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : out std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : out std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__11747\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \VCCG0\ : std_logic;
signal v33a_enn : std_logic;
signal vpp_ok : std_logic;
signal vddq_en : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_12_1_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_1_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_1_0\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_5_1_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_5\ : std_logic;
signal \PCH_PWRGD.curr_state_e_0Z0Z_0\ : std_logic;
signal \PCH_PWRGD.m4_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.N_580_i_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_7_1_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_e_0Z0Z_1\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_15\ : std_logic;
signal \PCH_PWRGD.count_0_sqmuxa_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_0\ : std_logic;
signal \PCH_PWRGD.count_rst_14\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_13\ : std_logic;
signal \PCH_PWRGD.count_rst_13_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_1\ : std_logic;
signal \bfn_4_10_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_0\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_1\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_2\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_3\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_4\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_5\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_7\ : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_8\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_9\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_10\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_11\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_12\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_13\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal v5s_enn : std_logic;
signal slp_s4n : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_9\ : std_logic;
signal \PCH_PWRGD.count_rst_10_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_4\ : std_logic;
signal \PCH_PWRGD.count_0_5\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_1\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0\ : std_logic;
signal \bfn_5_6_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_5\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8\ : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_11\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_12\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_13\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_14\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_14_c_RNICCRZ0Z7\ : std_logic;
signal \PCH_PWRGD.count_RNI1N0D1Z0Z_10\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_10\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_14\ : std_logic;
signal vr_ready_vccin : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8PZ0Z7\ : std_logic;
signal \PCH_PWRGD.countZ0Z_13\ : std_logic;
signal \PCH_PWRGD.count_rst_1_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_13\ : std_logic;
signal slp_s3n : std_logic;
signal \PCH_PWRGD.count_rst_0\ : std_logic;
signal \PCH_PWRGD.count_rst_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_9_c_RNIEQ4KZ0Z5\ : std_logic;
signal \tmp_1_RNIBJDJ_cascade_\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_okZ0\ : std_logic;
signal \N_600_i\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_ok_e_1\ : std_logic;
signal \PCH_PWRGD.N_3_i\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_ok_e_1_cascade_\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_ok_0\ : std_logic;
signal v1p8a_ok : std_logic;
signal v5a_ok : std_logic;
signal v33a_ok : std_logic;
signal slp_susn : std_logic;
signal \PCH_PWRGD.count_m2_0_a2_0\ : std_logic;
signal \PCH_PWRGD.N_580_i\ : std_logic;
signal rsmrstn : std_logic;
signal \VPP_VDDQ.countZ0Z_3\ : std_logic;
signal \VPP_VDDQ.countZ0Z_5\ : std_logic;
signal \VPP_VDDQ.countZ0Z_7\ : std_logic;
signal \VPP_VDDQ.countZ0Z_4\ : std_logic;
signal \VPP_VDDQ.countZ0Z_6\ : std_logic;
signal \VPP_VDDQ.countZ0Z_2\ : std_logic;
signal \VPP_VDDQ.countZ0Z_10\ : std_logic;
signal \VPP_VDDQ.countZ0Z_1\ : std_logic;
signal \VPP_VDDQ.countZ0Z_14\ : std_logic;
signal \VPP_VDDQ.countZ0Z_12\ : std_logic;
signal \VPP_VDDQ.countZ0Z_13\ : std_logic;
signal \VPP_VDDQ.countZ0Z_15\ : std_logic;
signal \VPP_VDDQ.un6_count_11\ : std_logic;
signal \VPP_VDDQ.un6_count_8_cascade_\ : std_logic;
signal \VPP_VDDQ.un6_count_9\ : std_logic;
signal \VPP_VDDQ_un6_count_cascade_\ : std_logic;
signal \VPP_VDDQ_curr_state12\ : std_logic;
signal \VPP_VDDQ.countZ0Z_9\ : std_logic;
signal \VPP_VDDQ.countZ0Z_8\ : std_logic;
signal \VPP_VDDQ.countZ0Z_11\ : std_logic;
signal \VPP_VDDQ.countZ0Z_0\ : std_logic;
signal \VPP_VDDQ.un6_count_10\ : std_logic;
signal \VPP_VDDQ.un1_curr_state13_0\ : std_logic;
signal \VPP_VDDQ_un6_count\ : std_logic;
signal \VPP_VDDQ_delayed_vddq_pwrgd_1_sqmuxa\ : std_logic;
signal \VPP_VDDQ_delayed_vddq_pwrgd_1_sqmuxa_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state11\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\ : std_logic;
signal \G_24\ : std_logic;
signal \VPP_VDDQ.N_9_1\ : std_logic;
signal \VPP_VDDQ.curr_stateZ1Z_0\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_1\ : std_logic;
signal \VPP_VDDQ.un1_curr_state12_0\ : std_logic;
signal \VPP_VDDQ.un1_vddq_pwrgdZ0\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgdZ0\ : std_logic;
signal vccst_en : std_logic;
signal vpp_en : std_logic;
signal pch_pwrok : std_logic;
signal vccst_pwrgd : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_6\ : std_logic;
signal \PCH_PWRGD.count_rst_8\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_2\ : std_logic;
signal \PCH_PWRGD.count_rst_12\ : std_logic;
signal \PCH_PWRGD.countZ0Z_2\ : std_logic;
signal \PCH_PWRGD_N_3\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \PCH_PWRGD.count_rst_11\ : std_logic;
signal \PCH_PWRGD.curr_state_e_0_RNI4GQL2Z0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_3\ : std_logic;
signal \PCH_PWRGD.countZ0Z_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \PCH_PWRGD.countZ0Z_5\ : std_logic;
signal \PCH_PWRGD.count_rst_9\ : std_logic;
signal \PCH_PWRGD.count_rst_3_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_11\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10_c_RNI84NZ0Z7\ : std_logic;
signal \PCH_PWRGD.count_0_11\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \PCH_PWRGD.count_rst_7_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_7\ : std_logic;
signal \PCH_PWRGD.countZ0Z_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \PCH_PWRGD.count_rst_6_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_8\ : std_logic;
signal \PCH_PWRGD.countZ0Z_8\ : std_logic;
signal \PCH_PWRGD.count_rst_5_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9_cascade_\ : std_logic;
signal \PCH_PWRGD.N_1_i\ : std_logic;
signal \PCH_PWRGD.count_0_9\ : std_logic;
signal \PCH_PWRGD.count_rst_2\ : std_logic;
signal \PCH_PWRGD.count_rst_2_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_12\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_11_c_RNI96OZ0Z7\ : std_logic;
signal \PCH_PWRGD.countZ0Z_12\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal \COUNTER.un4_counter_0\ : std_logic;
signal \COUNTER.un4_counter_1\ : std_logic;
signal \COUNTER.un4_counter_2\ : std_logic;
signal \COUNTER.un4_counter_3\ : std_logic;
signal \COUNTER.un4_counter_4\ : std_logic;
signal \COUNTER.un4_counter_5\ : std_logic;
signal \COUNTER.un4_counter_6\ : std_logic;
signal \COUNTER_un4_counter_7\ : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \COUNTER_un4_counter_7_THRU_CO_cascade_\ : std_logic;
signal \COUNTER.un4_counter_0_and\ : std_logic;
signal \COUNTER.un4_counter_1_and\ : std_logic;
signal \COUNTER.un4_counter_2_and\ : std_logic;
signal \COUNTER.un4_counter_3_and\ : std_logic;
signal \COUNTER.un4_counter_4_and\ : std_logic;
signal \COUNTER.un4_counter_5_and\ : std_logic;
signal \COUNTER.un4_counter_7_and\ : std_logic;
signal \COUNTER.un4_counter_6_and\ : std_logic;
signal \RSMRST_PWRGD.curr_state10\ : std_logic;
signal \PCH_PWRGD.count_0_sqmuxa\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7\ : std_logic;
signal \PCH_PWRGD.countZ0Z_14\ : std_logic;
signal \PCH_PWRGD.count_rst_4\ : std_logic;
signal \PCH_PWRGD.countZ0Z_10\ : std_logic;
signal \PCH_PWRGD.curr_state_e_0_RNI4GQL2Z0Z_0\ : std_logic;
signal \PCH_PWRGD.count_m2_0_a2_iso\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_6_cascade_\ : std_logic;
signal \VPP_VDDQ.g0_3_a3_0_1\ : std_logic;
signal \VPP_VDDQ.N_6\ : std_logic;
signal \VPP_VDDQ.count_2_1_9_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_9_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_9\ : std_logic;
signal \VPP_VDDQ.count_2_1_5\ : std_logic;
signal \VPP_VDDQ.count_2_0_10\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_6\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_4\ : std_logic;
signal \VPP_VDDQ.count_2_1_6\ : std_logic;
signal \VPP_VDDQ.count_2_1_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_4\ : std_logic;
signal \VPP_VDDQ.count_2_RNI25V3Z0Z_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIZ0_cascade_\ : std_logic;
signal \VPP_VDDQ.m4_1_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2_e_0_RNINUSCZ0Z_1\ : std_logic;
signal \VPP_VDDQ.count_2_1_1\ : std_logic;
signal \COUNTER.counterZ0Z_1\ : std_logic;
signal \COUNTER.counterZ0Z_0\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \COUNTER.counterZ0Z_2\ : std_logic;
signal \COUNTER.counter_1_cry_1_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_1\ : std_logic;
signal \COUNTER.counterZ0Z_3\ : std_logic;
signal \COUNTER.counter_1_cry_2_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_2\ : std_logic;
signal \COUNTER.counterZ0Z_4\ : std_logic;
signal \COUNTER.counter_1_cry_3_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_3\ : std_logic;
signal \COUNTER.counterZ0Z_5\ : std_logic;
signal \COUNTER.counter_1_cry_4_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_4\ : std_logic;
signal \COUNTER.counterZ0Z_6\ : std_logic;
signal \COUNTER.counter_1_cry_5_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_5\ : std_logic;
signal \COUNTER.counterZ0Z_7\ : std_logic;
signal \COUNTER.counter_1_cry_6\ : std_logic;
signal \COUNTER.counterZ0Z_8\ : std_logic;
signal \COUNTER.counter_1_cry_7\ : std_logic;
signal \COUNTER.counter_1_cry_8\ : std_logic;
signal \COUNTER.counterZ0Z_9\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \COUNTER.counterZ0Z_10\ : std_logic;
signal \COUNTER.counter_1_cry_9\ : std_logic;
signal \COUNTER.counterZ0Z_11\ : std_logic;
signal \COUNTER.counter_1_cry_10\ : std_logic;
signal \COUNTER.counterZ0Z_12\ : std_logic;
signal \COUNTER.counter_1_cry_11\ : std_logic;
signal \COUNTER.counterZ0Z_13\ : std_logic;
signal \COUNTER.counter_1_cry_12\ : std_logic;
signal \COUNTER.counterZ0Z_14\ : std_logic;
signal \COUNTER.counter_1_cry_13\ : std_logic;
signal \COUNTER.counterZ0Z_15\ : std_logic;
signal \COUNTER.counter_1_cry_14\ : std_logic;
signal \COUNTER.counterZ0Z_16\ : std_logic;
signal \COUNTER.counter_1_cry_15\ : std_logic;
signal \COUNTER.counter_1_cry_16\ : std_logic;
signal \COUNTER.counterZ0Z_17\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \COUNTER.counterZ0Z_18\ : std_logic;
signal \COUNTER.counter_1_cry_17\ : std_logic;
signal \COUNTER.counterZ0Z_19\ : std_logic;
signal \COUNTER.counter_1_cry_18\ : std_logic;
signal \COUNTER.counterZ0Z_20\ : std_logic;
signal \COUNTER.counter_1_cry_19\ : std_logic;
signal \COUNTER.counterZ0Z_21\ : std_logic;
signal \COUNTER.counter_1_cry_20\ : std_logic;
signal \COUNTER.counterZ0Z_22\ : std_logic;
signal \COUNTER.counter_1_cry_21\ : std_logic;
signal \COUNTER.counterZ0Z_23\ : std_logic;
signal \COUNTER.counter_1_cry_22\ : std_logic;
signal \COUNTER.counterZ0Z_24\ : std_logic;
signal \COUNTER.counter_1_cry_23\ : std_logic;
signal \COUNTER.counter_1_cry_24\ : std_logic;
signal \COUNTER.counterZ0Z_25\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \COUNTER.counterZ0Z_26\ : std_logic;
signal \COUNTER.counter_1_cry_25\ : std_logic;
signal \COUNTER.counterZ0Z_27\ : std_logic;
signal \COUNTER.counter_1_cry_26\ : std_logic;
signal \COUNTER.counterZ0Z_28\ : std_logic;
signal \COUNTER.counter_1_cry_27\ : std_logic;
signal \COUNTER.counterZ0Z_29\ : std_logic;
signal \COUNTER.counter_1_cry_28\ : std_logic;
signal \COUNTER.counterZ0Z_30\ : std_logic;
signal \COUNTER.counter_1_cry_29\ : std_logic;
signal \COUNTER.counter_1_cry_30\ : std_logic;
signal \COUNTER.counterZ0Z_31\ : std_logic;
signal \RSMRST_PWRGD.un4_count_11\ : std_logic;
signal \RSMRST_PWRGD.un4_count_8_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_1_i_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_6_cascade_\ : std_logic;
signal \RSMRST_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\ : std_logic;
signal \G_10_cascade_\ : std_logic;
signal \RSMRST_PWRGD.un4_count_9\ : std_logic;
signal \RSMRST_PWRGD.N_3_i\ : std_logic;
signal \RSMRST_PWRGD.N_1_i\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.i3_mux_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \VPP_VDDQ_delayed_vddq_ok\ : std_logic;
signal \RSMRST_PWRGD.un4_count_10\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_okZ0\ : std_logic;
signal \VPP_VDDQ.count_2_1_3_cascade_\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1_cZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2_cZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_4\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIRZ0Z9731\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3_cZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4_cZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_6\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIVFZ0Z931\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5_cZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6_cZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7_cZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8_cZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8_cZ0_THRU_CO\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9_THRU_CO\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_RNOZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7_cZ0_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_0_8\ : std_logic;
signal \VPP_VDDQ.count_2_1_8_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_clk_100khz_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_1\ : std_logic;
signal \VPP_VDDQ.count_2_RNI82TR_0Z0Z_1\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_en\ : std_logic;
signal \VPP_VDDQ.count_2_en_0_tz_cascade_\ : std_logic;
signal \COUNTER_un4_counter_7_THRU_CO\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNIZ0Z_0_cascade_\ : std_logic;
signal \clk_100Khz_signalkeep\ : std_logic;
signal \VPP_VDDQ.m6_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_RNI_0Z0Z_2\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_4_1\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.count_2_0_0\ : std_logic;
signal \VPP_VDDQ.g0_0_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.g0_2_a2_1\ : std_logic;
signal \VPP_VDDQ.g0_2_a2_7\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.N_9_0\ : std_logic;
signal \VPP_VDDQ.N_10\ : std_logic;
signal \VPP_VDDQ.g0_2_a2_9_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_RNIUPFQ6Z0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.m4_0\ : std_logic;
signal \RSMRST_PWRGD.un1_curr_state10_0\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_2\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_3\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_4\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_5\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_7\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_9\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_11\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_12\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_13\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \tmp_1_RNIBJDJ_0\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \GNDG0\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_15\ : std_logic;
signal \RSMRST_PWRGD.N_9_2\ : std_logic;
signal \G_10\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_11_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_11\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6_c_RNI1JAZ0Z31\ : std_logic;
signal \VPP_VDDQ.count_2_1_7\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_7\ : std_logic;
signal \VPP_VDDQ.count_2_1_7_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_14_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_0_14\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_13_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_0_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_0_15\ : std_logic;
signal \VPP_VDDQ.count_2_1_15_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2_cZ0_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_0_3\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_10\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_9\ : std_logic;
signal \VPP_VDDQ.N_1_i_12_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_11\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_8\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_14_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_3\ : std_logic;
signal \VPP_VDDQ.count_2_RNIZ0Z_3\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1_cZ0_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2\ : std_logic;
signal \VPP_VDDQ.count_2_1_2\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_13\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_15\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_14\ : std_logic;
signal \VPP_VDDQ.g0_2_a2_8\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.count_2_RNIUPFQ6Z0Z_1\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_0\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1\ : std_logic;
signal vddq_ok : std_logic;
signal \VPP_VDDQ.curr_state_2_RNIZ0Z_0\ : std_logic;
signal \VPP_VDDQ.curr_state_2_e_0Z0Z_1\ : std_logic;
signal \tmp_1_RNIBJDJ\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4_cZ0_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_0_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11_THRU_CO\ : std_logic;
signal \VPP_VDDQ.m4_1\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_12\ : std_logic;
signal \VPP_VDDQ.un5_clk_100khz\ : std_logic;
signal \VPP_VDDQ.count_2_0_12\ : std_logic;
signal fpga_osc : std_logic;
signal \VPP_VDDQ.count_2_en\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \VCCST_OVERRIDE_3V3_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \SLP_S0n_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \PWRBTNn_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \GPIO_FPGA_SoC_2_wire\ : std_logic;
signal \VCCIN_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \CPU_C10_GATE_N_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \TPM_GPIO_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \PLTRSTn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \FPGA_OSC_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \SPI_FP_IO2_wire\ : std_logic;
signal \SATAXPCIE1_FPGA_wire\ : std_logic;
signal \GPIO_FPGA_EXP_1_wire\ : std_logic;
signal \VCCINAUX_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \GPIO_FPGA_EXP_2_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSACK_N_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \GPIO_FPGA_SoC_3_wire\ : std_logic;
signal \VR_PROCHOT_FPGA_OUT_N_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \SOC_SPKR_wire\ : std_logic;
signal \SLP_S5n_wire\ : std_logic;
signal \V12_MAIN_MON_wire\ : std_logic;
signal \SPI_FP_IO3_wire\ : std_logic;
signal \SATAXPCIE0_FPGA_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \FPGA_SLP_WLAN_N_wire\ : std_logic;

begin
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    V33A_ENn <= \V33A_ENn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \VCCST_OVERRIDE_3V3_wire\ <= VCCST_OVERRIDE_3V3;
    \V5S_OK_wire\ <= V5S_OK;
    \SLP_S3n_wire\ <= SLP_S3n;
    \SLP_S0n_wire\ <= SLP_S0n;
    V5S_ENn <= \V5S_ENn_wire\;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \PWRBTNn_wire\ <= PWRBTNn;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \GPIO_FPGA_SoC_2_wire\ <= GPIO_FPGA_SoC_2;
    \VCCIN_VR_PROCHOT_FPGA_wire\ <= VCCIN_VR_PROCHOT_FPGA;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    \CPU_C10_GATE_N_wire\ <= CPU_C10_GATE_N;
    VCCST_EN <= \VCCST_EN_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \TPM_GPIO_wire\ <= TPM_GPIO;
    \SUSWARN_N_wire\ <= SUSWARN_N;
    \PLTRSTn_wire\ <= PLTRSTn;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    \V5A_OK_wire\ <= V5A_OK;
    RSMRSTn <= \RSMRSTn_wire\;
    \FPGA_OSC_wire\ <= FPGA_OSC;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \SPI_FP_IO2_wire\ <= SPI_FP_IO2;
    \SATAXPCIE1_FPGA_wire\ <= SATAXPCIE1_FPGA;
    \GPIO_FPGA_EXP_1_wire\ <= GPIO_FPGA_EXP_1;
    \VCCINAUX_VR_PROCHOT_FPGA_wire\ <= VCCINAUX_VR_PROCHOT_FPGA;
    VCCINAUX_VR_PE <= \VCCINAUX_VR_PE_wire\;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    \GPIO_FPGA_EXP_2_wire\ <= GPIO_FPGA_EXP_2;
    VPP_EN <= \VPP_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    \SUSACK_N_wire\ <= SUSACK_N;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    DSW_PWROK <= \DSW_PWROK_wire\;
    V5A_EN <= \V5A_EN_wire\;
    \GPIO_FPGA_SoC_3_wire\ <= GPIO_FPGA_SoC_3;
    \VR_PROCHOT_FPGA_OUT_N_wire\ <= VR_PROCHOT_FPGA_OUT_N;
    \VPP_OK_wire\ <= VPP_OK;
    VCCIN_VR_PE <= \VCCIN_VR_PE_wire\;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \SOC_SPKR_wire\ <= SOC_SPKR;
    \SLP_S5n_wire\ <= SLP_S5n;
    \V12_MAIN_MON_wire\ <= V12_MAIN_MON;
    \SPI_FP_IO3_wire\ <= SPI_FP_IO3;
    \SATAXPCIE0_FPGA_wire\ <= SATAXPCIE0_FPGA;
    \V33A_OK_wire\ <= V33A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    \FPGA_SLP_WLAN_N_wire\ <= FPGA_SLP_WLAN_N;

    \ipInertedIOPad_VR_READY_VCCINAUX_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11747\,
            DIN => \N__11746\,
            DOUT => \N__11745\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \ipInertedIOPad_VR_READY_VCCINAUX_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11747\,
            PADOUT => \N__11746\,
            PADIN => \N__11745\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11738\,
            DIN => \N__11737\,
            DOUT => \N__11736\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \ipInertedIOPad_V33A_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11738\,
            PADOUT => \N__11737\,
            PADIN => \N__11736\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__4633\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11729\,
            DIN => \N__11728\,
            DOUT => \N__11727\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \ipInertedIOPad_V1P8A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11729\,
            PADOUT => \N__11728\,
            PADIN => \N__11727\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__5589\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11720\,
            DIN => \N__11719\,
            DOUT => \N__11718\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \ipInertedIOPad_VDDQ_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11720\,
            PADOUT => \N__11719\,
            PADIN => \N__11718\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__4615\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11711\,
            DIN => \N__11710\,
            DOUT => \N__11709\,
            PACKAGEPIN => \VCCST_OVERRIDE_3V3_wire\
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11711\,
            PADOUT => \N__11710\,
            PADIN => \N__11709\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11702\,
            DIN => \N__11701\,
            DOUT => \N__11700\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \ipInertedIOPad_V5S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11702\,
            PADOUT => \N__11701\,
            PADIN => \N__11700\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S3n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11693\,
            DIN => \N__11692\,
            DOUT => \N__11691\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \ipInertedIOPad_SLP_S3n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11693\,
            PADOUT => \N__11692\,
            PADIN => \N__11691\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s3n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S0n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11684\,
            DIN => \N__11683\,
            DOUT => \N__11682\,
            PACKAGEPIN => \SLP_S0n_wire\
        );

    \ipInertedIOPad_SLP_S0n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11684\,
            PADOUT => \N__11683\,
            PADIN => \N__11682\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11675\,
            DIN => \N__11674\,
            DOUT => \N__11673\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \ipInertedIOPad_V5S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11675\,
            PADOUT => \N__11674\,
            PADIN => \N__11673\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__4822\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11666\,
            DIN => \N__11665\,
            DOUT => \N__11664\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \ipInertedIOPad_V1P8A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11666\,
            PADOUT => \N__11665\,
            PADIN => \N__11664\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v1p8a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTNn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11657\,
            DIN => \N__11656\,
            DOUT => \N__11655\,
            PACKAGEPIN => \PWRBTNn_wire\
        );

    \ipInertedIOPad_PWRBTNn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11657\,
            PADOUT => \N__11656\,
            PADIN => \N__11655\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTN_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11648\,
            DIN => \N__11647\,
            DOUT => \N__11646\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \ipInertedIOPad_PWRBTN_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11648\,
            PADOUT => \N__11647\,
            PADIN => \N__11646\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11639\,
            DIN => \N__11638\,
            DOUT => \N__11637\,
            PACKAGEPIN => \GPIO_FPGA_SoC_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11639\,
            PADOUT => \N__11638\,
            PADIN => \N__11637\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11630\,
            DIN => \N__11629\,
            DOUT => \N__11628\,
            PACKAGEPIN => \VCCIN_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11630\,
            PADOUT => \N__11629\,
            PADIN => \N__11628\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_SUSn_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11621\,
            DIN => \N__11620\,
            DOUT => \N__11619\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \ipInertedIOPad_SLP_SUSn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11621\,
            PADOUT => \N__11620\,
            PADIN => \N__11619\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_susn,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CPU_C10_GATE_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11612\,
            DIN => \N__11611\,
            DOUT => \N__11610\,
            PACKAGEPIN => \CPU_C10_GATE_N_wire\
        );

    \ipInertedIOPad_CPU_C10_GATE_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11612\,
            PADOUT => \N__11611\,
            PADIN => \N__11610\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11603\,
            DIN => \N__11602\,
            DOUT => \N__11601\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \ipInertedIOPad_VCCST_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11603\,
            PADOUT => \N__11602\,
            PADIN => \N__11601\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__5977\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33DSW_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11594\,
            DIN => \N__11593\,
            DOUT => \N__11592\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \ipInertedIOPad_V33DSW_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11594\,
            PADOUT => \N__11593\,
            PADIN => \N__11592\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TPM_GPIO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11585\,
            DIN => \N__11584\,
            DOUT => \N__11583\,
            PACKAGEPIN => \TPM_GPIO_wire\
        );

    \ipInertedIOPad_TPM_GPIO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11585\,
            PADOUT => \N__11584\,
            PADIN => \N__11583\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSWARN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11576\,
            DIN => \N__11575\,
            DOUT => \N__11574\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \ipInertedIOPad_SUSWARN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11576\,
            PADOUT => \N__11575\,
            PADIN => \N__11574\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PLTRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11567\,
            DIN => \N__11566\,
            DOUT => \N__11565\,
            PACKAGEPIN => \PLTRSTn_wire\
        );

    \ipInertedIOPad_PLTRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11567\,
            PADOUT => \N__11566\,
            PADIN => \N__11565\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11558\,
            DIN => \N__11557\,
            DOUT => \N__11556\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11558\,
            PADOUT => \N__11557\,
            PADIN => \N__11556\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_READY_VCCIN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11549\,
            DIN => \N__11548\,
            DOUT => \N__11547\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \ipInertedIOPad_VR_READY_VCCIN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11549\,
            PADOUT => \N__11548\,
            PADIN => \N__11547\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccin,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11540\,
            DIN => \N__11539\,
            DOUT => \N__11538\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \ipInertedIOPad_V5A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11540\,
            PADOUT => \N__11539\,
            PADIN => \N__11538\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RSMRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11531\,
            DIN => \N__11530\,
            DOUT => \N__11529\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \ipInertedIOPad_RSMRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11531\,
            PADOUT => \N__11530\,
            PADIN => \N__11529\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__5476\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_OSC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11522\,
            DIN => \N__11521\,
            DOUT => \N__11520\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \ipInertedIOPad_FPGA_OSC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11522\,
            PADOUT => \N__11521\,
            PADIN => \N__11520\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => fpga_osc,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_PWRGD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11513\,
            DIN => \N__11512\,
            DOUT => \N__11511\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \ipInertedIOPad_VCCST_PWRGD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11513\,
            PADOUT => \N__11512\,
            PADIN => \N__11511\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__5875\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SYS_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11504\,
            DIN => \N__11503\,
            DOUT => \N__11502\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \ipInertedIOPad_SYS_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11504\,
            PADOUT => \N__11503\,
            PADIN => \N__11502\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__5919\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11495\,
            DIN => \N__11494\,
            DOUT => \N__11493\,
            PACKAGEPIN => \SPI_FP_IO2_wire\
        );

    \ipInertedIOPad_SPI_FP_IO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11495\,
            PADOUT => \N__11494\,
            PADIN => \N__11493\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11486\,
            DIN => \N__11485\,
            DOUT => \N__11484\,
            PACKAGEPIN => \SATAXPCIE1_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11486\,
            PADOUT => \N__11485\,
            PADIN => \N__11484\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11477\,
            DIN => \N__11476\,
            DOUT => \N__11475\,
            PACKAGEPIN => \GPIO_FPGA_EXP_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11477\,
            PADOUT => \N__11476\,
            PADIN => \N__11475\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11468\,
            DIN => \N__11467\,
            DOUT => \N__11466\,
            PACKAGEPIN => \VCCINAUX_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11468\,
            PADOUT => \N__11467\,
            PADIN => \N__11466\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11459\,
            DIN => \N__11458\,
            DOUT => \N__11457\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11459\,
            PADOUT => \N__11458\,
            PADIN => \N__11457\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__10105\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_HDA_SDO_ATP_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11450\,
            DIN => \N__11449\,
            DOUT => \N__11448\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \ipInertedIOPad_HDA_SDO_ATP_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11450\,
            PADOUT => \N__11449\,
            PADIN => \N__11448\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11441\,
            DIN => \N__11440\,
            DOUT => \N__11439\,
            PACKAGEPIN => \GPIO_FPGA_EXP_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11441\,
            PADOUT => \N__11440\,
            PADIN => \N__11439\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11432\,
            DIN => \N__11431\,
            DOUT => \N__11430\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \ipInertedIOPad_VPP_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11432\,
            PADOUT => \N__11431\,
            PADIN => \N__11430\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__5932\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11423\,
            DIN => \N__11422\,
            DOUT => \N__11421\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \ipInertedIOPad_VDDQ_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11423\,
            PADOUT => \N__11422\,
            PADIN => \N__11421\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vddq_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSACK_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11414\,
            DIN => \N__11413\,
            DOUT => \N__11412\,
            PACKAGEPIN => \SUSACK_N_wire\
        );

    \ipInertedIOPad_SUSACK_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11414\,
            PADOUT => \N__11413\,
            PADIN => \N__11412\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S4n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11405\,
            DIN => \N__11404\,
            DOUT => \N__11403\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \ipInertedIOPad_SLP_S4n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11405\,
            PADOUT => \N__11404\,
            PADIN => \N__11403\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s4n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_CPU_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11396\,
            DIN => \N__11395\,
            DOUT => \N__11394\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \ipInertedIOPad_VCCST_CPU_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11396\,
            PADOUT => \N__11395\,
            PADIN => \N__11394\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11387\,
            DIN => \N__11386\,
            DOUT => \N__11385\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \ipInertedIOPad_VCCINAUX_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11387\,
            PADOUT => \N__11386\,
            PADIN => \N__11385\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__5644\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11378\,
            DIN => \N__11377\,
            DOUT => \N__11376\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \ipInertedIOPad_V33S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11378\,
            PADOUT => \N__11377\,
            PADIN => \N__11376\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11369\,
            DIN => \N__11368\,
            DOUT => \N__11367\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \ipInertedIOPad_V33S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11369\,
            PADOUT => \N__11368\,
            PADIN => \N__11367\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__4818\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11360\,
            DIN => \N__11359\,
            DOUT => \N__11358\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11360\,
            PADOUT => \N__11359\,
            PADIN => \N__11358\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DSW_PWROK_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11351\,
            DIN => \N__11350\,
            DOUT => \N__11349\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \ipInertedIOPad_DSW_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11351\,
            PADOUT => \N__11350\,
            PADIN => \N__11349\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__10112\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11342\,
            DIN => \N__11341\,
            DOUT => \N__11340\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \ipInertedIOPad_V5A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11342\,
            PADOUT => \N__11341\,
            PADIN => \N__11340\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__5596\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11333\,
            DIN => \N__11332\,
            DOUT => \N__11331\,
            PACKAGEPIN => \GPIO_FPGA_SoC_3_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11333\,
            PADOUT => \N__11332\,
            PADIN => \N__11331\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11324\,
            DIN => \N__11323\,
            DOUT => \N__11322\,
            PACKAGEPIN => \VR_PROCHOT_FPGA_OUT_N_wire\
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11324\,
            PADOUT => \N__11323\,
            PADIN => \N__11322\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11315\,
            DIN => \N__11314\,
            DOUT => \N__11313\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \ipInertedIOPad_VPP_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11315\,
            PADOUT => \N__11314\,
            PADIN => \N__11313\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vpp_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11306\,
            DIN => \N__11305\,
            DOUT => \N__11304\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11306\,
            PADOUT => \N__11305\,
            PADIN => \N__11304\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11297\,
            DIN => \N__11296\,
            DOUT => \N__11295\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \ipInertedIOPad_VCCIN_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11297\,
            PADOUT => \N__11296\,
            PADIN => \N__11295\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SOC_SPKR_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11288\,
            DIN => \N__11287\,
            DOUT => \N__11286\,
            PACKAGEPIN => \SOC_SPKR_wire\
        );

    \ipInertedIOPad_SOC_SPKR_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11288\,
            PADOUT => \N__11287\,
            PADIN => \N__11286\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S5n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11279\,
            DIN => \N__11278\,
            DOUT => \N__11277\,
            PACKAGEPIN => \SLP_S5n_wire\
        );

    \ipInertedIOPad_SLP_S5n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11279\,
            PADOUT => \N__11278\,
            PADIN => \N__11277\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V12_MAIN_MON_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11270\,
            DIN => \N__11269\,
            DOUT => \N__11268\,
            PACKAGEPIN => \V12_MAIN_MON_wire\
        );

    \ipInertedIOPad_V12_MAIN_MON_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11270\,
            PADOUT => \N__11269\,
            PADIN => \N__11268\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11261\,
            DIN => \N__11260\,
            DOUT => \N__11259\,
            PACKAGEPIN => \SPI_FP_IO3_wire\
        );

    \ipInertedIOPad_SPI_FP_IO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11261\,
            PADOUT => \N__11260\,
            PADIN => \N__11259\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11252\,
            DIN => \N__11251\,
            DOUT => \N__11250\,
            PACKAGEPIN => \SATAXPCIE0_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11252\,
            PADOUT => \N__11251\,
            PADIN => \N__11250\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11243\,
            DIN => \N__11242\,
            DOUT => \N__11241\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \ipInertedIOPad_V33A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11243\,
            PADOUT => \N__11242\,
            PADIN => \N__11241\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PCH_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11234\,
            DIN => \N__11233\,
            DOUT => \N__11232\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \ipInertedIOPad_PCH_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11234\,
            PADOUT => \N__11233\,
            PADIN => \N__11232\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__5923\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11225\,
            DIN => \N__11224\,
            DOUT => \N__11223\,
            PACKAGEPIN => \FPGA_SLP_WLAN_N_wire\
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__11225\,
            PADOUT => \N__11224\,
            PADIN => \N__11223\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__2591\ : InMux
    port map (
            O => \N__11206\,
            I => \N__11202\
        );

    \I__2590\ : InMux
    port map (
            O => \N__11205\,
            I => \N__11198\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__11202\,
            I => \N__11194\
        );

    \I__2588\ : InMux
    port map (
            O => \N__11201\,
            I => \N__11190\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__11198\,
            I => \N__11187\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__11197\,
            I => \N__11184\
        );

    \I__2585\ : Span4Mux_v
    port map (
            O => \N__11194\,
            I => \N__11181\
        );

    \I__2584\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11178\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__11190\,
            I => \N__11175\
        );

    \I__2582\ : Span4Mux_v
    port map (
            O => \N__11187\,
            I => \N__11172\
        );

    \I__2581\ : InMux
    port map (
            O => \N__11184\,
            I => \N__11169\
        );

    \I__2580\ : Odrv4
    port map (
            O => \N__11181\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__11178\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__2578\ : Odrv12
    port map (
            O => \N__11175\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__11172\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__11169\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__2575\ : CascadeMux
    port map (
            O => \N__11158\,
            I => \N__11155\
        );

    \I__2574\ : InMux
    port map (
            O => \N__11155\,
            I => \N__11152\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__11152\,
            I => \N__11148\
        );

    \I__2572\ : InMux
    port map (
            O => \N__11151\,
            I => \N__11145\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__11148\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4_cZ0_THRU_CO\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__11145\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4_cZ0_THRU_CO\
        );

    \I__2569\ : InMux
    port map (
            O => \N__11140\,
            I => \N__11137\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__11137\,
            I => \N__11134\
        );

    \I__2567\ : Odrv12
    port map (
            O => \N__11134\,
            I => \VPP_VDDQ.count_2_0_5\
        );

    \I__2566\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11128\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__11128\,
            I => \N__11124\
        );

    \I__2564\ : InMux
    port map (
            O => \N__11127\,
            I => \N__11121\
        );

    \I__2563\ : Odrv4
    port map (
            O => \N__11124\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11_THRU_CO\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__11121\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11_THRU_CO\
        );

    \I__2561\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11110\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__11115\,
            I => \N__11102\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__11114\,
            I => \N__11095\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__11113\,
            I => \N__11089\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__11110\,
            I => \N__11085\
        );

    \I__2556\ : InMux
    port map (
            O => \N__11109\,
            I => \N__11080\
        );

    \I__2555\ : InMux
    port map (
            O => \N__11108\,
            I => \N__11075\
        );

    \I__2554\ : InMux
    port map (
            O => \N__11107\,
            I => \N__11068\
        );

    \I__2553\ : InMux
    port map (
            O => \N__11106\,
            I => \N__11068\
        );

    \I__2552\ : InMux
    port map (
            O => \N__11105\,
            I => \N__11068\
        );

    \I__2551\ : InMux
    port map (
            O => \N__11102\,
            I => \N__11061\
        );

    \I__2550\ : InMux
    port map (
            O => \N__11101\,
            I => \N__11061\
        );

    \I__2549\ : InMux
    port map (
            O => \N__11100\,
            I => \N__11061\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__11099\,
            I => \N__11056\
        );

    \I__2547\ : InMux
    port map (
            O => \N__11098\,
            I => \N__11048\
        );

    \I__2546\ : InMux
    port map (
            O => \N__11095\,
            I => \N__11035\
        );

    \I__2545\ : InMux
    port map (
            O => \N__11094\,
            I => \N__11035\
        );

    \I__2544\ : InMux
    port map (
            O => \N__11093\,
            I => \N__11035\
        );

    \I__2543\ : InMux
    port map (
            O => \N__11092\,
            I => \N__11035\
        );

    \I__2542\ : InMux
    port map (
            O => \N__11089\,
            I => \N__11035\
        );

    \I__2541\ : InMux
    port map (
            O => \N__11088\,
            I => \N__11035\
        );

    \I__2540\ : Span4Mux_v
    port map (
            O => \N__11085\,
            I => \N__11031\
        );

    \I__2539\ : CascadeMux
    port map (
            O => \N__11084\,
            I => \N__11027\
        );

    \I__2538\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11024\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__11080\,
            I => \N__11021\
        );

    \I__2536\ : InMux
    port map (
            O => \N__11079\,
            I => \N__11016\
        );

    \I__2535\ : InMux
    port map (
            O => \N__11078\,
            I => \N__11016\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__11075\,
            I => \N__11011\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__11068\,
            I => \N__11006\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__11061\,
            I => \N__11006\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__11060\,
            I => \N__11001\
        );

    \I__2530\ : CascadeMux
    port map (
            O => \N__11059\,
            I => \N__10998\
        );

    \I__2529\ : InMux
    port map (
            O => \N__11056\,
            I => \N__10991\
        );

    \I__2528\ : InMux
    port map (
            O => \N__11055\,
            I => \N__10991\
        );

    \I__2527\ : InMux
    port map (
            O => \N__11054\,
            I => \N__10991\
        );

    \I__2526\ : InMux
    port map (
            O => \N__11053\,
            I => \N__10988\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__11052\,
            I => \N__10985\
        );

    \I__2524\ : InMux
    port map (
            O => \N__11051\,
            I => \N__10982\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__11048\,
            I => \N__10977\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__11035\,
            I => \N__10977\
        );

    \I__2521\ : InMux
    port map (
            O => \N__11034\,
            I => \N__10974\
        );

    \I__2520\ : Sp12to4
    port map (
            O => \N__11031\,
            I => \N__10971\
        );

    \I__2519\ : InMux
    port map (
            O => \N__11030\,
            I => \N__10968\
        );

    \I__2518\ : InMux
    port map (
            O => \N__11027\,
            I => \N__10965\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__11024\,
            I => \N__10958\
        );

    \I__2516\ : Span4Mux_v
    port map (
            O => \N__11021\,
            I => \N__10958\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__11016\,
            I => \N__10958\
        );

    \I__2514\ : InMux
    port map (
            O => \N__11015\,
            I => \N__10955\
        );

    \I__2513\ : InMux
    port map (
            O => \N__11014\,
            I => \N__10952\
        );

    \I__2512\ : Span4Mux_h
    port map (
            O => \N__11011\,
            I => \N__10947\
        );

    \I__2511\ : Span4Mux_h
    port map (
            O => \N__11006\,
            I => \N__10947\
        );

    \I__2510\ : InMux
    port map (
            O => \N__11005\,
            I => \N__10938\
        );

    \I__2509\ : InMux
    port map (
            O => \N__11004\,
            I => \N__10938\
        );

    \I__2508\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10938\
        );

    \I__2507\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10938\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__10991\,
            I => \N__10935\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__10988\,
            I => \N__10932\
        );

    \I__2504\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10929\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10982\,
            I => \N__10922\
        );

    \I__2502\ : Span4Mux_h
    port map (
            O => \N__10977\,
            I => \N__10922\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__10974\,
            I => \N__10922\
        );

    \I__2500\ : Odrv12
    port map (
            O => \N__10971\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__10968\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__10965\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__2497\ : Odrv4
    port map (
            O => \N__10958\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__10955\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__10952\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__10947\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__10938\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__10935\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__2491\ : Odrv4
    port map (
            O => \N__10932\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10929\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__2489\ : Odrv4
    port map (
            O => \N__10922\,
            I => \VPP_VDDQ.m4_1\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__10897\,
            I => \N__10894\
        );

    \I__2487\ : InMux
    port map (
            O => \N__10894\,
            I => \N__10890\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__10893\,
            I => \N__10887\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__10890\,
            I => \N__10881\
        );

    \I__2484\ : InMux
    port map (
            O => \N__10887\,
            I => \N__10876\
        );

    \I__2483\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10876\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__10885\,
            I => \N__10873\
        );

    \I__2481\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10870\
        );

    \I__2480\ : Span4Mux_v
    port map (
            O => \N__10881\,
            I => \N__10867\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__10876\,
            I => \N__10864\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10873\,
            I => \N__10861\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__10870\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__2476\ : Odrv4
    port map (
            O => \N__10867\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__10864\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__10861\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__10852\,
            I => \N__10843\
        );

    \I__2472\ : InMux
    port map (
            O => \N__10851\,
            I => \N__10836\
        );

    \I__2471\ : InMux
    port map (
            O => \N__10850\,
            I => \N__10833\
        );

    \I__2470\ : InMux
    port map (
            O => \N__10849\,
            I => \N__10830\
        );

    \I__2469\ : CascadeMux
    port map (
            O => \N__10848\,
            I => \N__10824\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__10847\,
            I => \N__10820\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__10846\,
            I => \N__10814\
        );

    \I__2466\ : InMux
    port map (
            O => \N__10843\,
            I => \N__10800\
        );

    \I__2465\ : InMux
    port map (
            O => \N__10842\,
            I => \N__10800\
        );

    \I__2464\ : InMux
    port map (
            O => \N__10841\,
            I => \N__10800\
        );

    \I__2463\ : InMux
    port map (
            O => \N__10840\,
            I => \N__10797\
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__10839\,
            I => \N__10794\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__10836\,
            I => \N__10789\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__10833\,
            I => \N__10784\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__10830\,
            I => \N__10784\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__10829\,
            I => \N__10781\
        );

    \I__2457\ : InMux
    port map (
            O => \N__10828\,
            I => \N__10766\
        );

    \I__2456\ : InMux
    port map (
            O => \N__10827\,
            I => \N__10766\
        );

    \I__2455\ : InMux
    port map (
            O => \N__10824\,
            I => \N__10766\
        );

    \I__2454\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10766\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10820\,
            I => \N__10766\
        );

    \I__2452\ : InMux
    port map (
            O => \N__10819\,
            I => \N__10759\
        );

    \I__2451\ : InMux
    port map (
            O => \N__10818\,
            I => \N__10759\
        );

    \I__2450\ : InMux
    port map (
            O => \N__10817\,
            I => \N__10759\
        );

    \I__2449\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10756\
        );

    \I__2448\ : InMux
    port map (
            O => \N__10813\,
            I => \N__10749\
        );

    \I__2447\ : InMux
    port map (
            O => \N__10812\,
            I => \N__10749\
        );

    \I__2446\ : InMux
    port map (
            O => \N__10811\,
            I => \N__10749\
        );

    \I__2445\ : InMux
    port map (
            O => \N__10810\,
            I => \N__10740\
        );

    \I__2444\ : InMux
    port map (
            O => \N__10809\,
            I => \N__10740\
        );

    \I__2443\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10740\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10807\,
            I => \N__10740\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__10800\,
            I => \N__10737\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__10797\,
            I => \N__10734\
        );

    \I__2439\ : InMux
    port map (
            O => \N__10794\,
            I => \N__10731\
        );

    \I__2438\ : InMux
    port map (
            O => \N__10793\,
            I => \N__10721\
        );

    \I__2437\ : InMux
    port map (
            O => \N__10792\,
            I => \N__10721\
        );

    \I__2436\ : Span4Mux_v
    port map (
            O => \N__10789\,
            I => \N__10718\
        );

    \I__2435\ : Span4Mux_s3_h
    port map (
            O => \N__10784\,
            I => \N__10715\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10781\,
            I => \N__10712\
        );

    \I__2433\ : InMux
    port map (
            O => \N__10780\,
            I => \N__10703\
        );

    \I__2432\ : InMux
    port map (
            O => \N__10779\,
            I => \N__10703\
        );

    \I__2431\ : InMux
    port map (
            O => \N__10778\,
            I => \N__10703\
        );

    \I__2430\ : InMux
    port map (
            O => \N__10777\,
            I => \N__10703\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__10766\,
            I => \N__10698\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__10759\,
            I => \N__10698\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__10756\,
            I => \N__10691\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__10749\,
            I => \N__10691\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__10740\,
            I => \N__10691\
        );

    \I__2424\ : Span4Mux_v
    port map (
            O => \N__10737\,
            I => \N__10688\
        );

    \I__2423\ : Sp12to4
    port map (
            O => \N__10734\,
            I => \N__10683\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__10731\,
            I => \N__10683\
        );

    \I__2421\ : InMux
    port map (
            O => \N__10730\,
            I => \N__10678\
        );

    \I__2420\ : InMux
    port map (
            O => \N__10729\,
            I => \N__10678\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10728\,
            I => \N__10673\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10727\,
            I => \N__10673\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10726\,
            I => \N__10670\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__10721\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__2415\ : Odrv4
    port map (
            O => \N__10718\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__10715\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__10712\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__10703\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__2411\ : Odrv4
    port map (
            O => \N__10698\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__2410\ : Odrv4
    port map (
            O => \N__10691\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__2409\ : Odrv4
    port map (
            O => \N__10688\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__2408\ : Odrv12
    port map (
            O => \N__10683\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__10678\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__10673\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__10670\,
            I => \VPP_VDDQ.un5_clk_100khz\
        );

    \I__2404\ : InMux
    port map (
            O => \N__10645\,
            I => \N__10642\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__10642\,
            I => \N__10639\
        );

    \I__2402\ : Span4Mux_h
    port map (
            O => \N__10639\,
            I => \N__10636\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__10636\,
            I => \VPP_VDDQ.count_2_0_12\
        );

    \I__2400\ : ClkMux
    port map (
            O => \N__10633\,
            I => \N__10628\
        );

    \I__2399\ : ClkMux
    port map (
            O => \N__10632\,
            I => \N__10622\
        );

    \I__2398\ : ClkMux
    port map (
            O => \N__10631\,
            I => \N__10619\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__10628\,
            I => \N__10604\
        );

    \I__2396\ : ClkMux
    port map (
            O => \N__10627\,
            I => \N__10601\
        );

    \I__2395\ : ClkMux
    port map (
            O => \N__10626\,
            I => \N__10598\
        );

    \I__2394\ : ClkMux
    port map (
            O => \N__10625\,
            I => \N__10594\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__10622\,
            I => \N__10585\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__10619\,
            I => \N__10585\
        );

    \I__2391\ : ClkMux
    port map (
            O => \N__10618\,
            I => \N__10582\
        );

    \I__2390\ : ClkMux
    port map (
            O => \N__10617\,
            I => \N__10579\
        );

    \I__2389\ : ClkMux
    port map (
            O => \N__10616\,
            I => \N__10576\
        );

    \I__2388\ : ClkMux
    port map (
            O => \N__10615\,
            I => \N__10573\
        );

    \I__2387\ : ClkMux
    port map (
            O => \N__10614\,
            I => \N__10568\
        );

    \I__2386\ : ClkMux
    port map (
            O => \N__10613\,
            I => \N__10565\
        );

    \I__2385\ : ClkMux
    port map (
            O => \N__10612\,
            I => \N__10561\
        );

    \I__2384\ : ClkMux
    port map (
            O => \N__10611\,
            I => \N__10558\
        );

    \I__2383\ : ClkMux
    port map (
            O => \N__10610\,
            I => \N__10555\
        );

    \I__2382\ : ClkMux
    port map (
            O => \N__10609\,
            I => \N__10551\
        );

    \I__2381\ : ClkMux
    port map (
            O => \N__10608\,
            I => \N__10547\
        );

    \I__2380\ : ClkMux
    port map (
            O => \N__10607\,
            I => \N__10542\
        );

    \I__2379\ : Span4Mux_v
    port map (
            O => \N__10604\,
            I => \N__10534\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10601\,
            I => \N__10534\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__10598\,
            I => \N__10534\
        );

    \I__2376\ : ClkMux
    port map (
            O => \N__10597\,
            I => \N__10531\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__10594\,
            I => \N__10528\
        );

    \I__2374\ : ClkMux
    port map (
            O => \N__10593\,
            I => \N__10525\
        );

    \I__2373\ : ClkMux
    port map (
            O => \N__10592\,
            I => \N__10522\
        );

    \I__2372\ : ClkMux
    port map (
            O => \N__10591\,
            I => \N__10519\
        );

    \I__2371\ : ClkMux
    port map (
            O => \N__10590\,
            I => \N__10516\
        );

    \I__2370\ : Span4Mux_v
    port map (
            O => \N__10585\,
            I => \N__10511\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__10582\,
            I => \N__10511\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__10579\,
            I => \N__10506\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10576\,
            I => \N__10506\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__10573\,
            I => \N__10503\
        );

    \I__2365\ : ClkMux
    port map (
            O => \N__10572\,
            I => \N__10500\
        );

    \I__2364\ : ClkMux
    port map (
            O => \N__10571\,
            I => \N__10497\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__10568\,
            I => \N__10488\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10565\,
            I => \N__10488\
        );

    \I__2361\ : ClkMux
    port map (
            O => \N__10564\,
            I => \N__10485\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__10561\,
            I => \N__10482\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__10558\,
            I => \N__10477\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__10555\,
            I => \N__10477\
        );

    \I__2357\ : ClkMux
    port map (
            O => \N__10554\,
            I => \N__10474\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10551\,
            I => \N__10471\
        );

    \I__2355\ : ClkMux
    port map (
            O => \N__10550\,
            I => \N__10468\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__10547\,
            I => \N__10465\
        );

    \I__2353\ : ClkMux
    port map (
            O => \N__10546\,
            I => \N__10462\
        );

    \I__2352\ : ClkMux
    port map (
            O => \N__10545\,
            I => \N__10459\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__10542\,
            I => \N__10456\
        );

    \I__2350\ : ClkMux
    port map (
            O => \N__10541\,
            I => \N__10451\
        );

    \I__2349\ : Span4Mux_v
    port map (
            O => \N__10534\,
            I => \N__10445\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__10531\,
            I => \N__10445\
        );

    \I__2347\ : Span4Mux_v
    port map (
            O => \N__10528\,
            I => \N__10436\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10525\,
            I => \N__10436\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10522\,
            I => \N__10436\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__10519\,
            I => \N__10436\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__10516\,
            I => \N__10433\
        );

    \I__2342\ : Span4Mux_v
    port map (
            O => \N__10511\,
            I => \N__10430\
        );

    \I__2341\ : Span4Mux_v
    port map (
            O => \N__10506\,
            I => \N__10421\
        );

    \I__2340\ : Span4Mux_h
    port map (
            O => \N__10503\,
            I => \N__10421\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__10500\,
            I => \N__10421\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__10497\,
            I => \N__10421\
        );

    \I__2337\ : ClkMux
    port map (
            O => \N__10496\,
            I => \N__10418\
        );

    \I__2336\ : ClkMux
    port map (
            O => \N__10495\,
            I => \N__10415\
        );

    \I__2335\ : ClkMux
    port map (
            O => \N__10494\,
            I => \N__10412\
        );

    \I__2334\ : ClkMux
    port map (
            O => \N__10493\,
            I => \N__10408\
        );

    \I__2333\ : Span4Mux_v
    port map (
            O => \N__10488\,
            I => \N__10402\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__10485\,
            I => \N__10402\
        );

    \I__2331\ : Span4Mux_h
    port map (
            O => \N__10482\,
            I => \N__10395\
        );

    \I__2330\ : Span4Mux_v
    port map (
            O => \N__10477\,
            I => \N__10395\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10474\,
            I => \N__10395\
        );

    \I__2328\ : Span4Mux_h
    port map (
            O => \N__10471\,
            I => \N__10390\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__10468\,
            I => \N__10390\
        );

    \I__2326\ : Span4Mux_v
    port map (
            O => \N__10465\,
            I => \N__10385\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__10462\,
            I => \N__10385\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__10459\,
            I => \N__10380\
        );

    \I__2323\ : Span4Mux_h
    port map (
            O => \N__10456\,
            I => \N__10380\
        );

    \I__2322\ : ClkMux
    port map (
            O => \N__10455\,
            I => \N__10377\
        );

    \I__2321\ : ClkMux
    port map (
            O => \N__10454\,
            I => \N__10374\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__10451\,
            I => \N__10371\
        );

    \I__2319\ : ClkMux
    port map (
            O => \N__10450\,
            I => \N__10368\
        );

    \I__2318\ : Span4Mux_v
    port map (
            O => \N__10445\,
            I => \N__10365\
        );

    \I__2317\ : Span4Mux_v
    port map (
            O => \N__10436\,
            I => \N__10362\
        );

    \I__2316\ : Span4Mux_v
    port map (
            O => \N__10433\,
            I => \N__10349\
        );

    \I__2315\ : Span4Mux_h
    port map (
            O => \N__10430\,
            I => \N__10349\
        );

    \I__2314\ : Span4Mux_v
    port map (
            O => \N__10421\,
            I => \N__10349\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__10418\,
            I => \N__10349\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__10415\,
            I => \N__10349\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__10412\,
            I => \N__10349\
        );

    \I__2310\ : ClkMux
    port map (
            O => \N__10411\,
            I => \N__10346\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__10408\,
            I => \N__10343\
        );

    \I__2308\ : ClkMux
    port map (
            O => \N__10407\,
            I => \N__10340\
        );

    \I__2307\ : Span4Mux_v
    port map (
            O => \N__10402\,
            I => \N__10337\
        );

    \I__2306\ : Span4Mux_v
    port map (
            O => \N__10395\,
            I => \N__10326\
        );

    \I__2305\ : Span4Mux_v
    port map (
            O => \N__10390\,
            I => \N__10326\
        );

    \I__2304\ : Span4Mux_h
    port map (
            O => \N__10385\,
            I => \N__10326\
        );

    \I__2303\ : Span4Mux_v
    port map (
            O => \N__10380\,
            I => \N__10326\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__10377\,
            I => \N__10326\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__10374\,
            I => \N__10323\
        );

    \I__2300\ : Span4Mux_h
    port map (
            O => \N__10371\,
            I => \N__10318\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__10368\,
            I => \N__10318\
        );

    \I__2298\ : IoSpan4Mux
    port map (
            O => \N__10365\,
            I => \N__10309\
        );

    \I__2297\ : Span4Mux_h
    port map (
            O => \N__10362\,
            I => \N__10309\
        );

    \I__2296\ : Span4Mux_v
    port map (
            O => \N__10349\,
            I => \N__10309\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__10346\,
            I => \N__10309\
        );

    \I__2294\ : Span12Mux_s5_h
    port map (
            O => \N__10343\,
            I => \N__10304\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__10340\,
            I => \N__10304\
        );

    \I__2292\ : Span4Mux_v
    port map (
            O => \N__10337\,
            I => \N__10299\
        );

    \I__2291\ : Span4Mux_v
    port map (
            O => \N__10326\,
            I => \N__10299\
        );

    \I__2290\ : Span4Mux_v
    port map (
            O => \N__10323\,
            I => \N__10294\
        );

    \I__2289\ : Span4Mux_v
    port map (
            O => \N__10318\,
            I => \N__10294\
        );

    \I__2288\ : IoSpan4Mux
    port map (
            O => \N__10309\,
            I => \N__10291\
        );

    \I__2287\ : Odrv12
    port map (
            O => \N__10304\,
            I => fpga_osc
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__10299\,
            I => fpga_osc
        );

    \I__2285\ : Odrv4
    port map (
            O => \N__10294\,
            I => fpga_osc
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__10291\,
            I => fpga_osc
        );

    \I__2283\ : CEMux
    port map (
            O => \N__10282\,
            I => \N__10264\
        );

    \I__2282\ : CEMux
    port map (
            O => \N__10281\,
            I => \N__10261\
        );

    \I__2281\ : CEMux
    port map (
            O => \N__10280\,
            I => \N__10257\
        );

    \I__2280\ : CEMux
    port map (
            O => \N__10279\,
            I => \N__10254\
        );

    \I__2279\ : CEMux
    port map (
            O => \N__10278\,
            I => \N__10251\
        );

    \I__2278\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10244\
        );

    \I__2277\ : InMux
    port map (
            O => \N__10276\,
            I => \N__10244\
        );

    \I__2276\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10244\
        );

    \I__2275\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10235\
        );

    \I__2274\ : InMux
    port map (
            O => \N__10273\,
            I => \N__10235\
        );

    \I__2273\ : InMux
    port map (
            O => \N__10272\,
            I => \N__10235\
        );

    \I__2272\ : InMux
    port map (
            O => \N__10271\,
            I => \N__10235\
        );

    \I__2271\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10232\
        );

    \I__2270\ : CEMux
    port map (
            O => \N__10269\,
            I => \N__10227\
        );

    \I__2269\ : CEMux
    port map (
            O => \N__10268\,
            I => \N__10224\
        );

    \I__2268\ : CEMux
    port map (
            O => \N__10267\,
            I => \N__10221\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__10264\,
            I => \N__10216\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__10261\,
            I => \N__10216\
        );

    \I__2265\ : CEMux
    port map (
            O => \N__10260\,
            I => \N__10213\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__10257\,
            I => \N__10208\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__10254\,
            I => \N__10208\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__10251\,
            I => \N__10201\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__10244\,
            I => \N__10198\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__10235\,
            I => \N__10193\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__10232\,
            I => \N__10193\
        );

    \I__2258\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10188\
        );

    \I__2257\ : InMux
    port map (
            O => \N__10230\,
            I => \N__10188\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__10227\,
            I => \N__10182\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__10224\,
            I => \N__10179\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__10221\,
            I => \N__10176\
        );

    \I__2253\ : Span4Mux_h
    port map (
            O => \N__10216\,
            I => \N__10171\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__10213\,
            I => \N__10171\
        );

    \I__2251\ : Span4Mux_s3_h
    port map (
            O => \N__10208\,
            I => \N__10168\
        );

    \I__2250\ : InMux
    port map (
            O => \N__10207\,
            I => \N__10163\
        );

    \I__2249\ : InMux
    port map (
            O => \N__10206\,
            I => \N__10163\
        );

    \I__2248\ : InMux
    port map (
            O => \N__10205\,
            I => \N__10160\
        );

    \I__2247\ : InMux
    port map (
            O => \N__10204\,
            I => \N__10157\
        );

    \I__2246\ : Span4Mux_h
    port map (
            O => \N__10201\,
            I => \N__10152\
        );

    \I__2245\ : Span4Mux_s3_h
    port map (
            O => \N__10198\,
            I => \N__10152\
        );

    \I__2244\ : Span4Mux_v
    port map (
            O => \N__10193\,
            I => \N__10147\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__10188\,
            I => \N__10147\
        );

    \I__2242\ : InMux
    port map (
            O => \N__10187\,
            I => \N__10144\
        );

    \I__2241\ : InMux
    port map (
            O => \N__10186\,
            I => \N__10139\
        );

    \I__2240\ : InMux
    port map (
            O => \N__10185\,
            I => \N__10139\
        );

    \I__2239\ : Odrv12
    port map (
            O => \N__10182\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__10179\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__2237\ : Odrv4
    port map (
            O => \N__10176\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__2236\ : Odrv4
    port map (
            O => \N__10171\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__10168\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__10163\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__10160\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__10157\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__10152\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__10147\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__10144\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__10139\,
            I => \VPP_VDDQ.count_2_en\
        );

    \I__2227\ : InMux
    port map (
            O => \N__10114\,
            I => \N__10109\
        );

    \I__2226\ : InMux
    port map (
            O => \N__10113\,
            I => \N__10106\
        );

    \I__2225\ : IoInMux
    port map (
            O => \N__10112\,
            I => \N__10102\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__10109\,
            I => \N__10099\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__10106\,
            I => \N__10096\
        );

    \I__2222\ : IoInMux
    port map (
            O => \N__10105\,
            I => \N__10093\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__10102\,
            I => \N__10090\
        );

    \I__2220\ : Span4Mux_v
    port map (
            O => \N__10099\,
            I => \N__10087\
        );

    \I__2219\ : Span4Mux_h
    port map (
            O => \N__10096\,
            I => \N__10084\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__10093\,
            I => \N__10081\
        );

    \I__2217\ : Span12Mux_s8_h
    port map (
            O => \N__10090\,
            I => \N__10078\
        );

    \I__2216\ : Span4Mux_h
    port map (
            O => \N__10087\,
            I => \N__10075\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__10084\,
            I => \N__10070\
        );

    \I__2214\ : IoSpan4Mux
    port map (
            O => \N__10081\,
            I => \N__10070\
        );

    \I__2213\ : Odrv12
    port map (
            O => \N__10078\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__10075\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__10070\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__10063\,
            I => \N__10060\
        );

    \I__2209\ : InMux
    port map (
            O => \N__10060\,
            I => \N__10057\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__10057\,
            I => \N__10054\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__10054\,
            I => \N__10050\
        );

    \I__2206\ : InMux
    port map (
            O => \N__10053\,
            I => \N__10047\
        );

    \I__2205\ : Odrv4
    port map (
            O => \N__10050\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_cZ0_THRU_CO\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__10047\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_cZ0_THRU_CO\
        );

    \I__2203\ : InMux
    port map (
            O => \N__10042\,
            I => \N__10039\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__10039\,
            I => \N__10036\
        );

    \I__2201\ : Span4Mux_h
    port map (
            O => \N__10036\,
            I => \N__10033\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__10033\,
            I => \VPP_VDDQ.count_2_0_3\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__10030\,
            I => \N__10026\
        );

    \I__2198\ : InMux
    port map (
            O => \N__10029\,
            I => \N__10023\
        );

    \I__2197\ : InMux
    port map (
            O => \N__10026\,
            I => \N__10019\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__10023\,
            I => \N__10015\
        );

    \I__2195\ : CascadeMux
    port map (
            O => \N__10022\,
            I => \N__10012\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__10019\,
            I => \N__10008\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__10018\,
            I => \N__10005\
        );

    \I__2192\ : Span4Mux_v
    port map (
            O => \N__10015\,
            I => \N__10002\
        );

    \I__2191\ : InMux
    port map (
            O => \N__10012\,
            I => \N__9999\
        );

    \I__2190\ : InMux
    port map (
            O => \N__10011\,
            I => \N__9996\
        );

    \I__2189\ : Span4Mux_v
    port map (
            O => \N__10008\,
            I => \N__9993\
        );

    \I__2188\ : InMux
    port map (
            O => \N__10005\,
            I => \N__9990\
        );

    \I__2187\ : Odrv4
    port map (
            O => \N__10002\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9999\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__9996\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__9993\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__9990\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9979\,
            I => \N__9976\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9976\,
            I => \N__9971\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9975\,
            I => \N__9968\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9974\,
            I => \N__9965\
        );

    \I__2178\ : Span4Mux_h
    port map (
            O => \N__9971\,
            I => \N__9957\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__9968\,
            I => \N__9957\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9965\,
            I => \N__9957\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9954\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__9957\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__9954\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__2172\ : CascadeMux
    port map (
            O => \N__9949\,
            I => \VPP_VDDQ.N_1_i_12_cascade_\
        );

    \I__2171\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9941\
        );

    \I__2170\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9938\
        );

    \I__2169\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9934\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__9941\,
            I => \N__9929\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9938\,
            I => \N__9929\
        );

    \I__2166\ : CascadeMux
    port map (
            O => \N__9937\,
            I => \N__9926\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9934\,
            I => \N__9923\
        );

    \I__2164\ : Span4Mux_v
    port map (
            O => \N__9929\,
            I => \N__9920\
        );

    \I__2163\ : InMux
    port map (
            O => \N__9926\,
            I => \N__9917\
        );

    \I__2162\ : Odrv12
    port map (
            O => \N__9923\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__9920\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__9917\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__9910\,
            I => \N__9906\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__9909\,
            I => \N__9902\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9906\,
            I => \N__9897\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9905\,
            I => \N__9894\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9902\,
            I => \N__9891\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9901\,
            I => \N__9888\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9900\,
            I => \N__9885\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__9897\,
            I => \N__9882\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__9894\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__9891\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__9888\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9885\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__9882\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__9871\,
            I => \VPP_VDDQ.un9_clk_100khz_14_1_cascade_\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9868\,
            I => \N__9865\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__9865\,
            I => \N__9858\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9864\,
            I => \N__9855\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9863\,
            I => \N__9852\
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__9862\,
            I => \N__9849\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9861\,
            I => \N__9846\
        );

    \I__2139\ : Span4Mux_v
    port map (
            O => \N__9858\,
            I => \N__9841\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9855\,
            I => \N__9841\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9852\,
            I => \N__9838\
        );

    \I__2136\ : InMux
    port map (
            O => \N__9849\,
            I => \N__9835\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__9846\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__2134\ : Odrv4
    port map (
            O => \N__9841\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__2133\ : Odrv12
    port map (
            O => \N__9838\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9835\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__2131\ : InMux
    port map (
            O => \N__9826\,
            I => \N__9823\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__9823\,
            I => \VPP_VDDQ.count_2_RNIZ0Z_3\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9820\,
            I => \N__9817\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__9817\,
            I => \N__9813\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9816\,
            I => \N__9810\
        );

    \I__2126\ : Span4Mux_v
    port map (
            O => \N__9813\,
            I => \N__9805\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__9810\,
            I => \N__9805\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__9805\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1_cZ0_THRU_CO\
        );

    \I__2123\ : CascadeMux
    port map (
            O => \N__9802\,
            I => \N__9798\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9801\,
            I => \N__9795\
        );

    \I__2121\ : InMux
    port map (
            O => \N__9798\,
            I => \N__9790\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9795\,
            I => \N__9787\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9794\,
            I => \N__9782\
        );

    \I__2118\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9782\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9790\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__9787\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9782\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__9775\,
            I => \N__9772\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9772\,
            I => \N__9769\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__9769\,
            I => \VPP_VDDQ.count_2_1_2\
        );

    \I__2111\ : InMux
    port map (
            O => \N__9766\,
            I => \N__9758\
        );

    \I__2110\ : InMux
    port map (
            O => \N__9765\,
            I => \N__9758\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__9764\,
            I => \N__9755\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9763\,
            I => \N__9752\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__9758\,
            I => \N__9749\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9746\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__9752\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__9749\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__9746\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__9739\,
            I => \N__9733\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9738\,
            I => \N__9730\
        );

    \I__2100\ : InMux
    port map (
            O => \N__9737\,
            I => \N__9727\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9736\,
            I => \N__9722\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9733\,
            I => \N__9722\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__9730\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__9727\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__9722\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9715\,
            I => \N__9707\
        );

    \I__2093\ : InMux
    port map (
            O => \N__9714\,
            I => \N__9707\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__9713\,
            I => \N__9704\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9712\,
            I => \N__9701\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9707\,
            I => \N__9698\
        );

    \I__2089\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9695\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__9701\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__9698\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9695\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__2085\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9685\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__9685\,
            I => \VPP_VDDQ.g0_2_a2_8\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9682\,
            I => \N__9678\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9681\,
            I => \N__9675\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__9678\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9675\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__2079\ : InMux
    port map (
            O => \N__9670\,
            I => \N__9667\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__9667\,
            I => \VPP_VDDQ.count_2_RNIUPFQ6Z0Z_1\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9664\,
            I => \N__9661\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9661\,
            I => \VPP_VDDQ.curr_state_2_0_0\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9658\,
            I => \N__9653\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__9657\,
            I => \N__9649\
        );

    \I__2073\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9645\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__9653\,
            I => \N__9642\
        );

    \I__2071\ : InMux
    port map (
            O => \N__9652\,
            I => \N__9638\
        );

    \I__2070\ : InMux
    port map (
            O => \N__9649\,
            I => \N__9635\
        );

    \I__2069\ : InMux
    port map (
            O => \N__9648\,
            I => \N__9632\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__9645\,
            I => \N__9627\
        );

    \I__2067\ : Span4Mux_h
    port map (
            O => \N__9642\,
            I => \N__9627\
        );

    \I__2066\ : InMux
    port map (
            O => \N__9641\,
            I => \N__9624\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9638\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__9635\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__9632\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__9627\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__9624\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__9613\,
            I => \N__9609\
        );

    \I__2059\ : InMux
    port map (
            O => \N__9612\,
            I => \N__9603\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9609\,
            I => \N__9598\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9608\,
            I => \N__9595\
        );

    \I__2056\ : CascadeMux
    port map (
            O => \N__9607\,
            I => \N__9591\
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__9606\,
            I => \N__9588\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__9603\,
            I => \N__9584\
        );

    \I__2053\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9581\
        );

    \I__2052\ : InMux
    port map (
            O => \N__9601\,
            I => \N__9577\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__9598\,
            I => \N__9574\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__9595\,
            I => \N__9570\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9594\,
            I => \N__9561\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9591\,
            I => \N__9561\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9561\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9561\
        );

    \I__2045\ : Span4Mux_v
    port map (
            O => \N__9584\,
            I => \N__9556\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__9581\,
            I => \N__9556\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9580\,
            I => \N__9553\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9577\,
            I => \N__9548\
        );

    \I__2041\ : Span4Mux_h
    port map (
            O => \N__9574\,
            I => \N__9545\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9573\,
            I => \N__9542\
        );

    \I__2039\ : Span4Mux_v
    port map (
            O => \N__9570\,
            I => \N__9537\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__9561\,
            I => \N__9537\
        );

    \I__2037\ : Span4Mux_v
    port map (
            O => \N__9556\,
            I => \N__9532\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9553\,
            I => \N__9532\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9552\,
            I => \N__9527\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9551\,
            I => \N__9527\
        );

    \I__2033\ : Span4Mux_v
    port map (
            O => \N__9548\,
            I => \N__9520\
        );

    \I__2032\ : Span4Mux_s3_h
    port map (
            O => \N__9545\,
            I => \N__9520\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9542\,
            I => \N__9520\
        );

    \I__2030\ : Span4Mux_v
    port map (
            O => \N__9537\,
            I => \N__9513\
        );

    \I__2029\ : Span4Mux_h
    port map (
            O => \N__9532\,
            I => \N__9513\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9527\,
            I => \N__9513\
        );

    \I__2027\ : Span4Mux_v
    port map (
            O => \N__9520\,
            I => \N__9510\
        );

    \I__2026\ : IoSpan4Mux
    port map (
            O => \N__9513\,
            I => \N__9507\
        );

    \I__2025\ : Odrv4
    port map (
            O => \N__9510\,
            I => vddq_ok
        );

    \I__2024\ : Odrv4
    port map (
            O => \N__9507\,
            I => vddq_ok
        );

    \I__2023\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9497\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__9501\,
            I => \N__9494\
        );

    \I__2021\ : CascadeMux
    port map (
            O => \N__9500\,
            I => \N__9491\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__9497\,
            I => \N__9488\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9481\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9491\,
            I => \N__9478\
        );

    \I__2017\ : Span4Mux_h
    port map (
            O => \N__9488\,
            I => \N__9475\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9468\
        );

    \I__2015\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9468\
        );

    \I__2014\ : InMux
    port map (
            O => \N__9485\,
            I => \N__9468\
        );

    \I__2013\ : InMux
    port map (
            O => \N__9484\,
            I => \N__9465\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__9481\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_0\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__9478\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_0\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__9475\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_0\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__9468\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_0\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__9465\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_0\
        );

    \I__2007\ : InMux
    port map (
            O => \N__9454\,
            I => \N__9451\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__9451\,
            I => \VPP_VDDQ.curr_state_2_e_0Z0Z_1\
        );

    \I__2005\ : CEMux
    port map (
            O => \N__9448\,
            I => \N__9441\
        );

    \I__2004\ : CEMux
    port map (
            O => \N__9447\,
            I => \N__9438\
        );

    \I__2003\ : CEMux
    port map (
            O => \N__9446\,
            I => \N__9435\
        );

    \I__2002\ : InMux
    port map (
            O => \N__9445\,
            I => \N__9432\
        );

    \I__2001\ : InMux
    port map (
            O => \N__9444\,
            I => \N__9429\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9441\,
            I => \N__9426\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__9438\,
            I => \N__9423\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__9435\,
            I => \N__9420\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__9432\,
            I => \N__9416\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__9429\,
            I => \N__9413\
        );

    \I__1995\ : Span12Mux_s7_v
    port map (
            O => \N__9426\,
            I => \N__9410\
        );

    \I__1994\ : Sp12to4
    port map (
            O => \N__9423\,
            I => \N__9405\
        );

    \I__1993\ : Sp12to4
    port map (
            O => \N__9420\,
            I => \N__9405\
        );

    \I__1992\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9402\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__9416\,
            I => \N__9399\
        );

    \I__1990\ : Span4Mux_h
    port map (
            O => \N__9413\,
            I => \N__9396\
        );

    \I__1989\ : Odrv12
    port map (
            O => \N__9410\,
            I => \tmp_1_RNIBJDJ\
        );

    \I__1988\ : Odrv12
    port map (
            O => \N__9405\,
            I => \tmp_1_RNIBJDJ\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__9402\,
            I => \tmp_1_RNIBJDJ\
        );

    \I__1986\ : Odrv4
    port map (
            O => \N__9399\,
            I => \tmp_1_RNIBJDJ\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__9396\,
            I => \tmp_1_RNIBJDJ\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__9385\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0_cascade_\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__9382\,
            I => \VPP_VDDQ.count_2Z0Z_14_cascade_\
        );

    \I__1982\ : InMux
    port map (
            O => \N__9379\,
            I => \N__9373\
        );

    \I__1981\ : InMux
    port map (
            O => \N__9378\,
            I => \N__9373\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__9373\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13_THRU_CO\
        );

    \I__1979\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9367\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__9367\,
            I => \VPP_VDDQ.count_2_0_14\
        );

    \I__1977\ : CascadeMux
    port map (
            O => \N__9364\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0_cascade_\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__9361\,
            I => \VPP_VDDQ.count_2Z0Z_13_cascade_\
        );

    \I__1975\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9352\
        );

    \I__1974\ : InMux
    port map (
            O => \N__9357\,
            I => \N__9352\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__9352\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12_THRU_CO\
        );

    \I__1972\ : InMux
    port map (
            O => \N__9349\,
            I => \N__9346\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__9346\,
            I => \VPP_VDDQ.count_2_0_13\
        );

    \I__1970\ : InMux
    port map (
            O => \N__9343\,
            I => \N__9339\
        );

    \I__1969\ : InMux
    port map (
            O => \N__9342\,
            I => \N__9336\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__9339\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_THRU_CO\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__9336\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_THRU_CO\
        );

    \I__1966\ : InMux
    port map (
            O => \N__9331\,
            I => \N__9328\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__9328\,
            I => \VPP_VDDQ.count_2_0_15\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__9325\,
            I => \VPP_VDDQ.count_2_1_15_cascade_\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__9322\,
            I => \VPP_VDDQ.count_2Z0Z_2_cascade_\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9319\,
            I => \N__9316\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__9316\,
            I => \VPP_VDDQ.count_2_0_2\
        );

    \I__1960\ : SRMux
    port map (
            O => \N__9313\,
            I => \N__9310\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__9310\,
            I => \N__9306\
        );

    \I__1958\ : SRMux
    port map (
            O => \N__9309\,
            I => \N__9303\
        );

    \I__1957\ : Span4Mux_v
    port map (
            O => \N__9306\,
            I => \N__9298\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__9303\,
            I => \N__9298\
        );

    \I__1955\ : Span4Mux_v
    port map (
            O => \N__9298\,
            I => \N__9294\
        );

    \I__1954\ : SRMux
    port map (
            O => \N__9297\,
            I => \N__9291\
        );

    \I__1953\ : Sp12to4
    port map (
            O => \N__9294\,
            I => \N__9286\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__9291\,
            I => \N__9286\
        );

    \I__1951\ : Odrv12
    port map (
            O => \N__9286\,
            I => \G_10\
        );

    \I__1950\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9280\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__9280\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\
        );

    \I__1948\ : InMux
    port map (
            O => \N__9277\,
            I => \N__9273\
        );

    \I__1947\ : InMux
    port map (
            O => \N__9276\,
            I => \N__9270\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__9273\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10_THRU_CO\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__9270\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10_THRU_CO\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__9265\,
            I => \VPP_VDDQ.count_2Z0Z_11_cascade_\
        );

    \I__1943\ : InMux
    port map (
            O => \N__9262\,
            I => \N__9259\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__9259\,
            I => \VPP_VDDQ.count_2_0_11\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9256\,
            I => \N__9251\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9255\,
            I => \N__9246\
        );

    \I__1939\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9246\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__9251\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNI1JAZ0Z31\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__9246\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNI1JAZ0Z31\
        );

    \I__1936\ : InMux
    port map (
            O => \N__9241\,
            I => \N__9238\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__9238\,
            I => \N__9235\
        );

    \I__1934\ : Span4Mux_h
    port map (
            O => \N__9235\,
            I => \N__9232\
        );

    \I__1933\ : Odrv4
    port map (
            O => \N__9232\,
            I => \VPP_VDDQ.count_2_1_7\
        );

    \I__1932\ : InMux
    port map (
            O => \N__9229\,
            I => \N__9225\
        );

    \I__1931\ : InMux
    port map (
            O => \N__9228\,
            I => \N__9222\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__9225\,
            I => \N__9216\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__9222\,
            I => \N__9216\
        );

    \I__1928\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9213\
        );

    \I__1927\ : Span4Mux_v
    port map (
            O => \N__9216\,
            I => \N__9210\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__9213\,
            I => \VPP_VDDQ.count_2Z0Z_7\
        );

    \I__1925\ : Odrv4
    port map (
            O => \N__9210\,
            I => \VPP_VDDQ.count_2Z0Z_7\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__9205\,
            I => \VPP_VDDQ.count_2_1_7_cascade_\
        );

    \I__1923\ : InMux
    port map (
            O => \N__9202\,
            I => \N__9199\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__9199\,
            I => \VPP_VDDQ.un1_count_2_1_axb_7\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__9196\,
            I => \N__9193\
        );

    \I__1920\ : InMux
    port map (
            O => \N__9193\,
            I => \N__9190\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__9190\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\
        );

    \I__1918\ : CascadeMux
    port map (
            O => \N__9187\,
            I => \N__9184\
        );

    \I__1917\ : InMux
    port map (
            O => \N__9184\,
            I => \N__9180\
        );

    \I__1916\ : InMux
    port map (
            O => \N__9183\,
            I => \N__9177\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__9180\,
            I => \N__9174\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__9177\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__1913\ : Odrv4
    port map (
            O => \N__9174\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__1912\ : InMux
    port map (
            O => \N__9169\,
            I => \RSMRST_PWRGD.un1_count_1_cry_8\
        );

    \I__1911\ : InMux
    port map (
            O => \N__9166\,
            I => \N__9162\
        );

    \I__1910\ : InMux
    port map (
            O => \N__9165\,
            I => \N__9159\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__9162\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__9159\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__1907\ : InMux
    port map (
            O => \N__9154\,
            I => \RSMRST_PWRGD.un1_count_1_cry_9\
        );

    \I__1906\ : InMux
    port map (
            O => \N__9151\,
            I => \N__9147\
        );

    \I__1905\ : InMux
    port map (
            O => \N__9150\,
            I => \N__9144\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__9147\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__9144\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__1902\ : InMux
    port map (
            O => \N__9139\,
            I => \RSMRST_PWRGD.un1_count_1_cry_10\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__9136\,
            I => \N__9132\
        );

    \I__1900\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9129\
        );

    \I__1899\ : InMux
    port map (
            O => \N__9132\,
            I => \N__9126\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__9129\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__9126\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__1896\ : InMux
    port map (
            O => \N__9121\,
            I => \RSMRST_PWRGD.un1_count_1_cry_11\
        );

    \I__1895\ : InMux
    port map (
            O => \N__9118\,
            I => \N__9114\
        );

    \I__1894\ : InMux
    port map (
            O => \N__9117\,
            I => \N__9111\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__9114\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__9111\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1891\ : InMux
    port map (
            O => \N__9106\,
            I => \RSMRST_PWRGD.un1_count_1_cry_12\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__9103\,
            I => \N__9091\
        );

    \I__1889\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9081\
        );

    \I__1888\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9065\
        );

    \I__1887\ : InMux
    port map (
            O => \N__9100\,
            I => \N__9065\
        );

    \I__1886\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9065\
        );

    \I__1885\ : InMux
    port map (
            O => \N__9098\,
            I => \N__9065\
        );

    \I__1884\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9056\
        );

    \I__1883\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9056\
        );

    \I__1882\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9056\
        );

    \I__1881\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9056\
        );

    \I__1880\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9050\
        );

    \I__1879\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9041\
        );

    \I__1878\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9041\
        );

    \I__1877\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9041\
        );

    \I__1876\ : InMux
    port map (
            O => \N__9087\,
            I => \N__9041\
        );

    \I__1875\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9034\
        );

    \I__1874\ : InMux
    port map (
            O => \N__9085\,
            I => \N__9034\
        );

    \I__1873\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9034\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__9081\,
            I => \N__9022\
        );

    \I__1871\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9010\
        );

    \I__1870\ : InMux
    port map (
            O => \N__9079\,
            I => \N__9010\
        );

    \I__1869\ : InMux
    port map (
            O => \N__9078\,
            I => \N__9010\
        );

    \I__1868\ : InMux
    port map (
            O => \N__9077\,
            I => \N__9010\
        );

    \I__1867\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9003\
        );

    \I__1866\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9003\
        );

    \I__1865\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9003\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__9065\,
            I => \N__9000\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__9056\,
            I => \N__8997\
        );

    \I__1862\ : InMux
    port map (
            O => \N__9055\,
            I => \N__8990\
        );

    \I__1861\ : InMux
    port map (
            O => \N__9054\,
            I => \N__8990\
        );

    \I__1860\ : InMux
    port map (
            O => \N__9053\,
            I => \N__8990\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__9050\,
            I => \N__8987\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__9041\,
            I => \N__8982\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__9034\,
            I => \N__8982\
        );

    \I__1856\ : InMux
    port map (
            O => \N__9033\,
            I => \N__8979\
        );

    \I__1855\ : InMux
    port map (
            O => \N__9032\,
            I => \N__8970\
        );

    \I__1854\ : InMux
    port map (
            O => \N__9031\,
            I => \N__8970\
        );

    \I__1853\ : InMux
    port map (
            O => \N__9030\,
            I => \N__8970\
        );

    \I__1852\ : InMux
    port map (
            O => \N__9029\,
            I => \N__8970\
        );

    \I__1851\ : InMux
    port map (
            O => \N__9028\,
            I => \N__8961\
        );

    \I__1850\ : InMux
    port map (
            O => \N__9027\,
            I => \N__8961\
        );

    \I__1849\ : InMux
    port map (
            O => \N__9026\,
            I => \N__8961\
        );

    \I__1848\ : InMux
    port map (
            O => \N__9025\,
            I => \N__8961\
        );

    \I__1847\ : Span4Mux_h
    port map (
            O => \N__9022\,
            I => \N__8958\
        );

    \I__1846\ : InMux
    port map (
            O => \N__9021\,
            I => \N__8951\
        );

    \I__1845\ : InMux
    port map (
            O => \N__9020\,
            I => \N__8951\
        );

    \I__1844\ : InMux
    port map (
            O => \N__9019\,
            I => \N__8951\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__9010\,
            I => \N__8938\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__9003\,
            I => \N__8938\
        );

    \I__1841\ : Span4Mux_v
    port map (
            O => \N__9000\,
            I => \N__8938\
        );

    \I__1840\ : Span4Mux_v
    port map (
            O => \N__8997\,
            I => \N__8938\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8990\,
            I => \N__8938\
        );

    \I__1838\ : Span4Mux_v
    port map (
            O => \N__8987\,
            I => \N__8931\
        );

    \I__1837\ : Span4Mux_h
    port map (
            O => \N__8982\,
            I => \N__8931\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__8979\,
            I => \N__8931\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8970\,
            I => \N__8926\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__8961\,
            I => \N__8926\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__8958\,
            I => \N__8921\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8951\,
            I => \N__8921\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8950\,
            I => \N__8916\
        );

    \I__1830\ : InMux
    port map (
            O => \N__8949\,
            I => \N__8916\
        );

    \I__1829\ : Span4Mux_h
    port map (
            O => \N__8938\,
            I => \N__8913\
        );

    \I__1828\ : Odrv4
    port map (
            O => \N__8931\,
            I => \tmp_1_RNIBJDJ_0\
        );

    \I__1827\ : Odrv4
    port map (
            O => \N__8926\,
            I => \tmp_1_RNIBJDJ_0\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__8921\,
            I => \tmp_1_RNIBJDJ_0\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__8916\,
            I => \tmp_1_RNIBJDJ_0\
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__8913\,
            I => \tmp_1_RNIBJDJ_0\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8902\,
            I => \N__8898\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8901\,
            I => \N__8895\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8898\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8895\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8890\,
            I => \RSMRST_PWRGD.un1_count_1_cry_13\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8887\,
            I => \bfn_9_7_0_\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__8884\,
            I => \N__8880\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8883\,
            I => \N__8877\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8880\,
            I => \N__8874\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8877\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8874\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__1812\ : CEMux
    port map (
            O => \N__8869\,
            I => \N__8866\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8866\,
            I => \RSMRST_PWRGD.N_9_2\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8863\,
            I => \N__8859\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8862\,
            I => \N__8856\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8859\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8856\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8851\,
            I => \RSMRST_PWRGD.un1_count_1_cry_0\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8848\,
            I => \N__8844\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8841\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8844\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8841\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8836\,
            I => \RSMRST_PWRGD.un1_count_1_cry_1\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8833\,
            I => \N__8829\
        );

    \I__1799\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8826\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8829\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8826\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8821\,
            I => \RSMRST_PWRGD.un1_count_1_cry_2\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8818\,
            I => \N__8814\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8817\,
            I => \N__8811\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8814\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__8811\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8806\,
            I => \RSMRST_PWRGD.un1_count_1_cry_3\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8803\,
            I => \N__8799\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8802\,
            I => \N__8796\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8799\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__8796\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8791\,
            I => \RSMRST_PWRGD.un1_count_1_cry_4\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8788\,
            I => \N__8784\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8787\,
            I => \N__8781\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8784\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8781\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__1781\ : InMux
    port map (
            O => \N__8776\,
            I => \RSMRST_PWRGD.un1_count_1_cry_5\
        );

    \I__1780\ : CascadeMux
    port map (
            O => \N__8773\,
            I => \N__8769\
        );

    \I__1779\ : InMux
    port map (
            O => \N__8772\,
            I => \N__8766\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8763\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__8766\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__8763\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8758\,
            I => \RSMRST_PWRGD.un1_count_1_cry_6\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8755\,
            I => \N__8751\
        );

    \I__1773\ : InMux
    port map (
            O => \N__8754\,
            I => \N__8748\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8751\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__8748\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8743\,
            I => \bfn_9_6_0_\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8740\,
            I => \N__8737\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8737\,
            I => \N__8734\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__8734\,
            I => \VPP_VDDQ.un9_clk_100khz_4_1\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__8731\,
            I => \N__8728\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8728\,
            I => \N__8725\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8725\,
            I => \N__8722\
        );

    \I__1763\ : Span4Mux_h
    port map (
            O => \N__8722\,
            I => \N__8717\
        );

    \I__1762\ : InMux
    port map (
            O => \N__8721\,
            I => \N__8712\
        );

    \I__1761\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8712\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__8717\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__8712\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8707\,
            I => \N__8704\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__8704\,
            I => \VPP_VDDQ.count_2_0_0\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__8701\,
            I => \VPP_VDDQ.g0_0_0_cascade_\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8698\,
            I => \N__8691\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8688\
        );

    \I__1753\ : InMux
    port map (
            O => \N__8696\,
            I => \N__8685\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8695\,
            I => \N__8680\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8680\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__8691\,
            I => \N__8677\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__8688\,
            I => \N__8674\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8685\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8680\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__1746\ : Odrv12
    port map (
            O => \N__8677\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__8674\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8665\,
            I => \N__8662\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8662\,
            I => \VPP_VDDQ.g0_2_a2_1\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8659\,
            I => \N__8656\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__8656\,
            I => \VPP_VDDQ.g0_2_a2_7\
        );

    \I__1740\ : CascadeMux
    port map (
            O => \N__8653\,
            I => \VPP_VDDQ.count_2Z0Z_0_cascade_\
        );

    \I__1739\ : InMux
    port map (
            O => \N__8650\,
            I => \N__8647\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8647\,
            I => \N__8644\
        );

    \I__1737\ : Odrv4
    port map (
            O => \N__8644\,
            I => \VPP_VDDQ.N_9_0\
        );

    \I__1736\ : InMux
    port map (
            O => \N__8641\,
            I => \N__8638\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8638\,
            I => \N__8635\
        );

    \I__1734\ : Span4Mux_v
    port map (
            O => \N__8635\,
            I => \N__8632\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__8632\,
            I => \VPP_VDDQ.N_10\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__8629\,
            I => \VPP_VDDQ.g0_2_a2_9_cascade_\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__8626\,
            I => \VPP_VDDQ.count_2_RNIUPFQ6Z0Z_1_cascade_\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8623\,
            I => \N__8620\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8620\,
            I => \VPP_VDDQ.m4_0\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__8617\,
            I => \N__8613\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8610\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8613\,
            I => \N__8607\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8610\,
            I => \RSMRST_PWRGD.un1_curr_state10_0\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8607\,
            I => \RSMRST_PWRGD.un1_curr_state10_0\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8602\,
            I => \N__8598\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8601\,
            I => \N__8595\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__8598\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8595\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__8590\,
            I => \VPP_VDDQ.count_2_en_0_tz_cascade_\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8587\,
            I => \N__8582\
        );

    \I__1717\ : InMux
    port map (
            O => \N__8586\,
            I => \N__8574\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8571\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8582\,
            I => \N__8563\
        );

    \I__1714\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8560\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8580\,
            I => \N__8551\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8551\
        );

    \I__1711\ : InMux
    port map (
            O => \N__8578\,
            I => \N__8551\
        );

    \I__1710\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8551\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__8574\,
            I => \N__8548\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__8571\,
            I => \N__8545\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8538\
        );

    \I__1706\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8538\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8538\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8567\,
            I => \N__8535\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8566\,
            I => \N__8532\
        );

    \I__1702\ : Span4Mux_v
    port map (
            O => \N__8563\,
            I => \N__8527\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8560\,
            I => \N__8527\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8551\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__8548\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__8545\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__8538\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__8535\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8532\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__8527\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__8512\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__8509\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_0_cascade_\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__8506\,
            I => \N__8499\
        );

    \I__1690\ : InMux
    port map (
            O => \N__8505\,
            I => \N__8490\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8504\,
            I => \N__8490\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__8503\,
            I => \N__8487\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8502\,
            I => \N__8482\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8499\,
            I => \N__8482\
        );

    \I__1685\ : InMux
    port map (
            O => \N__8498\,
            I => \N__8475\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8497\,
            I => \N__8475\
        );

    \I__1683\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8469\
        );

    \I__1682\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8469\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__8490\,
            I => \N__8466\
        );

    \I__1680\ : InMux
    port map (
            O => \N__8487\,
            I => \N__8463\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8482\,
            I => \N__8460\
        );

    \I__1678\ : InMux
    port map (
            O => \N__8481\,
            I => \N__8457\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8454\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__8475\,
            I => \N__8451\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8448\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8469\,
            I => \N__8445\
        );

    \I__1673\ : Span4Mux_h
    port map (
            O => \N__8466\,
            I => \N__8442\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8463\,
            I => \N__8437\
        );

    \I__1671\ : Span4Mux_h
    port map (
            O => \N__8460\,
            I => \N__8437\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8457\,
            I => \clk_100Khz_signalkeep\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8454\,
            I => \clk_100Khz_signalkeep\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__8451\,
            I => \clk_100Khz_signalkeep\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__8448\,
            I => \clk_100Khz_signalkeep\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__8445\,
            I => \clk_100Khz_signalkeep\
        );

    \I__1665\ : Odrv4
    port map (
            O => \N__8442\,
            I => \clk_100Khz_signalkeep\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__8437\,
            I => \clk_100Khz_signalkeep\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__8422\,
            I => \VPP_VDDQ.m6_cascade_\
        );

    \I__1662\ : CascadeMux
    port map (
            O => \N__8419\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\
        );

    \I__1661\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8413\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__8413\,
            I => \VPP_VDDQ.count_2_RNI_0Z0Z_2\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8410\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13\
        );

    \I__1658\ : InMux
    port map (
            O => \N__8407\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14\
        );

    \I__1657\ : SRMux
    port map (
            O => \N__8404\,
            I => \N__8401\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__8401\,
            I => \N__8398\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__8398\,
            I => \VPP_VDDQ.delayed_vddq_ok_RNOZ0\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__8395\,
            I => \N__8391\
        );

    \I__1653\ : InMux
    port map (
            O => \N__8394\,
            I => \N__8388\
        );

    \I__1652\ : InMux
    port map (
            O => \N__8391\,
            I => \N__8385\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8388\,
            I => \N__8382\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__8385\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7_cZ0_THRU_CO\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__8382\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7_cZ0_THRU_CO\
        );

    \I__1648\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8374\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__8374\,
            I => \VPP_VDDQ.count_2_0_8\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__8371\,
            I => \VPP_VDDQ.count_2_1_8_cascade_\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__8368\,
            I => \N__8365\
        );

    \I__1644\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8361\
        );

    \I__1643\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8358\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__8361\,
            I => \N__8353\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__8358\,
            I => \N__8353\
        );

    \I__1640\ : Odrv12
    port map (
            O => \N__8353\,
            I => \VPP_VDDQ.un1_clk_100khz_1\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__8350\,
            I => \N__8347\
        );

    \I__1638\ : InMux
    port map (
            O => \N__8347\,
            I => \N__8343\
        );

    \I__1637\ : InMux
    port map (
            O => \N__8346\,
            I => \N__8340\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__8343\,
            I => \N__8337\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__8340\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__8337\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1\
        );

    \I__1633\ : InMux
    port map (
            O => \N__8332\,
            I => \N__8329\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__8329\,
            I => \N__8325\
        );

    \I__1631\ : InMux
    port map (
            O => \N__8328\,
            I => \N__8321\
        );

    \I__1630\ : Span4Mux_h
    port map (
            O => \N__8325\,
            I => \N__8318\
        );

    \I__1629\ : InMux
    port map (
            O => \N__8324\,
            I => \N__8315\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__8321\,
            I => \VPP_VDDQ.count_2_RNI82TR_0Z0Z_1\
        );

    \I__1627\ : Odrv4
    port map (
            O => \N__8318\,
            I => \VPP_VDDQ.count_2_RNI82TR_0Z0Z_1\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__8315\,
            I => \VPP_VDDQ.count_2_RNI82TR_0Z0Z_1\
        );

    \I__1625\ : InMux
    port map (
            O => \N__8308\,
            I => \N__8304\
        );

    \I__1624\ : InMux
    port map (
            O => \N__8307\,
            I => \N__8301\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8304\,
            I => \N__8296\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__8301\,
            I => \N__8296\
        );

    \I__1621\ : Odrv12
    port map (
            O => \N__8296\,
            I => \VPP_VDDQ.delayed_vddq_ok_en\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8293\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4_cZ0\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__8290\,
            I => \N__8287\
        );

    \I__1618\ : InMux
    port map (
            O => \N__8287\,
            I => \N__8284\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__8284\,
            I => \VPP_VDDQ.un1_count_2_1_axb_6\
        );

    \I__1616\ : InMux
    port map (
            O => \N__8281\,
            I => \N__8278\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__8278\,
            I => \N__8273\
        );

    \I__1614\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8268\
        );

    \I__1613\ : InMux
    port map (
            O => \N__8276\,
            I => \N__8268\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__8273\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIVFZ0Z931\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__8268\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIVFZ0Z931\
        );

    \I__1610\ : InMux
    port map (
            O => \N__8263\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5_cZ0\
        );

    \I__1609\ : InMux
    port map (
            O => \N__8260\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6_cZ0\
        );

    \I__1608\ : InMux
    port map (
            O => \N__8257\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7_cZ0\
        );

    \I__1607\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8248\
        );

    \I__1606\ : InMux
    port map (
            O => \N__8253\,
            I => \N__8248\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__8248\,
            I => \VPP_VDDQ.un1_count_2_1_cry_8_cZ0_THRU_CO\
        );

    \I__1604\ : InMux
    port map (
            O => \N__8245\,
            I => \bfn_8_9_0_\
        );

    \I__1603\ : InMux
    port map (
            O => \N__8242\,
            I => \N__8238\
        );

    \I__1602\ : InMux
    port map (
            O => \N__8241\,
            I => \N__8235\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__8238\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9_THRU_CO\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__8235\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9_THRU_CO\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8230\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9\
        );

    \I__1598\ : InMux
    port map (
            O => \N__8227\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10\
        );

    \I__1597\ : InMux
    port map (
            O => \N__8224\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11\
        );

    \I__1596\ : InMux
    port map (
            O => \N__8221\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12\
        );

    \I__1595\ : InMux
    port map (
            O => \N__8218\,
            I => \N__8215\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__8215\,
            I => \N__8212\
        );

    \I__1593\ : Span12Mux_s5_v
    port map (
            O => \N__8212\,
            I => \N__8209\
        );

    \I__1592\ : Odrv12
    port map (
            O => \N__8209\,
            I => \VPP_VDDQ_delayed_vddq_ok\
        );

    \I__1591\ : InMux
    port map (
            O => \N__8206\,
            I => \N__8203\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__8203\,
            I => \RSMRST_PWRGD.un4_count_10\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__8200\,
            I => \N__8196\
        );

    \I__1588\ : InMux
    port map (
            O => \N__8199\,
            I => \N__8193\
        );

    \I__1587\ : InMux
    port map (
            O => \N__8196\,
            I => \N__8190\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__8193\,
            I => \VPP_VDDQ.delayed_vddq_okZ0\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__8190\,
            I => \VPP_VDDQ.delayed_vddq_okZ0\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__8185\,
            I => \VPP_VDDQ.count_2_1_3_cascade_\
        );

    \I__1583\ : InMux
    port map (
            O => \N__8182\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1_cZ0\
        );

    \I__1582\ : InMux
    port map (
            O => \N__8179\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_cZ0\
        );

    \I__1581\ : CascadeMux
    port map (
            O => \N__8176\,
            I => \N__8173\
        );

    \I__1580\ : InMux
    port map (
            O => \N__8173\,
            I => \N__8170\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__8170\,
            I => \VPP_VDDQ.un1_count_2_1_axb_4\
        );

    \I__1578\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8162\
        );

    \I__1577\ : InMux
    port map (
            O => \N__8166\,
            I => \N__8157\
        );

    \I__1576\ : InMux
    port map (
            O => \N__8165\,
            I => \N__8157\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__8162\,
            I => \N__8152\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__8157\,
            I => \N__8152\
        );

    \I__1573\ : Odrv4
    port map (
            O => \N__8152\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIRZ0Z9731\
        );

    \I__1572\ : InMux
    port map (
            O => \N__8149\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3_cZ0\
        );

    \I__1571\ : InMux
    port map (
            O => \N__8146\,
            I => \N__8143\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__8143\,
            I => \RSMRST_PWRGD.un4_count_11\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__8140\,
            I => \RSMRST_PWRGD.un4_count_8_cascade_\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__8137\,
            I => \RSMRST_PWRGD.N_1_i_cascade_\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__8134\,
            I => \RSMRST_PWRGD.N_6_cascade_\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__8131\,
            I => \RSMRST_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\
        );

    \I__1565\ : CascadeMux
    port map (
            O => \N__8128\,
            I => \G_10_cascade_\
        );

    \I__1564\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8122\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__8122\,
            I => \RSMRST_PWRGD.un4_count_9\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__8119\,
            I => \N__8114\
        );

    \I__1561\ : InMux
    port map (
            O => \N__8118\,
            I => \N__8108\
        );

    \I__1560\ : InMux
    port map (
            O => \N__8117\,
            I => \N__8108\
        );

    \I__1559\ : InMux
    port map (
            O => \N__8114\,
            I => \N__8103\
        );

    \I__1558\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8103\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__8108\,
            I => \N__8100\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__8103\,
            I => \N__8097\
        );

    \I__1555\ : Span4Mux_v
    port map (
            O => \N__8100\,
            I => \N__8093\
        );

    \I__1554\ : Span4Mux_h
    port map (
            O => \N__8097\,
            I => \N__8090\
        );

    \I__1553\ : InMux
    port map (
            O => \N__8096\,
            I => \N__8087\
        );

    \I__1552\ : Span4Mux_v
    port map (
            O => \N__8093\,
            I => \N__8084\
        );

    \I__1551\ : Span4Mux_h
    port map (
            O => \N__8090\,
            I => \N__8079\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__8087\,
            I => \N__8079\
        );

    \I__1549\ : Odrv4
    port map (
            O => \N__8084\,
            I => \RSMRST_PWRGD.N_3_i\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__8079\,
            I => \RSMRST_PWRGD.N_3_i\
        );

    \I__1547\ : InMux
    port map (
            O => \N__8074\,
            I => \N__8068\
        );

    \I__1546\ : InMux
    port map (
            O => \N__8073\,
            I => \N__8068\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__8068\,
            I => \RSMRST_PWRGD.N_1_i\
        );

    \I__1544\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8057\
        );

    \I__1543\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8050\
        );

    \I__1542\ : InMux
    port map (
            O => \N__8063\,
            I => \N__8050\
        );

    \I__1541\ : InMux
    port map (
            O => \N__8062\,
            I => \N__8050\
        );

    \I__1540\ : InMux
    port map (
            O => \N__8061\,
            I => \N__8045\
        );

    \I__1539\ : InMux
    port map (
            O => \N__8060\,
            I => \N__8045\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__8057\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__8050\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__8045\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__8038\,
            I => \RSMRST_PWRGD.i3_mux_0_cascade_\
        );

    \I__1534\ : InMux
    port map (
            O => \N__8035\,
            I => \N__8027\
        );

    \I__1533\ : InMux
    port map (
            O => \N__8034\,
            I => \N__8024\
        );

    \I__1532\ : InMux
    port map (
            O => \N__8033\,
            I => \N__8017\
        );

    \I__1531\ : InMux
    port map (
            O => \N__8032\,
            I => \N__8017\
        );

    \I__1530\ : InMux
    port map (
            O => \N__8031\,
            I => \N__8017\
        );

    \I__1529\ : InMux
    port map (
            O => \N__8030\,
            I => \N__8014\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__8027\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__8024\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__8017\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__8014\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__1524\ : InMux
    port map (
            O => \N__8005\,
            I => \N__8001\
        );

    \I__1523\ : InMux
    port map (
            O => \N__8004\,
            I => \N__7998\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__8001\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7998\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__1520\ : InMux
    port map (
            O => \N__7993\,
            I => \COUNTER.counter_1_cry_25\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__7990\,
            I => \N__7986\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7989\,
            I => \N__7983\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7986\,
            I => \N__7980\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__7983\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__7980\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7975\,
            I => \COUNTER.counter_1_cry_26\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7972\,
            I => \N__7968\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7971\,
            I => \N__7965\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7968\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7965\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7960\,
            I => \COUNTER.counter_1_cry_27\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7957\,
            I => \N__7953\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7956\,
            I => \N__7950\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7953\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7950\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7945\,
            I => \COUNTER.counter_1_cry_28\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7942\,
            I => \N__7938\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7935\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7938\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7935\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7930\,
            I => \COUNTER.counter_1_cry_29\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7927\,
            I => \COUNTER.counter_1_cry_30\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__7924\,
            I => \N__7920\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7923\,
            I => \N__7917\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7914\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7917\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__7914\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7905\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7902\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__7905\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7902\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7897\,
            I => \COUNTER.counter_1_cry_17\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__7894\,
            I => \N__7890\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7893\,
            I => \N__7887\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7890\,
            I => \N__7884\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7887\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7884\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7879\,
            I => \COUNTER.counter_1_cry_18\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7872\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7869\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7872\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7869\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7864\,
            I => \COUNTER.counter_1_cry_19\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7861\,
            I => \N__7857\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7860\,
            I => \N__7854\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7857\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7854\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7849\,
            I => \COUNTER.counter_1_cry_20\
        );

    \I__1471\ : CascadeMux
    port map (
            O => \N__7846\,
            I => \N__7842\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7845\,
            I => \N__7839\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7842\,
            I => \N__7836\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7839\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__7836\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7831\,
            I => \COUNTER.counter_1_cry_21\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7828\,
            I => \N__7824\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7827\,
            I => \N__7821\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7824\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7821\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7816\,
            I => \COUNTER.counter_1_cry_22\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7813\,
            I => \N__7809\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7806\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7809\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7806\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7801\,
            I => \COUNTER.counter_1_cry_23\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7794\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7797\,
            I => \N__7791\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7794\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__7791\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7786\,
            I => \bfn_7_14_0_\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__7783\,
            I => \N__7779\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7782\,
            I => \N__7776\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7779\,
            I => \N__7773\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7776\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7773\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7768\,
            I => \bfn_7_12_0_\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7765\,
            I => \N__7761\
        );

    \I__1443\ : InMux
    port map (
            O => \N__7764\,
            I => \N__7758\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__7761\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7758\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__1440\ : InMux
    port map (
            O => \N__7753\,
            I => \COUNTER.counter_1_cry_9\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7746\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7749\,
            I => \N__7743\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7746\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7743\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7738\,
            I => \COUNTER.counter_1_cry_10\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7735\,
            I => \N__7731\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7734\,
            I => \N__7728\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7731\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__7728\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7723\,
            I => \COUNTER.counter_1_cry_11\
        );

    \I__1429\ : InMux
    port map (
            O => \N__7720\,
            I => \N__7716\
        );

    \I__1428\ : InMux
    port map (
            O => \N__7719\,
            I => \N__7713\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__7716\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__7713\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__1425\ : InMux
    port map (
            O => \N__7708\,
            I => \COUNTER.counter_1_cry_12\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__7705\,
            I => \N__7701\
        );

    \I__1423\ : InMux
    port map (
            O => \N__7704\,
            I => \N__7698\
        );

    \I__1422\ : InMux
    port map (
            O => \N__7701\,
            I => \N__7695\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7698\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7695\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7690\,
            I => \COUNTER.counter_1_cry_13\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7687\,
            I => \N__7683\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7686\,
            I => \N__7680\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7683\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__7680\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__1414\ : InMux
    port map (
            O => \N__7675\,
            I => \COUNTER.counter_1_cry_14\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7672\,
            I => \N__7668\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7671\,
            I => \N__7665\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__7668\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__7665\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7660\,
            I => \COUNTER.counter_1_cry_15\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7657\,
            I => \N__7653\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7656\,
            I => \N__7650\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7653\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7650\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7645\,
            I => \bfn_7_13_0_\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__7642\,
            I => \N__7638\
        );

    \I__1402\ : InMux
    port map (
            O => \N__7641\,
            I => \N__7634\
        );

    \I__1401\ : InMux
    port map (
            O => \N__7638\,
            I => \N__7629\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7637\,
            I => \N__7629\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7634\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__7629\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__7624\,
            I => \N__7621\
        );

    \I__1396\ : InMux
    port map (
            O => \N__7621\,
            I => \N__7615\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7620\,
            I => \N__7608\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7619\,
            I => \N__7608\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7618\,
            I => \N__7608\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7615\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7608\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7603\,
            I => \N__7598\
        );

    \I__1389\ : InMux
    port map (
            O => \N__7602\,
            I => \N__7595\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7601\,
            I => \N__7592\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7598\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7595\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7592\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7585\,
            I => \N__7582\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__7582\,
            I => \COUNTER.counter_1_cry_1_THRU_CO\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7579\,
            I => \COUNTER.counter_1_cry_1\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7576\,
            I => \N__7571\
        );

    \I__1380\ : InMux
    port map (
            O => \N__7575\,
            I => \N__7566\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7574\,
            I => \N__7566\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__7571\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7566\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7561\,
            I => \N__7558\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__7558\,
            I => \COUNTER.counter_1_cry_2_THRU_CO\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7555\,
            I => \COUNTER.counter_1_cry_2\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__7552\,
            I => \N__7547\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7551\,
            I => \N__7544\
        );

    \I__1371\ : InMux
    port map (
            O => \N__7550\,
            I => \N__7541\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7547\,
            I => \N__7538\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__7544\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7541\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7538\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__7531\,
            I => \N__7528\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7528\,
            I => \N__7525\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7525\,
            I => \COUNTER.counter_1_cry_3_THRU_CO\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7522\,
            I => \COUNTER.counter_1_cry_3\
        );

    \I__1362\ : CascadeMux
    port map (
            O => \N__7519\,
            I => \N__7514\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7518\,
            I => \N__7511\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7517\,
            I => \N__7508\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7514\,
            I => \N__7505\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__7511\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7508\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7505\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7498\,
            I => \N__7495\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7495\,
            I => \COUNTER.counter_1_cry_4_THRU_CO\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7492\,
            I => \COUNTER.counter_1_cry_4\
        );

    \I__1352\ : InMux
    port map (
            O => \N__7489\,
            I => \N__7484\
        );

    \I__1351\ : InMux
    port map (
            O => \N__7488\,
            I => \N__7481\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7487\,
            I => \N__7478\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__7484\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__7481\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__7478\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__7471\,
            I => \N__7468\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7468\,
            I => \N__7465\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7465\,
            I => \COUNTER.counter_1_cry_5_THRU_CO\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7462\,
            I => \COUNTER.counter_1_cry_5\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7459\,
            I => \N__7455\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7458\,
            I => \N__7452\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__7455\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__7452\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7447\,
            I => \COUNTER.counter_1_cry_6\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7444\,
            I => \N__7440\
        );

    \I__1336\ : InMux
    port map (
            O => \N__7443\,
            I => \N__7437\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7440\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7437\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__1333\ : InMux
    port map (
            O => \N__7432\,
            I => \COUNTER.counter_1_cry_7\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7429\,
            I => \N__7426\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__7426\,
            I => \VPP_VDDQ.count_2_1_5\
        );

    \I__1330\ : InMux
    port map (
            O => \N__7423\,
            I => \N__7420\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__7420\,
            I => \N__7417\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__7417\,
            I => \VPP_VDDQ.count_2_0_10\
        );

    \I__1327\ : InMux
    port map (
            O => \N__7414\,
            I => \N__7409\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7413\,
            I => \N__7406\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7412\,
            I => \N__7403\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__7409\,
            I => \N__7400\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__7406\,
            I => \N__7395\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__7403\,
            I => \N__7395\
        );

    \I__1321\ : Odrv12
    port map (
            O => \N__7400\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__1320\ : Odrv4
    port map (
            O => \N__7395\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__7390\,
            I => \N__7386\
        );

    \I__1318\ : InMux
    port map (
            O => \N__7389\,
            I => \N__7383\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7379\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__7383\,
            I => \N__7376\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7382\,
            I => \N__7373\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__7379\,
            I => \N__7370\
        );

    \I__1313\ : Odrv12
    port map (
            O => \N__7376\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__7373\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__1311\ : Odrv4
    port map (
            O => \N__7370\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__1310\ : InMux
    port map (
            O => \N__7363\,
            I => \N__7360\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__7360\,
            I => \N__7357\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__7357\,
            I => \VPP_VDDQ.count_2_1_6\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__7354\,
            I => \VPP_VDDQ.count_2_1_1_cascade_\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7351\,
            I => \N__7348\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__7348\,
            I => \N__7344\
        );

    \I__1304\ : InMux
    port map (
            O => \N__7347\,
            I => \N__7341\
        );

    \I__1303\ : Odrv4
    port map (
            O => \N__7344\,
            I => \VPP_VDDQ.count_2_1_4\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__7341\,
            I => \VPP_VDDQ.count_2_1_4\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7336\,
            I => \N__7333\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__7333\,
            I => \VPP_VDDQ.count_2_RNI25V3Z0Z_1\
        );

    \I__1299\ : CascadeMux
    port map (
            O => \N__7330\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIZ0_cascade_\
        );

    \I__1298\ : CascadeMux
    port map (
            O => \N__7327\,
            I => \VPP_VDDQ.m4_1_cascade_\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__7324\,
            I => \N__7320\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__7323\,
            I => \N__7317\
        );

    \I__1295\ : InMux
    port map (
            O => \N__7320\,
            I => \N__7314\
        );

    \I__1294\ : InMux
    port map (
            O => \N__7317\,
            I => \N__7310\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7314\,
            I => \N__7307\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__7313\,
            I => \N__7304\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__7310\,
            I => \N__7301\
        );

    \I__1290\ : Span4Mux_h
    port map (
            O => \N__7307\,
            I => \N__7298\
        );

    \I__1289\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7295\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__7301\,
            I => \VPP_VDDQ.curr_state_2_e_0_RNINUSCZ0Z_1\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__7298\,
            I => \VPP_VDDQ.curr_state_2_e_0_RNINUSCZ0Z_1\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__7295\,
            I => \VPP_VDDQ.curr_state_2_e_0_RNINUSCZ0Z_1\
        );

    \I__1285\ : InMux
    port map (
            O => \N__7288\,
            I => \N__7285\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__7285\,
            I => \VPP_VDDQ.count_2_1_1\
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__7282\,
            I => \VPP_VDDQ.count_2_1_6_cascade_\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__7279\,
            I => \N__7276\
        );

    \I__1281\ : InMux
    port map (
            O => \N__7276\,
            I => \N__7273\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__7273\,
            I => \VPP_VDDQ.g0_3_a3_0_1\
        );

    \I__1279\ : InMux
    port map (
            O => \N__7270\,
            I => \N__7267\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__7267\,
            I => \VPP_VDDQ.N_6\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__7264\,
            I => \VPP_VDDQ.count_2_1_9_cascade_\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__7261\,
            I => \VPP_VDDQ.count_2Z0Z_9_cascade_\
        );

    \I__1275\ : InMux
    port map (
            O => \N__7258\,
            I => \N__7255\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__7255\,
            I => \VPP_VDDQ.count_2_0_9\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__7252\,
            I => \N__7249\
        );

    \I__1272\ : InMux
    port map (
            O => \N__7249\,
            I => \N__7246\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__7246\,
            I => \N__7243\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__7243\,
            I => \COUNTER.un4_counter_5_and\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__7240\,
            I => \N__7237\
        );

    \I__1268\ : InMux
    port map (
            O => \N__7237\,
            I => \N__7234\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__7234\,
            I => \N__7231\
        );

    \I__1266\ : Span4Mux_h
    port map (
            O => \N__7231\,
            I => \N__7228\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__7228\,
            I => \COUNTER.un4_counter_7_and\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__7225\,
            I => \N__7222\
        );

    \I__1263\ : InMux
    port map (
            O => \N__7222\,
            I => \N__7219\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__7219\,
            I => \N__7216\
        );

    \I__1261\ : Odrv12
    port map (
            O => \N__7216\,
            I => \COUNTER.un4_counter_6_and\
        );

    \I__1260\ : InMux
    port map (
            O => \N__7213\,
            I => \N__7210\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__7210\,
            I => \N__7207\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__7207\,
            I => \N__7204\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__7204\,
            I => \RSMRST_PWRGD.curr_state10\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__7201\,
            I => \N__7186\
        );

    \I__1255\ : InMux
    port map (
            O => \N__7200\,
            I => \N__7175\
        );

    \I__1254\ : InMux
    port map (
            O => \N__7199\,
            I => \N__7164\
        );

    \I__1253\ : InMux
    port map (
            O => \N__7198\,
            I => \N__7164\
        );

    \I__1252\ : InMux
    port map (
            O => \N__7197\,
            I => \N__7164\
        );

    \I__1251\ : InMux
    port map (
            O => \N__7196\,
            I => \N__7164\
        );

    \I__1250\ : InMux
    port map (
            O => \N__7195\,
            I => \N__7164\
        );

    \I__1249\ : InMux
    port map (
            O => \N__7194\,
            I => \N__7161\
        );

    \I__1248\ : CascadeMux
    port map (
            O => \N__7193\,
            I => \N__7156\
        );

    \I__1247\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7149\
        );

    \I__1246\ : InMux
    port map (
            O => \N__7191\,
            I => \N__7149\
        );

    \I__1245\ : InMux
    port map (
            O => \N__7190\,
            I => \N__7146\
        );

    \I__1244\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7137\
        );

    \I__1243\ : InMux
    port map (
            O => \N__7186\,
            I => \N__7137\
        );

    \I__1242\ : InMux
    port map (
            O => \N__7185\,
            I => \N__7137\
        );

    \I__1241\ : InMux
    port map (
            O => \N__7184\,
            I => \N__7137\
        );

    \I__1240\ : InMux
    port map (
            O => \N__7183\,
            I => \N__7130\
        );

    \I__1239\ : InMux
    port map (
            O => \N__7182\,
            I => \N__7119\
        );

    \I__1238\ : InMux
    port map (
            O => \N__7181\,
            I => \N__7119\
        );

    \I__1237\ : InMux
    port map (
            O => \N__7180\,
            I => \N__7119\
        );

    \I__1236\ : InMux
    port map (
            O => \N__7179\,
            I => \N__7119\
        );

    \I__1235\ : InMux
    port map (
            O => \N__7178\,
            I => \N__7119\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__7175\,
            I => \N__7112\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__7164\,
            I => \N__7112\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__7161\,
            I => \N__7112\
        );

    \I__1231\ : InMux
    port map (
            O => \N__7160\,
            I => \N__7109\
        );

    \I__1230\ : InMux
    port map (
            O => \N__7159\,
            I => \N__7106\
        );

    \I__1229\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7103\
        );

    \I__1228\ : InMux
    port map (
            O => \N__7155\,
            I => \N__7098\
        );

    \I__1227\ : InMux
    port map (
            O => \N__7154\,
            I => \N__7098\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__7149\,
            I => \N__7095\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__7146\,
            I => \N__7092\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__7137\,
            I => \N__7089\
        );

    \I__1223\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7084\
        );

    \I__1222\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7084\
        );

    \I__1221\ : InMux
    port map (
            O => \N__7134\,
            I => \N__7079\
        );

    \I__1220\ : InMux
    port map (
            O => \N__7133\,
            I => \N__7079\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__7130\,
            I => \N__7072\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__7119\,
            I => \N__7072\
        );

    \I__1217\ : Span4Mux_v
    port map (
            O => \N__7112\,
            I => \N__7072\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__7109\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__7106\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__7103\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__7098\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1212\ : Odrv4
    port map (
            O => \N__7095\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__7092\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__7089\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__7084\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__7079\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__7072\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__1206\ : InMux
    port map (
            O => \N__7051\,
            I => \N__7047\
        );

    \I__1205\ : InMux
    port map (
            O => \N__7050\,
            I => \N__7044\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__7047\,
            I => \N__7041\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__7044\,
            I => \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7\
        );

    \I__1202\ : Odrv4
    port map (
            O => \N__7041\,
            I => \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__7036\,
            I => \N__7033\
        );

    \I__1200\ : InMux
    port map (
            O => \N__7033\,
            I => \N__7027\
        );

    \I__1199\ : InMux
    port map (
            O => \N__7032\,
            I => \N__7027\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__7027\,
            I => \N__7024\
        );

    \I__1197\ : Span4Mux_h
    port map (
            O => \N__7024\,
            I => \N__7021\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__7021\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__1195\ : InMux
    port map (
            O => \N__7018\,
            I => \N__7013\
        );

    \I__1194\ : CascadeMux
    port map (
            O => \N__7017\,
            I => \N__7010\
        );

    \I__1193\ : InMux
    port map (
            O => \N__7016\,
            I => \N__7007\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__7013\,
            I => \N__7004\
        );

    \I__1191\ : InMux
    port map (
            O => \N__7010\,
            I => \N__7001\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__7007\,
            I => \N__6998\
        );

    \I__1189\ : Odrv12
    port map (
            O => \N__7004\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__7001\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__6998\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__6991\,
            I => \N__6987\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6990\,
            I => \N__6982\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6987\,
            I => \N__6982\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6982\,
            I => \N__6979\
        );

    \I__1182\ : Span4Mux_h
    port map (
            O => \N__6979\,
            I => \N__6976\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__6976\,
            I => \PCH_PWRGD.countZ0Z_10\
        );

    \I__1180\ : CEMux
    port map (
            O => \N__6973\,
            I => \N__6969\
        );

    \I__1179\ : CEMux
    port map (
            O => \N__6972\,
            I => \N__6957\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6969\,
            I => \N__6954\
        );

    \I__1177\ : CEMux
    port map (
            O => \N__6968\,
            I => \N__6951\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6967\,
            I => \N__6946\
        );

    \I__1175\ : CEMux
    port map (
            O => \N__6966\,
            I => \N__6946\
        );

    \I__1174\ : CEMux
    port map (
            O => \N__6965\,
            I => \N__6943\
        );

    \I__1173\ : CascadeMux
    port map (
            O => \N__6964\,
            I => \N__6937\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6963\,
            I => \N__6933\
        );

    \I__1171\ : CEMux
    port map (
            O => \N__6962\,
            I => \N__6929\
        );

    \I__1170\ : CEMux
    port map (
            O => \N__6961\,
            I => \N__6926\
        );

    \I__1169\ : CEMux
    port map (
            O => \N__6960\,
            I => \N__6923\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6957\,
            I => \N__6920\
        );

    \I__1167\ : Span4Mux_h
    port map (
            O => \N__6954\,
            I => \N__6906\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6951\,
            I => \N__6906\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6946\,
            I => \N__6906\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__6943\,
            I => \N__6906\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6942\,
            I => \N__6899\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6899\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6899\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6894\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6936\,
            I => \N__6894\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6933\,
            I => \N__6891\
        );

    \I__1157\ : CEMux
    port map (
            O => \N__6932\,
            I => \N__6888\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6929\,
            I => \N__6883\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6926\,
            I => \N__6876\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6923\,
            I => \N__6873\
        );

    \I__1153\ : Span4Mux_s3_v
    port map (
            O => \N__6920\,
            I => \N__6870\
        );

    \I__1152\ : InMux
    port map (
            O => \N__6919\,
            I => \N__6865\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6918\,
            I => \N__6865\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6917\,
            I => \N__6858\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6916\,
            I => \N__6858\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6915\,
            I => \N__6858\
        );

    \I__1147\ : Span4Mux_v
    port map (
            O => \N__6906\,
            I => \N__6855\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6899\,
            I => \N__6852\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6894\,
            I => \N__6847\
        );

    \I__1144\ : Span4Mux_v
    port map (
            O => \N__6891\,
            I => \N__6847\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6888\,
            I => \N__6844\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6887\,
            I => \N__6839\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6886\,
            I => \N__6839\
        );

    \I__1140\ : Span4Mux_h
    port map (
            O => \N__6883\,
            I => \N__6836\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6882\,
            I => \N__6831\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6831\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6826\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6879\,
            I => \N__6826\
        );

    \I__1135\ : Span4Mux_h
    port map (
            O => \N__6876\,
            I => \N__6815\
        );

    \I__1134\ : Span4Mux_h
    port map (
            O => \N__6873\,
            I => \N__6815\
        );

    \I__1133\ : Span4Mux_h
    port map (
            O => \N__6870\,
            I => \N__6815\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6865\,
            I => \N__6815\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6858\,
            I => \N__6815\
        );

    \I__1130\ : Span4Mux_s2_v
    port map (
            O => \N__6855\,
            I => \N__6810\
        );

    \I__1129\ : Span4Mux_h
    port map (
            O => \N__6852\,
            I => \N__6810\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__6847\,
            I => \PCH_PWRGD.curr_state_e_0_RNI4GQL2Z0Z_0\
        );

    \I__1127\ : Odrv12
    port map (
            O => \N__6844\,
            I => \PCH_PWRGD.curr_state_e_0_RNI4GQL2Z0Z_0\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6839\,
            I => \PCH_PWRGD.curr_state_e_0_RNI4GQL2Z0Z_0\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__6836\,
            I => \PCH_PWRGD.curr_state_e_0_RNI4GQL2Z0Z_0\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6831\,
            I => \PCH_PWRGD.curr_state_e_0_RNI4GQL2Z0Z_0\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6826\,
            I => \PCH_PWRGD.curr_state_e_0_RNI4GQL2Z0Z_0\
        );

    \I__1122\ : Odrv4
    port map (
            O => \N__6815\,
            I => \PCH_PWRGD.curr_state_e_0_RNI4GQL2Z0Z_0\
        );

    \I__1121\ : Odrv4
    port map (
            O => \N__6810\,
            I => \PCH_PWRGD.curr_state_e_0_RNI4GQL2Z0Z_0\
        );

    \I__1120\ : SRMux
    port map (
            O => \N__6793\,
            I => \N__6783\
        );

    \I__1119\ : SRMux
    port map (
            O => \N__6792\,
            I => \N__6780\
        );

    \I__1118\ : SRMux
    port map (
            O => \N__6791\,
            I => \N__6777\
        );

    \I__1117\ : SRMux
    port map (
            O => \N__6790\,
            I => \N__6774\
        );

    \I__1116\ : SRMux
    port map (
            O => \N__6789\,
            I => \N__6771\
        );

    \I__1115\ : SRMux
    port map (
            O => \N__6788\,
            I => \N__6768\
        );

    \I__1114\ : SRMux
    port map (
            O => \N__6787\,
            I => \N__6764\
        );

    \I__1113\ : SRMux
    port map (
            O => \N__6786\,
            I => \N__6761\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6783\,
            I => \N__6758\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__6780\,
            I => \N__6755\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6777\,
            I => \N__6748\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6774\,
            I => \N__6748\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6771\,
            I => \N__6748\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6768\,
            I => \N__6745\
        );

    \I__1106\ : SRMux
    port map (
            O => \N__6767\,
            I => \N__6742\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6764\,
            I => \N__6739\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6761\,
            I => \N__6736\
        );

    \I__1103\ : Span4Mux_v
    port map (
            O => \N__6758\,
            I => \N__6733\
        );

    \I__1102\ : Span4Mux_v
    port map (
            O => \N__6755\,
            I => \N__6728\
        );

    \I__1101\ : Span4Mux_v
    port map (
            O => \N__6748\,
            I => \N__6728\
        );

    \I__1100\ : Span4Mux_v
    port map (
            O => \N__6745\,
            I => \N__6723\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6742\,
            I => \N__6723\
        );

    \I__1098\ : Span4Mux_h
    port map (
            O => \N__6739\,
            I => \N__6720\
        );

    \I__1097\ : Odrv12
    port map (
            O => \N__6736\,
            I => \PCH_PWRGD.count_m2_0_a2_iso\
        );

    \I__1096\ : Odrv4
    port map (
            O => \N__6733\,
            I => \PCH_PWRGD.count_m2_0_a2_iso\
        );

    \I__1095\ : Odrv4
    port map (
            O => \N__6728\,
            I => \PCH_PWRGD.count_m2_0_a2_iso\
        );

    \I__1094\ : Odrv4
    port map (
            O => \N__6723\,
            I => \PCH_PWRGD.count_m2_0_a2_iso\
        );

    \I__1093\ : Odrv4
    port map (
            O => \N__6720\,
            I => \PCH_PWRGD.count_m2_0_a2_iso\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__6709\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7_cascade_\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__6706\,
            I => \N__6703\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6703\,
            I => \N__6700\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__6700\,
            I => \N__6697\
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__6697\,
            I => \COUNTER.un4_counter_2_and\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__6694\,
            I => \N__6691\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6688\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6688\,
            I => \N__6685\
        );

    \I__1084\ : Odrv4
    port map (
            O => \N__6685\,
            I => \COUNTER.un4_counter_3_and\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__6682\,
            I => \N__6679\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6676\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__6676\,
            I => \N__6673\
        );

    \I__1080\ : Odrv4
    port map (
            O => \N__6673\,
            I => \COUNTER.un4_counter_4_and\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6670\,
            I => \bfn_6_10_0_\
        );

    \I__1078\ : CascadeMux
    port map (
            O => \N__6667\,
            I => \COUNTER_un4_counter_7_THRU_CO_cascade_\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__6664\,
            I => \N__6661\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6658\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6658\,
            I => \COUNTER.un4_counter_0_and\
        );

    \I__1074\ : CascadeMux
    port map (
            O => \N__6655\,
            I => \N__6652\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6652\,
            I => \N__6649\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__6649\,
            I => \COUNTER.un4_counter_1_and\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6646\,
            I => \N__6640\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6645\,
            I => \N__6640\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6640\,
            I => \PCH_PWRGD.un2_count_1_cry_11_c_RNI96OZ0Z7\
        );

    \I__1068\ : InMux
    port map (
            O => \N__6637\,
            I => \N__6633\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6630\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6633\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__6630\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__6625\,
            I => \PCH_PWRGD.count_rst_7_cascade_\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6622\,
            I => \N__6619\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__6619\,
            I => \N__6616\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__6616\,
            I => \PCH_PWRGD.count_0_7\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6607\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6612\,
            I => \N__6604\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6611\,
            I => \N__6601\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6598\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6607\,
            I => \N__6595\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__6604\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__6601\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__6598\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__1052\ : Odrv4
    port map (
            O => \N__6595\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__6586\,
            I => \N__6582\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__6585\,
            I => \N__6579\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6576\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6579\,
            I => \N__6573\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__6576\,
            I => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6573\,
            I => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__6568\,
            I => \PCH_PWRGD.count_rst_6_cascade_\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6565\,
            I => \N__6562\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6562\,
            I => \PCH_PWRGD.count_0_8\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6559\,
            I => \N__6556\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__6556\,
            I => \N__6553\
        );

    \I__1040\ : Span4Mux_v
    port map (
            O => \N__6553\,
            I => \N__6547\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6552\,
            I => \N__6544\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6551\,
            I => \N__6541\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6538\
        );

    \I__1036\ : Odrv4
    port map (
            O => \N__6547\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6544\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6541\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6538\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__6529\,
            I => \PCH_PWRGD.count_rst_5_cascade_\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__6526\,
            I => \N__6523\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6523\,
            I => \N__6520\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6520\,
            I => \N__6516\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__6519\,
            I => \N__6512\
        );

    \I__1027\ : Span4Mux_v
    port map (
            O => \N__6516\,
            I => \N__6509\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6515\,
            I => \N__6506\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6512\,
            I => \N__6503\
        );

    \I__1024\ : Odrv4
    port map (
            O => \N__6509\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__6506\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6503\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6490\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6495\,
            I => \N__6490\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6490\,
            I => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\
        );

    \I__1018\ : CascadeMux
    port map (
            O => \N__6487\,
            I => \PCH_PWRGD.countZ0Z_9_cascade_\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6469\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6483\,
            I => \N__6469\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6482\,
            I => \N__6469\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6481\,
            I => \N__6457\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6457\
        );

    \I__1012\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6457\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6457\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6477\,
            I => \N__6457\
        );

    \I__1009\ : CascadeMux
    port map (
            O => \N__6476\,
            I => \N__6451\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6469\,
            I => \N__6443\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6440\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6457\,
            I => \N__6437\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6456\,
            I => \N__6434\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6455\,
            I => \N__6427\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6454\,
            I => \N__6427\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6451\,
            I => \N__6424\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6450\,
            I => \N__6421\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6449\,
            I => \N__6412\
        );

    \I__999\ : InMux
    port map (
            O => \N__6448\,
            I => \N__6412\
        );

    \I__998\ : InMux
    port map (
            O => \N__6447\,
            I => \N__6412\
        );

    \I__997\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6412\
        );

    \I__996\ : Span4Mux_v
    port map (
            O => \N__6443\,
            I => \N__6409\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__6440\,
            I => \N__6404\
        );

    \I__994\ : Span4Mux_h
    port map (
            O => \N__6437\,
            I => \N__6404\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__6434\,
            I => \N__6401\
        );

    \I__992\ : InMux
    port map (
            O => \N__6433\,
            I => \N__6396\
        );

    \I__991\ : InMux
    port map (
            O => \N__6432\,
            I => \N__6396\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__6427\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__6424\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__6421\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__6412\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__6409\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__985\ : Odrv4
    port map (
            O => \N__6404\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__984\ : Odrv4
    port map (
            O => \N__6401\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__6396\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__982\ : InMux
    port map (
            O => \N__6379\,
            I => \N__6376\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__6376\,
            I => \N__6373\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__6373\,
            I => \PCH_PWRGD.count_0_9\
        );

    \I__979\ : InMux
    port map (
            O => \N__6370\,
            I => \N__6367\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__6367\,
            I => \N__6364\
        );

    \I__977\ : Odrv4
    port map (
            O => \N__6364\,
            I => \PCH_PWRGD.count_rst_2\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__6361\,
            I => \PCH_PWRGD.count_rst_2_cascade_\
        );

    \I__975\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6355\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__6355\,
            I => \PCH_PWRGD.un2_count_1_axb_12\
        );

    \I__973\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6347\
        );

    \I__972\ : InMux
    port map (
            O => \N__6351\,
            I => \N__6342\
        );

    \I__971\ : InMux
    port map (
            O => \N__6350\,
            I => \N__6342\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__6347\,
            I => \PCH_PWRGD.count_rst_12\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__6342\,
            I => \PCH_PWRGD.count_rst_12\
        );

    \I__968\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6334\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__6334\,
            I => \N__6330\
        );

    \I__966\ : InMux
    port map (
            O => \N__6333\,
            I => \N__6327\
        );

    \I__965\ : Odrv4
    port map (
            O => \N__6330\,
            I => \PCH_PWRGD.countZ0Z_2\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__6327\,
            I => \PCH_PWRGD.countZ0Z_2\
        );

    \I__963\ : InMux
    port map (
            O => \N__6322\,
            I => \N__6319\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__6319\,
            I => \N__6316\
        );

    \I__961\ : Span4Mux_h
    port map (
            O => \N__6316\,
            I => \N__6313\
        );

    \I__960\ : Odrv4
    port map (
            O => \N__6313\,
            I => \PCH_PWRGD_N_3\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__6310\,
            I => \N__6307\
        );

    \I__958\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6302\
        );

    \I__957\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6298\
        );

    \I__956\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6295\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__6302\,
            I => \N__6292\
        );

    \I__954\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6289\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__6298\,
            I => \N__6286\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__6295\,
            I => \N__6283\
        );

    \I__951\ : Span4Mux_h
    port map (
            O => \N__6292\,
            I => \N__6280\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__6289\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__949\ : Odrv4
    port map (
            O => \N__6286\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__948\ : Odrv4
    port map (
            O => \N__6283\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__947\ : Odrv4
    port map (
            O => \N__6280\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__946\ : InMux
    port map (
            O => \N__6271\,
            I => \N__6268\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__6268\,
            I => \PCH_PWRGD.count_rst_11\
        );

    \I__944\ : CascadeMux
    port map (
            O => \N__6265\,
            I => \PCH_PWRGD.curr_state_e_0_RNI4GQL2Z0Z_0_cascade_\
        );

    \I__943\ : InMux
    port map (
            O => \N__6262\,
            I => \N__6259\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__6259\,
            I => \PCH_PWRGD.count_0_3\
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__6256\,
            I => \N__6253\
        );

    \I__940\ : InMux
    port map (
            O => \N__6253\,
            I => \N__6250\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__6250\,
            I => \N__6244\
        );

    \I__938\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6239\
        );

    \I__937\ : InMux
    port map (
            O => \N__6248\,
            I => \N__6239\
        );

    \I__936\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6236\
        );

    \I__935\ : Odrv4
    port map (
            O => \N__6244\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__6239\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__6236\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__932\ : CascadeMux
    port map (
            O => \N__6229\,
            I => \N__6226\
        );

    \I__931\ : InMux
    port map (
            O => \N__6226\,
            I => \N__6223\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__6223\,
            I => \N__6219\
        );

    \I__929\ : InMux
    port map (
            O => \N__6222\,
            I => \N__6216\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__6219\,
            I => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__6216\,
            I => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\
        );

    \I__926\ : CascadeMux
    port map (
            O => \N__6211\,
            I => \N__6207\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__6210\,
            I => \N__6204\
        );

    \I__924\ : InMux
    port map (
            O => \N__6207\,
            I => \N__6199\
        );

    \I__923\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6196\
        );

    \I__922\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6193\
        );

    \I__921\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6190\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__6199\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__6196\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__6193\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__6190\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__916\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6178\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__6178\,
            I => \PCH_PWRGD.count_rst_9\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__6175\,
            I => \PCH_PWRGD.count_rst_3_cascade_\
        );

    \I__913\ : InMux
    port map (
            O => \N__6172\,
            I => \N__6169\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__6169\,
            I => \N__6166\
        );

    \I__911\ : Span4Mux_v
    port map (
            O => \N__6166\,
            I => \N__6162\
        );

    \I__910\ : InMux
    port map (
            O => \N__6165\,
            I => \N__6159\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__6162\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__6159\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__907\ : InMux
    port map (
            O => \N__6154\,
            I => \N__6148\
        );

    \I__906\ : InMux
    port map (
            O => \N__6153\,
            I => \N__6148\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__6148\,
            I => \PCH_PWRGD.un2_count_1_cry_10_c_RNI84NZ0Z7\
        );

    \I__904\ : InMux
    port map (
            O => \N__6145\,
            I => \N__6142\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__6142\,
            I => \PCH_PWRGD.count_0_11\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__6139\,
            I => \N__6136\
        );

    \I__901\ : InMux
    port map (
            O => \N__6136\,
            I => \N__6132\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__6135\,
            I => \N__6129\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__6132\,
            I => \N__6126\
        );

    \I__898\ : InMux
    port map (
            O => \N__6129\,
            I => \N__6123\
        );

    \I__897\ : Odrv4
    port map (
            O => \N__6126\,
            I => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__6123\,
            I => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__895\ : SRMux
    port map (
            O => \N__6118\,
            I => \N__6114\
        );

    \I__894\ : SRMux
    port map (
            O => \N__6117\,
            I => \N__6111\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__6114\,
            I => \N__6107\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__6111\,
            I => \N__6104\
        );

    \I__891\ : SRMux
    port map (
            O => \N__6110\,
            I => \N__6101\
        );

    \I__890\ : Span4Mux_h
    port map (
            O => \N__6107\,
            I => \N__6097\
        );

    \I__889\ : Span4Mux_h
    port map (
            O => \N__6104\,
            I => \N__6092\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__6101\,
            I => \N__6092\
        );

    \I__887\ : InMux
    port map (
            O => \N__6100\,
            I => \N__6089\
        );

    \I__886\ : Odrv4
    port map (
            O => \N__6097\,
            I => \G_24\
        );

    \I__885\ : Odrv4
    port map (
            O => \N__6092\,
            I => \G_24\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__6089\,
            I => \G_24\
        );

    \I__883\ : CEMux
    port map (
            O => \N__6082\,
            I => \N__6079\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__6079\,
            I => \N__6076\
        );

    \I__881\ : Sp12to4
    port map (
            O => \N__6076\,
            I => \N__6073\
        );

    \I__880\ : Odrv12
    port map (
            O => \N__6073\,
            I => \VPP_VDDQ.N_9_1\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__6070\,
            I => \N__6064\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__6069\,
            I => \N__6060\
        );

    \I__877\ : InMux
    port map (
            O => \N__6068\,
            I => \N__6050\
        );

    \I__876\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6050\
        );

    \I__875\ : InMux
    port map (
            O => \N__6064\,
            I => \N__6050\
        );

    \I__874\ : InMux
    port map (
            O => \N__6063\,
            I => \N__6050\
        );

    \I__873\ : InMux
    port map (
            O => \N__6060\,
            I => \N__6045\
        );

    \I__872\ : InMux
    port map (
            O => \N__6059\,
            I => \N__6045\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__6050\,
            I => \VPP_VDDQ.curr_stateZ1Z_0\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__6045\,
            I => \VPP_VDDQ.curr_stateZ1Z_0\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__6040\,
            I => \N__6031\
        );

    \I__868\ : InMux
    port map (
            O => \N__6039\,
            I => \N__6022\
        );

    \I__867\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6022\
        );

    \I__866\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6022\
        );

    \I__865\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6022\
        );

    \I__864\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6015\
        );

    \I__863\ : InMux
    port map (
            O => \N__6034\,
            I => \N__6015\
        );

    \I__862\ : InMux
    port map (
            O => \N__6031\,
            I => \N__6015\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__6022\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__6015\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__859\ : InMux
    port map (
            O => \N__6010\,
            I => \N__6007\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__6007\,
            I => \VPP_VDDQ.un1_curr_state12_0\
        );

    \I__857\ : InMux
    port map (
            O => \N__6004\,
            I => \N__5992\
        );

    \I__856\ : InMux
    port map (
            O => \N__6003\,
            I => \N__5992\
        );

    \I__855\ : InMux
    port map (
            O => \N__6002\,
            I => \N__5992\
        );

    \I__854\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5992\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5992\,
            I => \VPP_VDDQ.un1_vddq_pwrgdZ0\
        );

    \I__852\ : InMux
    port map (
            O => \N__5989\,
            I => \N__5985\
        );

    \I__851\ : InMux
    port map (
            O => \N__5988\,
            I => \N__5982\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5985\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5982\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__848\ : IoInMux
    port map (
            O => \N__5977\,
            I => \N__5974\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__5974\,
            I => \N__5970\
        );

    \I__846\ : InMux
    port map (
            O => \N__5973\,
            I => \N__5966\
        );

    \I__845\ : IoSpan4Mux
    port map (
            O => \N__5970\,
            I => \N__5961\
        );

    \I__844\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5958\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__5966\,
            I => \N__5955\
        );

    \I__842\ : InMux
    port map (
            O => \N__5965\,
            I => \N__5950\
        );

    \I__841\ : InMux
    port map (
            O => \N__5964\,
            I => \N__5950\
        );

    \I__840\ : Span4Mux_s3_h
    port map (
            O => \N__5961\,
            I => \N__5947\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5958\,
            I => \N__5944\
        );

    \I__838\ : Span4Mux_v
    port map (
            O => \N__5955\,
            I => \N__5939\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5950\,
            I => \N__5939\
        );

    \I__836\ : Odrv4
    port map (
            O => \N__5947\,
            I => vccst_en
        );

    \I__835\ : Odrv12
    port map (
            O => \N__5944\,
            I => vccst_en
        );

    \I__834\ : Odrv4
    port map (
            O => \N__5939\,
            I => vccst_en
        );

    \I__833\ : IoInMux
    port map (
            O => \N__5932\,
            I => \N__5929\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5929\,
            I => \N__5926\
        );

    \I__831\ : Odrv12
    port map (
            O => \N__5926\,
            I => vpp_en
        );

    \I__830\ : IoInMux
    port map (
            O => \N__5923\,
            I => \N__5920\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__5920\,
            I => \N__5916\
        );

    \I__828\ : IoInMux
    port map (
            O => \N__5919\,
            I => \N__5913\
        );

    \I__827\ : IoSpan4Mux
    port map (
            O => \N__5916\,
            I => \N__5910\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5913\,
            I => \N__5906\
        );

    \I__825\ : Span4Mux_s0_v
    port map (
            O => \N__5910\,
            I => \N__5903\
        );

    \I__824\ : InMux
    port map (
            O => \N__5909\,
            I => \N__5900\
        );

    \I__823\ : IoSpan4Mux
    port map (
            O => \N__5906\,
            I => \N__5897\
        );

    \I__822\ : Span4Mux_h
    port map (
            O => \N__5903\,
            I => \N__5892\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5900\,
            I => \N__5892\
        );

    \I__820\ : Span4Mux_s3_h
    port map (
            O => \N__5897\,
            I => \N__5889\
        );

    \I__819\ : Span4Mux_v
    port map (
            O => \N__5892\,
            I => \N__5886\
        );

    \I__818\ : Span4Mux_v
    port map (
            O => \N__5889\,
            I => \N__5883\
        );

    \I__817\ : Span4Mux_v
    port map (
            O => \N__5886\,
            I => \N__5880\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__5883\,
            I => pch_pwrok
        );

    \I__815\ : Odrv4
    port map (
            O => \N__5880\,
            I => pch_pwrok
        );

    \I__814\ : IoInMux
    port map (
            O => \N__5875\,
            I => \N__5872\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5872\,
            I => \N__5869\
        );

    \I__812\ : Odrv12
    port map (
            O => \N__5869\,
            I => vccst_pwrgd
        );

    \I__811\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5863\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__5863\,
            I => \PCH_PWRGD.un2_count_1_axb_6\
        );

    \I__809\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5857\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5857\,
            I => \N__5852\
        );

    \I__807\ : InMux
    port map (
            O => \N__5856\,
            I => \N__5847\
        );

    \I__806\ : InMux
    port map (
            O => \N__5855\,
            I => \N__5847\
        );

    \I__805\ : Odrv4
    port map (
            O => \N__5852\,
            I => \PCH_PWRGD.count_rst_8\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5847\,
            I => \PCH_PWRGD.count_rst_8\
        );

    \I__803\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5839\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5839\,
            I => \N__5835\
        );

    \I__801\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5832\
        );

    \I__800\ : Odrv4
    port map (
            O => \N__5835\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__5832\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__798\ : InMux
    port map (
            O => \N__5827\,
            I => \N__5824\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5824\,
            I => \PCH_PWRGD.un2_count_1_axb_2\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__5821\,
            I => \VPP_VDDQ_un6_count_cascade_\
        );

    \I__795\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5815\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__5815\,
            I => \VPP_VDDQ_curr_state12\
        );

    \I__793\ : InMux
    port map (
            O => \N__5812\,
            I => \N__5808\
        );

    \I__792\ : InMux
    port map (
            O => \N__5811\,
            I => \N__5805\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__5808\,
            I => \N__5800\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5805\,
            I => \N__5800\
        );

    \I__789\ : Odrv4
    port map (
            O => \N__5800\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__788\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5793\
        );

    \I__787\ : InMux
    port map (
            O => \N__5796\,
            I => \N__5790\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5793\,
            I => \N__5787\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5790\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__784\ : Odrv12
    port map (
            O => \N__5787\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__5782\,
            I => \N__5778\
        );

    \I__782\ : InMux
    port map (
            O => \N__5781\,
            I => \N__5775\
        );

    \I__781\ : InMux
    port map (
            O => \N__5778\,
            I => \N__5772\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5775\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5772\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__778\ : InMux
    port map (
            O => \N__5767\,
            I => \N__5763\
        );

    \I__777\ : InMux
    port map (
            O => \N__5766\,
            I => \N__5760\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__5763\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5760\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__774\ : InMux
    port map (
            O => \N__5755\,
            I => \N__5752\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__5752\,
            I => \VPP_VDDQ.un6_count_10\
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__5749\,
            I => \N__5745\
        );

    \I__771\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5742\
        );

    \I__770\ : InMux
    port map (
            O => \N__5745\,
            I => \N__5739\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5742\,
            I => \VPP_VDDQ.un1_curr_state13_0\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5739\,
            I => \VPP_VDDQ.un1_curr_state13_0\
        );

    \I__767\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5731\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5731\,
            I => \VPP_VDDQ_un6_count\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__764\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5719\
        );

    \I__763\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5719\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__5719\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_1_sqmuxa\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__5716\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_1_sqmuxa_cascade_\
        );

    \I__760\ : InMux
    port map (
            O => \N__5713\,
            I => \N__5710\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5710\,
            I => \VPP_VDDQ.curr_state11\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__5707\,
            I => \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__5704\,
            I => \N__5700\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__5703\,
            I => \N__5695\
        );

    \I__755\ : InMux
    port map (
            O => \N__5700\,
            I => \N__5691\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__5699\,
            I => \N__5686\
        );

    \I__753\ : InMux
    port map (
            O => \N__5698\,
            I => \N__5679\
        );

    \I__752\ : InMux
    port map (
            O => \N__5695\,
            I => \N__5679\
        );

    \I__751\ : InMux
    port map (
            O => \N__5694\,
            I => \N__5679\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__5691\,
            I => \N__5676\
        );

    \I__749\ : InMux
    port map (
            O => \N__5690\,
            I => \N__5669\
        );

    \I__748\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5669\
        );

    \I__747\ : InMux
    port map (
            O => \N__5686\,
            I => \N__5669\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__5679\,
            I => \N__5666\
        );

    \I__745\ : Span4Mux_v
    port map (
            O => \N__5676\,
            I => \N__5659\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5669\,
            I => \N__5659\
        );

    \I__743\ : Span4Mux_h
    port map (
            O => \N__5666\,
            I => \N__5659\
        );

    \I__742\ : Odrv4
    port map (
            O => \N__5659\,
            I => \PCH_PWRGD.N_3_i\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__5656\,
            I => \PCH_PWRGD.delayed_vccin_ok_e_1_cascade_\
        );

    \I__740\ : InMux
    port map (
            O => \N__5653\,
            I => \N__5647\
        );

    \I__739\ : InMux
    port map (
            O => \N__5652\,
            I => \N__5647\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__5647\,
            I => \PCH_PWRGD.delayed_vccin_ok_0\
        );

    \I__737\ : IoInMux
    port map (
            O => \N__5644\,
            I => \N__5641\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__5641\,
            I => \N__5638\
        );

    \I__735\ : IoSpan4Mux
    port map (
            O => \N__5638\,
            I => \N__5635\
        );

    \I__734\ : Span4Mux_s3_h
    port map (
            O => \N__5635\,
            I => \N__5631\
        );

    \I__733\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5628\
        );

    \I__732\ : Span4Mux_h
    port map (
            O => \N__5631\,
            I => \N__5623\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__5628\,
            I => \N__5623\
        );

    \I__730\ : Span4Mux_v
    port map (
            O => \N__5623\,
            I => \N__5620\
        );

    \I__729\ : Span4Mux_h
    port map (
            O => \N__5620\,
            I => \N__5617\
        );

    \I__728\ : Odrv4
    port map (
            O => \N__5617\,
            I => v1p8a_ok
        );

    \I__727\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5611\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5611\,
            I => \N__5608\
        );

    \I__725\ : Span4Mux_v
    port map (
            O => \N__5608\,
            I => \N__5605\
        );

    \I__724\ : Span4Mux_h
    port map (
            O => \N__5605\,
            I => \N__5602\
        );

    \I__723\ : Span4Mux_v
    port map (
            O => \N__5602\,
            I => \N__5599\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__5599\,
            I => v5a_ok
        );

    \I__721\ : IoInMux
    port map (
            O => \N__5596\,
            I => \N__5593\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5593\,
            I => \N__5590\
        );

    \I__719\ : IoSpan4Mux
    port map (
            O => \N__5590\,
            I => \N__5585\
        );

    \I__718\ : IoInMux
    port map (
            O => \N__5589\,
            I => \N__5582\
        );

    \I__717\ : CascadeMux
    port map (
            O => \N__5588\,
            I => \N__5579\
        );

    \I__716\ : IoSpan4Mux
    port map (
            O => \N__5585\,
            I => \N__5574\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5582\,
            I => \N__5574\
        );

    \I__714\ : InMux
    port map (
            O => \N__5579\,
            I => \N__5571\
        );

    \I__713\ : IoSpan4Mux
    port map (
            O => \N__5574\,
            I => \N__5568\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__5571\,
            I => \N__5565\
        );

    \I__711\ : Span4Mux_s1_h
    port map (
            O => \N__5568\,
            I => \N__5562\
        );

    \I__710\ : Span4Mux_v
    port map (
            O => \N__5565\,
            I => \N__5559\
        );

    \I__709\ : Span4Mux_h
    port map (
            O => \N__5562\,
            I => \N__5554\
        );

    \I__708\ : Span4Mux_v
    port map (
            O => \N__5559\,
            I => \N__5554\
        );

    \I__707\ : Span4Mux_h
    port map (
            O => \N__5554\,
            I => \N__5551\
        );

    \I__706\ : Odrv4
    port map (
            O => \N__5551\,
            I => v33a_ok
        );

    \I__705\ : InMux
    port map (
            O => \N__5548\,
            I => \N__5545\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5545\,
            I => \N__5541\
        );

    \I__703\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5538\
        );

    \I__702\ : Span4Mux_h
    port map (
            O => \N__5541\,
            I => \N__5533\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5538\,
            I => \N__5533\
        );

    \I__700\ : Span4Mux_h
    port map (
            O => \N__5533\,
            I => \N__5530\
        );

    \I__699\ : Span4Mux_v
    port map (
            O => \N__5530\,
            I => \N__5527\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__5527\,
            I => slp_susn
        );

    \I__697\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5521\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5521\,
            I => \N__5517\
        );

    \I__695\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5514\
        );

    \I__694\ : Odrv4
    port map (
            O => \N__5517\,
            I => \PCH_PWRGD.count_m2_0_a2_0\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__5514\,
            I => \PCH_PWRGD.count_m2_0_a2_0\
        );

    \I__692\ : InMux
    port map (
            O => \N__5509\,
            I => \N__5506\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__5506\,
            I => \N__5502\
        );

    \I__690\ : InMux
    port map (
            O => \N__5505\,
            I => \N__5499\
        );

    \I__689\ : Span4Mux_v
    port map (
            O => \N__5502\,
            I => \N__5493\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__5499\,
            I => \N__5493\
        );

    \I__687\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5489\
        );

    \I__686\ : Span4Mux_v
    port map (
            O => \N__5493\,
            I => \N__5486\
        );

    \I__685\ : InMux
    port map (
            O => \N__5492\,
            I => \N__5483\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__5489\,
            I => \PCH_PWRGD.N_580_i\
        );

    \I__683\ : Odrv4
    port map (
            O => \N__5486\,
            I => \PCH_PWRGD.N_580_i\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5483\,
            I => \PCH_PWRGD.N_580_i\
        );

    \I__681\ : IoInMux
    port map (
            O => \N__5476\,
            I => \N__5473\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5473\,
            I => \N__5470\
        );

    \I__679\ : IoSpan4Mux
    port map (
            O => \N__5470\,
            I => \N__5464\
        );

    \I__678\ : InMux
    port map (
            O => \N__5469\,
            I => \N__5459\
        );

    \I__677\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5456\
        );

    \I__676\ : CascadeMux
    port map (
            O => \N__5467\,
            I => \N__5452\
        );

    \I__675\ : Span4Mux_s2_v
    port map (
            O => \N__5464\,
            I => \N__5449\
        );

    \I__674\ : InMux
    port map (
            O => \N__5463\,
            I => \N__5446\
        );

    \I__673\ : InMux
    port map (
            O => \N__5462\,
            I => \N__5443\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__5459\,
            I => \N__5438\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__5456\,
            I => \N__5438\
        );

    \I__670\ : CascadeMux
    port map (
            O => \N__5455\,
            I => \N__5435\
        );

    \I__669\ : InMux
    port map (
            O => \N__5452\,
            I => \N__5430\
        );

    \I__668\ : Sp12to4
    port map (
            O => \N__5449\,
            I => \N__5421\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__5446\,
            I => \N__5421\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__5443\,
            I => \N__5421\
        );

    \I__665\ : Sp12to4
    port map (
            O => \N__5438\,
            I => \N__5421\
        );

    \I__664\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5418\
        );

    \I__663\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5415\
        );

    \I__662\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5412\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5430\,
            I => rsmrstn
        );

    \I__660\ : Odrv12
    port map (
            O => \N__5421\,
            I => rsmrstn
        );

    \I__659\ : LocalMux
    port map (
            O => \N__5418\,
            I => rsmrstn
        );

    \I__658\ : LocalMux
    port map (
            O => \N__5415\,
            I => rsmrstn
        );

    \I__657\ : LocalMux
    port map (
            O => \N__5412\,
            I => rsmrstn
        );

    \I__656\ : InMux
    port map (
            O => \N__5401\,
            I => \N__5397\
        );

    \I__655\ : InMux
    port map (
            O => \N__5400\,
            I => \N__5394\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__5397\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__5394\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__652\ : InMux
    port map (
            O => \N__5389\,
            I => \N__5385\
        );

    \I__651\ : InMux
    port map (
            O => \N__5388\,
            I => \N__5382\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__5385\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__5382\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__5377\,
            I => \N__5373\
        );

    \I__647\ : InMux
    port map (
            O => \N__5376\,
            I => \N__5370\
        );

    \I__646\ : InMux
    port map (
            O => \N__5373\,
            I => \N__5367\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__5370\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__5367\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__643\ : InMux
    port map (
            O => \N__5362\,
            I => \N__5358\
        );

    \I__642\ : InMux
    port map (
            O => \N__5361\,
            I => \N__5355\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__5358\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__5355\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__639\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5346\
        );

    \I__638\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5343\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__5346\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__5343\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__635\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5334\
        );

    \I__634\ : InMux
    port map (
            O => \N__5337\,
            I => \N__5331\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__5334\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__5331\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__631\ : CascadeMux
    port map (
            O => \N__5326\,
            I => \N__5322\
        );

    \I__630\ : InMux
    port map (
            O => \N__5325\,
            I => \N__5319\
        );

    \I__629\ : InMux
    port map (
            O => \N__5322\,
            I => \N__5316\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__5319\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__5316\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__626\ : InMux
    port map (
            O => \N__5311\,
            I => \N__5307\
        );

    \I__625\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5304\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__5307\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__5304\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__622\ : InMux
    port map (
            O => \N__5299\,
            I => \N__5295\
        );

    \I__621\ : InMux
    port map (
            O => \N__5298\,
            I => \N__5292\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__5295\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__5292\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__618\ : InMux
    port map (
            O => \N__5287\,
            I => \N__5283\
        );

    \I__617\ : InMux
    port map (
            O => \N__5286\,
            I => \N__5280\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__5283\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__5280\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__5275\,
            I => \N__5272\
        );

    \I__613\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5268\
        );

    \I__612\ : InMux
    port map (
            O => \N__5271\,
            I => \N__5265\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__5268\,
            I => \N__5262\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__5265\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__609\ : Odrv4
    port map (
            O => \N__5262\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__608\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5253\
        );

    \I__607\ : InMux
    port map (
            O => \N__5256\,
            I => \N__5250\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__5253\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__5250\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__604\ : InMux
    port map (
            O => \N__5245\,
            I => \N__5242\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__5242\,
            I => \N__5239\
        );

    \I__602\ : Odrv4
    port map (
            O => \N__5239\,
            I => \VPP_VDDQ.un6_count_11\
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__5236\,
            I => \VPP_VDDQ.un6_count_8_cascade_\
        );

    \I__600\ : InMux
    port map (
            O => \N__5233\,
            I => \N__5230\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__5230\,
            I => \VPP_VDDQ.un6_count_9\
        );

    \I__598\ : InMux
    port map (
            O => \N__5227\,
            I => \N__5223\
        );

    \I__597\ : InMux
    port map (
            O => \N__5226\,
            I => \N__5220\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__5223\,
            I => \N__5215\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__5220\,
            I => \N__5215\
        );

    \I__594\ : Span4Mux_v
    port map (
            O => \N__5215\,
            I => \N__5211\
        );

    \I__593\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5208\
        );

    \I__592\ : Sp12to4
    port map (
            O => \N__5211\,
            I => \N__5203\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__5208\,
            I => \N__5203\
        );

    \I__590\ : Odrv12
    port map (
            O => \N__5203\,
            I => vr_ready_vccin
        );

    \I__589\ : InMux
    port map (
            O => \N__5200\,
            I => \N__5196\
        );

    \I__588\ : InMux
    port map (
            O => \N__5199\,
            I => \N__5193\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__5196\,
            I => \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8PZ0Z7\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__5193\,
            I => \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8PZ0Z7\
        );

    \I__585\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5182\
        );

    \I__584\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5182\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__5182\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__5179\,
            I => \PCH_PWRGD.count_rst_1_cascade_\
        );

    \I__581\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5173\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__5173\,
            I => \PCH_PWRGD.un2_count_1_axb_13\
        );

    \I__579\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5165\
        );

    \I__578\ : InMux
    port map (
            O => \N__5169\,
            I => \N__5162\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__5168\,
            I => \N__5159\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__5165\,
            I => \N__5154\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__5162\,
            I => \N__5154\
        );

    \I__574\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5149\
        );

    \I__573\ : Span4Mux_v
    port map (
            O => \N__5154\,
            I => \N__5146\
        );

    \I__572\ : InMux
    port map (
            O => \N__5153\,
            I => \N__5143\
        );

    \I__571\ : InMux
    port map (
            O => \N__5152\,
            I => \N__5140\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__5149\,
            I => \N__5133\
        );

    \I__569\ : Sp12to4
    port map (
            O => \N__5146\,
            I => \N__5133\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__5143\,
            I => \N__5133\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__5140\,
            I => \N__5130\
        );

    \I__566\ : Span12Mux_s10_h
    port map (
            O => \N__5133\,
            I => \N__5127\
        );

    \I__565\ : Span12Mux_s10_h
    port map (
            O => \N__5130\,
            I => \N__5124\
        );

    \I__564\ : Odrv12
    port map (
            O => \N__5127\,
            I => slp_s3n
        );

    \I__563\ : Odrv12
    port map (
            O => \N__5124\,
            I => slp_s3n
        );

    \I__562\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5115\
        );

    \I__561\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5112\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__5115\,
            I => \PCH_PWRGD.count_rst_0\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__5112\,
            I => \PCH_PWRGD.count_rst_0\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__5107\,
            I => \N__5104\
        );

    \I__557\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5101\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__5101\,
            I => \PCH_PWRGD.count_rst_1\
        );

    \I__555\ : InMux
    port map (
            O => \N__5098\,
            I => \N__5095\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__5095\,
            I => \N__5092\
        );

    \I__553\ : Span4Mux_h
    port map (
            O => \N__5092\,
            I => \N__5089\
        );

    \I__552\ : Odrv4
    port map (
            O => \N__5089\,
            I => \PCH_PWRGD.un2_count_1_cry_9_c_RNIEQ4KZ0Z5\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__5086\,
            I => \tmp_1_RNIBJDJ_cascade_\
        );

    \I__550\ : InMux
    port map (
            O => \N__5083\,
            I => \N__5080\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__5080\,
            I => \PCH_PWRGD.delayed_vccin_okZ0\
        );

    \I__548\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5073\
        );

    \I__547\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5070\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__5073\,
            I => \N__5066\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__5070\,
            I => \N__5063\
        );

    \I__544\ : InMux
    port map (
            O => \N__5069\,
            I => \N__5060\
        );

    \I__543\ : Odrv4
    port map (
            O => \N__5066\,
            I => \N_600_i\
        );

    \I__542\ : Odrv4
    port map (
            O => \N__5063\,
            I => \N_600_i\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__5060\,
            I => \N_600_i\
        );

    \I__540\ : InMux
    port map (
            O => \N__5053\,
            I => \N__5050\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__5050\,
            I => \PCH_PWRGD.delayed_vccin_ok_e_1\
        );

    \I__538\ : InMux
    port map (
            O => \N__5047\,
            I => \PCH_PWRGD.un2_count_1_cry_11\
        );

    \I__537\ : InMux
    port map (
            O => \N__5044\,
            I => \PCH_PWRGD.un2_count_1_cry_12\
        );

    \I__536\ : InMux
    port map (
            O => \N__5041\,
            I => \PCH_PWRGD.un2_count_1_cry_13\
        );

    \I__535\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5034\
        );

    \I__534\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5031\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__5034\,
            I => \N__5028\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__5031\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__5028\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__530\ : InMux
    port map (
            O => \N__5023\,
            I => \PCH_PWRGD.un2_count_1_cry_14\
        );

    \I__529\ : InMux
    port map (
            O => \N__5020\,
            I => \N__5016\
        );

    \I__528\ : InMux
    port map (
            O => \N__5019\,
            I => \N__5013\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__5016\,
            I => \PCH_PWRGD.un2_count_1_cry_14_c_RNICCRZ0Z7\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__5013\,
            I => \PCH_PWRGD.un2_count_1_cry_14_c_RNICCRZ0Z7\
        );

    \I__525\ : InMux
    port map (
            O => \N__5008\,
            I => \N__5005\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__5005\,
            I => \N__5002\
        );

    \I__523\ : Odrv4
    port map (
            O => \N__5002\,
            I => \PCH_PWRGD.count_RNI1N0D1Z0Z_10\
        );

    \I__522\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4996\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4996\,
            I => \PCH_PWRGD.un2_count_1_axb_10\
        );

    \I__520\ : InMux
    port map (
            O => \N__4993\,
            I => \N__4990\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4990\,
            I => \PCH_PWRGD.un2_count_1_axb_14\
        );

    \I__518\ : CascadeMux
    port map (
            O => \N__4987\,
            I => \N__4984\
        );

    \I__517\ : InMux
    port map (
            O => \N__4984\,
            I => \N__4978\
        );

    \I__516\ : InMux
    port map (
            O => \N__4983\,
            I => \N__4978\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4978\,
            I => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\
        );

    \I__514\ : InMux
    port map (
            O => \N__4975\,
            I => \PCH_PWRGD.un2_count_1_cry_2\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__4972\,
            I => \N__4968\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__4971\,
            I => \N__4965\
        );

    \I__511\ : InMux
    port map (
            O => \N__4968\,
            I => \N__4961\
        );

    \I__510\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4956\
        );

    \I__509\ : InMux
    port map (
            O => \N__4964\,
            I => \N__4956\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4961\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__4956\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__506\ : InMux
    port map (
            O => \N__4951\,
            I => \N__4945\
        );

    \I__505\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4945\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__4945\,
            I => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\
        );

    \I__503\ : InMux
    port map (
            O => \N__4942\,
            I => \PCH_PWRGD.un2_count_1_cry_3\
        );

    \I__502\ : InMux
    port map (
            O => \N__4939\,
            I => \PCH_PWRGD.un2_count_1_cry_4\
        );

    \I__501\ : InMux
    port map (
            O => \N__4936\,
            I => \PCH_PWRGD.un2_count_1_cry_5\
        );

    \I__500\ : InMux
    port map (
            O => \N__4933\,
            I => \PCH_PWRGD.un2_count_1_cry_6\
        );

    \I__499\ : InMux
    port map (
            O => \N__4930\,
            I => \PCH_PWRGD.un2_count_1_cry_7\
        );

    \I__498\ : InMux
    port map (
            O => \N__4927\,
            I => \bfn_5_7_0_\
        );

    \I__497\ : InMux
    port map (
            O => \N__4924\,
            I => \PCH_PWRGD.un2_count_1_cry_9\
        );

    \I__496\ : InMux
    port map (
            O => \N__4921\,
            I => \PCH_PWRGD.un2_count_1_cry_10\
        );

    \I__495\ : InMux
    port map (
            O => \N__4918\,
            I => \N__4915\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4915\,
            I => \PCH_PWRGD.un12_clk_100khz_9\
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__4912\,
            I => \PCH_PWRGD.count_rst_10_cascade_\
        );

    \I__492\ : CascadeMux
    port map (
            O => \N__4909\,
            I => \PCH_PWRGD.countZ0Z_4_cascade_\
        );

    \I__491\ : InMux
    port map (
            O => \N__4906\,
            I => \N__4903\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4903\,
            I => \PCH_PWRGD.count_0_4\
        );

    \I__489\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4897\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4897\,
            I => \PCH_PWRGD.count_0_5\
        );

    \I__487\ : InMux
    port map (
            O => \N__4894\,
            I => \N__4889\
        );

    \I__486\ : InMux
    port map (
            O => \N__4893\,
            I => \N__4886\
        );

    \I__485\ : InMux
    port map (
            O => \N__4892\,
            I => \N__4883\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4889\,
            I => \PCH_PWRGD.un2_count_1_axb_1\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__4886\,
            I => \PCH_PWRGD.un2_count_1_axb_1\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4883\,
            I => \PCH_PWRGD.un2_count_1_axb_1\
        );

    \I__481\ : InMux
    port map (
            O => \N__4876\,
            I => \N__4870\
        );

    \I__480\ : InMux
    port map (
            O => \N__4875\,
            I => \N__4867\
        );

    \I__479\ : CascadeMux
    port map (
            O => \N__4874\,
            I => \N__4863\
        );

    \I__478\ : InMux
    port map (
            O => \N__4873\,
            I => \N__4860\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4870\,
            I => \N__4855\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4867\,
            I => \N__4855\
        );

    \I__475\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4852\
        );

    \I__474\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4849\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__4860\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__472\ : Odrv4
    port map (
            O => \N__4855\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4852\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4849\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__469\ : InMux
    port map (
            O => \N__4840\,
            I => \PCH_PWRGD.un2_count_1_cry_1\
        );

    \I__468\ : InMux
    port map (
            O => \N__4837\,
            I => \VPP_VDDQ.un1_count_1_cry_10\
        );

    \I__467\ : InMux
    port map (
            O => \N__4834\,
            I => \VPP_VDDQ.un1_count_1_cry_11\
        );

    \I__466\ : InMux
    port map (
            O => \N__4831\,
            I => \VPP_VDDQ.un1_count_1_cry_12\
        );

    \I__465\ : InMux
    port map (
            O => \N__4828\,
            I => \VPP_VDDQ.un1_count_1_cry_13\
        );

    \I__464\ : InMux
    port map (
            O => \N__4825\,
            I => \bfn_4_12_0_\
        );

    \I__463\ : IoInMux
    port map (
            O => \N__4822\,
            I => \N__4819\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4819\,
            I => \N__4815\
        );

    \I__461\ : IoInMux
    port map (
            O => \N__4818\,
            I => \N__4812\
        );

    \I__460\ : Span4Mux_s3_h
    port map (
            O => \N__4815\,
            I => \N__4809\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__4812\,
            I => \N__4806\
        );

    \I__458\ : Sp12to4
    port map (
            O => \N__4809\,
            I => \N__4801\
        );

    \I__457\ : Span12Mux_s3_h
    port map (
            O => \N__4806\,
            I => \N__4801\
        );

    \I__456\ : Odrv12
    port map (
            O => \N__4801\,
            I => v5s_enn
        );

    \I__455\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4795\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__4795\,
            I => slp_s4n
        );

    \I__453\ : InMux
    port map (
            O => \N__4792\,
            I => \VPP_VDDQ.un1_count_1_cry_1\
        );

    \I__452\ : InMux
    port map (
            O => \N__4789\,
            I => \VPP_VDDQ.un1_count_1_cry_2\
        );

    \I__451\ : InMux
    port map (
            O => \N__4786\,
            I => \VPP_VDDQ.un1_count_1_cry_3\
        );

    \I__450\ : InMux
    port map (
            O => \N__4783\,
            I => \VPP_VDDQ.un1_count_1_cry_4\
        );

    \I__449\ : InMux
    port map (
            O => \N__4780\,
            I => \VPP_VDDQ.un1_count_1_cry_5\
        );

    \I__448\ : InMux
    port map (
            O => \N__4777\,
            I => \VPP_VDDQ.un1_count_1_cry_6\
        );

    \I__447\ : InMux
    port map (
            O => \N__4774\,
            I => \bfn_4_11_0_\
        );

    \I__446\ : InMux
    port map (
            O => \N__4771\,
            I => \VPP_VDDQ.un1_count_1_cry_8\
        );

    \I__445\ : InMux
    port map (
            O => \N__4768\,
            I => \VPP_VDDQ.un1_count_1_cry_9\
        );

    \I__444\ : InMux
    port map (
            O => \N__4765\,
            I => \N__4762\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4762\,
            I => \N__4759\
        );

    \I__442\ : Odrv4
    port map (
            O => \N__4759\,
            I => \PCH_PWRGD.count_0_0\
        );

    \I__441\ : InMux
    port map (
            O => \N__4756\,
            I => \N__4753\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4753\,
            I => \PCH_PWRGD.count_rst_14\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__4750\,
            I => \PCH_PWRGD.countZ0Z_0_cascade_\
        );

    \I__438\ : InMux
    port map (
            O => \N__4747\,
            I => \N__4744\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__4744\,
            I => \N__4741\
        );

    \I__436\ : Span4Mux_v
    port map (
            O => \N__4741\,
            I => \N__4738\
        );

    \I__435\ : Odrv4
    port map (
            O => \N__4738\,
            I => \PCH_PWRGD.count_rst_13\
        );

    \I__434\ : CascadeMux
    port map (
            O => \N__4735\,
            I => \PCH_PWRGD.count_rst_13_cascade_\
        );

    \I__433\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4729\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__4729\,
            I => \N__4725\
        );

    \I__431\ : InMux
    port map (
            O => \N__4728\,
            I => \N__4722\
        );

    \I__430\ : Odrv12
    port map (
            O => \N__4725\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4722\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__428\ : InMux
    port map (
            O => \N__4717\,
            I => \VPP_VDDQ.un1_count_1_cry_0\
        );

    \I__427\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4711\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__4711\,
            I => \N__4708\
        );

    \I__425\ : Odrv4
    port map (
            O => \N__4708\,
            I => \PCH_PWRGD.curr_state_e_0Z0Z_0\
        );

    \I__424\ : CascadeMux
    port map (
            O => \N__4705\,
            I => \PCH_PWRGD.m4_cascade_\
        );

    \I__423\ : CascadeMux
    port map (
            O => \N__4702\,
            I => \PCH_PWRGD.curr_stateZ0Z_0_cascade_\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__4699\,
            I => \PCH_PWRGD.N_580_i_cascade_\
        );

    \I__421\ : CascadeMux
    port map (
            O => \N__4696\,
            I => \PCH_PWRGD.curr_state_7_1_cascade_\
        );

    \I__420\ : InMux
    port map (
            O => \N__4693\,
            I => \N__4690\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__4690\,
            I => \PCH_PWRGD.curr_state_e_0Z0Z_1\
        );

    \I__418\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4684\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__4684\,
            I => \N__4678\
        );

    \I__416\ : InMux
    port map (
            O => \N__4683\,
            I => \N__4671\
        );

    \I__415\ : InMux
    port map (
            O => \N__4682\,
            I => \N__4671\
        );

    \I__414\ : InMux
    port map (
            O => \N__4681\,
            I => \N__4671\
        );

    \I__413\ : Odrv12
    port map (
            O => \N__4678\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__4671\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__4666\,
            I => \PCH_PWRGD.curr_stateZ0Z_1_cascade_\
        );

    \I__410\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4660\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__4660\,
            I => \PCH_PWRGD.count_0_15\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__4657\,
            I => \PCH_PWRGD.count_0_sqmuxa_cascade_\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__4654\,
            I => \PCH_PWRGD.un12_clk_100khz_12_1_cascade_\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__4651\,
            I => \PCH_PWRGD.un12_clk_100khz_1_cascade_\
        );

    \I__405\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4645\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4645\,
            I => \PCH_PWRGD.un12_clk_100khz_1_0\
        );

    \I__403\ : CascadeMux
    port map (
            O => \N__4642\,
            I => \PCH_PWRGD.un12_clk_100khz_5_1_cascade_\
        );

    \I__402\ : InMux
    port map (
            O => \N__4639\,
            I => \N__4636\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__4636\,
            I => \PCH_PWRGD.un12_clk_100khz_5\
        );

    \I__400\ : IoInMux
    port map (
            O => \N__4633\,
            I => \N__4630\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__4630\,
            I => v33a_enn
        );

    \I__398\ : InMux
    port map (
            O => \N__4627\,
            I => \N__4624\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__4624\,
            I => \N__4621\
        );

    \I__396\ : Span4Mux_s3_v
    port map (
            O => \N__4621\,
            I => \N__4618\
        );

    \I__395\ : Odrv4
    port map (
            O => \N__4618\,
            I => vpp_ok
        );

    \I__394\ : IoInMux
    port map (
            O => \N__4615\,
            I => \N__4612\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__4612\,
            I => vddq_en
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_2_1_cry_8_cZ0\,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_5_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_6_0_\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un2_count_1_cry_8\,
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER_un4_counter_7\,
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_8\,
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_16\,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_24\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_4_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_10_0_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_7\,
            carryinitout => \bfn_4_11_0_\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_9_7_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \SLP_SUSn_RNIN4K9_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5548\,
            lcout => v33a_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_vddq_en_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4627\,
            in2 => \_gnd_net_\,
            in3 => \N__5969\,
            lcout => vddq_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_e_0_0_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__6306\,
            in1 => \N__6468\,
            in2 => \N__5704\,
            in3 => \N__4687\,
            lcout => \PCH_PWRGD.curr_state_e_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10411\,
            ce => \N__9447\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4875\,
            in1 => \N__7190\,
            in2 => \_gnd_net_\,
            in3 => \N__6450\,
            lcout => \PCH_PWRGD.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10495\,
            ce => \N__6960\,
            sr => \N__6788\
        );

    \PCH_PWRGD.count_RNI_8_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4918\,
            in1 => \N__6559\,
            in2 => \N__6526\,
            in3 => \N__6172\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un12_clk_100khz_12_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI21JO2_0_1_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__6963\,
            in1 => \N__4732\,
            in2 => \N__4654\,
            in3 => \N__4747\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un12_clk_100khz_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNINULCI_1_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__4876\,
            in1 => \N__4639\,
            in2 => \N__4651\,
            in3 => \N__4648\,
            lcout => \PCH_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIJ10N9_10_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100011"
        )
    port map (
            in0 => \N__5098\,
            in1 => \N__5008\,
            in2 => \N__6964\,
            in3 => \N__5038\,
            lcout => \PCH_PWRGD.un12_clk_100khz_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI28H5_2_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6337\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5842\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un12_clk_100khz_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI2S2T5_2_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__6352\,
            in1 => \N__5860\,
            in2 => \N__4642\,
            in3 => \N__6936\,
            lcout => \PCH_PWRGD.un12_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_e_0_1_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110000001000"
        )
    port map (
            in0 => \N__4682\,
            in1 => \N__5498\,
            in2 => \N__6476\,
            in3 => \N__5698\,
            lcout => \PCH_PWRGD.curr_state_e_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10496\,
            ce => \N__9446\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m4_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__6433\,
            in1 => \N__6301\,
            in2 => \N__5703\,
            in3 => \N__4681\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.m4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_e_0_RNI7LVE1_0_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4714\,
            in2 => \N__4705\,
            in3 => \N__8498\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_0\,
            ltout => \PCH_PWRGD.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_e_0_RNI_0_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4702\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.N_580_i\,
            ltout => \PCH_PWRGD.N_580_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m6_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011100000"
        )
    port map (
            in0 => \N__4683\,
            in1 => \N__5694\,
            in2 => \N__4699\,
            in3 => \N__6432\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.curr_state_7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_e_0_RNI8MVE1_1_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__8497\,
            in1 => \_gnd_net_\,
            in2 => \N__4696\,
            in3 => \N__4693\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_1\,
            ltout => \PCH_PWRGD.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_e_0_RNI_1_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4666\,
            in3 => \_gnd_net_\,
            lcout => \N_600_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI76RC4_15_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__6942\,
            in1 => \N__5019\,
            in2 => \N__7193\,
            in3 => \N__4663\,
            lcout => \PCH_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_15_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5020\,
            lcout => \PCH_PWRGD.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10626\,
            ce => \N__6973\,
            sr => \N__6767\
        );

    \PCH_PWRGD.curr_state_e_0_RNI41T31_0_0_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5520\,
            in1 => \N__5492\,
            in2 => \N__5455\,
            in3 => \N__8480\,
            lcout => \PCH_PWRGD.count_0_sqmuxa\,
            ltout => \PCH_PWRGD.count_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI41T31_0_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__4873\,
            in1 => \_gnd_net_\,
            in2 => \N__4657\,
            in3 => \N__6456\,
            lcout => \PCH_PWRGD.count_rst_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI51GS3_0_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4765\,
            in1 => \N__4756\,
            in2 => \_gnd_net_\,
            in3 => \N__6940\,
            lcout => \PCH_PWRGD.countZ0Z_0\,
            ltout => \PCH_PWRGD.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI62GS3_1_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4894\,
            in2 => \N__4750\,
            in3 => \N__7133\,
            lcout => \PCH_PWRGD.count_rst_13\,
            ltout => \PCH_PWRGD.count_rst_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI21JO2_1_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4728\,
            in2 => \N__4735\,
            in3 => \N__6941\,
            lcout => \PCH_PWRGD.un2_count_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_13_c_RNIFBNB1_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__7050\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7159\,
            lcout => \PCH_PWRGD.count_rst_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_13_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5199\,
            in2 => \_gnd_net_\,
            in3 => \N__7155\,
            lcout => \PCH_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10572\,
            ce => \N__6961\,
            sr => \N__6787\
        );

    \PCH_PWRGD.count_1_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7154\,
            in1 => \N__4866\,
            in2 => \_gnd_net_\,
            in3 => \N__4893\,
            lcout => \PCH_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10572\,
            ce => \N__6961\,
            sr => \N__6787\
        );

    \PCH_PWRGD_PCH_PWRGD_un1_count_1_sqmuxa_0_0_a3_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5214\,
            in1 => \N__5434\,
            in2 => \N__5168\,
            in3 => \N__5076\,
            lcout => \PCH_PWRGD_N_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_0_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9029\,
            in1 => \N__5767\,
            in2 => \N__5749\,
            in3 => \N__5748\,
            lcout => \VPP_VDDQ.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_10_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_0\,
            clk => \N__10609\,
            ce => 'H',
            sr => \N__6117\
        );

    \VPP_VDDQ.count_1_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9025\,
            in1 => \N__5311\,
            in2 => \_gnd_net_\,
            in3 => \N__4717\,
            lcout => \VPP_VDDQ.countZ0Z_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_0\,
            carryout => \VPP_VDDQ.un1_count_1_cry_1\,
            clk => \N__10609\,
            ce => 'H',
            sr => \N__6117\
        );

    \VPP_VDDQ.count_2_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9030\,
            in1 => \N__5338\,
            in2 => \_gnd_net_\,
            in3 => \N__4792\,
            lcout => \VPP_VDDQ.countZ0Z_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_1_cry_2\,
            clk => \N__10609\,
            ce => 'H',
            sr => \N__6117\
        );

    \VPP_VDDQ.count_3_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9026\,
            in1 => \N__5401\,
            in2 => \_gnd_net_\,
            in3 => \N__4789\,
            lcout => \VPP_VDDQ.countZ0Z_3\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_1_cry_3\,
            clk => \N__10609\,
            ce => 'H',
            sr => \N__6117\
        );

    \VPP_VDDQ.count_4_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9031\,
            in1 => \N__5362\,
            in2 => \_gnd_net_\,
            in3 => \N__4786\,
            lcout => \VPP_VDDQ.countZ0Z_4\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_1_cry_4\,
            clk => \N__10609\,
            ce => 'H',
            sr => \N__6117\
        );

    \VPP_VDDQ.count_5_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9027\,
            in1 => \N__5389\,
            in2 => \_gnd_net_\,
            in3 => \N__4783\,
            lcout => \VPP_VDDQ.countZ0Z_5\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_1_cry_5\,
            clk => \N__10609\,
            ce => 'H',
            sr => \N__6117\
        );

    \VPP_VDDQ.count_6_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9032\,
            in1 => \N__5350\,
            in2 => \_gnd_net_\,
            in3 => \N__4780\,
            lcout => \VPP_VDDQ.countZ0Z_6\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_1_cry_6\,
            clk => \N__10609\,
            ce => 'H',
            sr => \N__6117\
        );

    \VPP_VDDQ.count_7_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9028\,
            in1 => \N__5376\,
            in2 => \_gnd_net_\,
            in3 => \N__4777\,
            lcout => \VPP_VDDQ.countZ0Z_7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_1_cry_7\,
            clk => \N__10609\,
            ce => 'H',
            sr => \N__6117\
        );

    \VPP_VDDQ.count_8_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9090\,
            in1 => \N__5796\,
            in2 => \_gnd_net_\,
            in3 => \N__4774\,
            lcout => \VPP_VDDQ.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_4_11_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_8\,
            clk => \N__10633\,
            ce => 'H',
            sr => \N__6110\
        );

    \VPP_VDDQ.count_9_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9086\,
            in1 => \N__5812\,
            in2 => \_gnd_net_\,
            in3 => \N__4771\,
            lcout => \VPP_VDDQ.countZ0Z_9\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_8\,
            carryout => \VPP_VDDQ.un1_count_1_cry_9\,
            clk => \N__10633\,
            ce => 'H',
            sr => \N__6110\
        );

    \VPP_VDDQ.count_10_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9087\,
            in1 => \N__5325\,
            in2 => \_gnd_net_\,
            in3 => \N__4768\,
            lcout => \VPP_VDDQ.countZ0Z_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_1_cry_10\,
            clk => \N__10633\,
            ce => 'H',
            sr => \N__6110\
        );

    \VPP_VDDQ.count_11_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9084\,
            in1 => \N__5781\,
            in2 => \_gnd_net_\,
            in3 => \N__4837\,
            lcout => \VPP_VDDQ.countZ0Z_11\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_1_cry_11\,
            clk => \N__10633\,
            ce => 'H',
            sr => \N__6110\
        );

    \VPP_VDDQ.count_12_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9088\,
            in1 => \N__5287\,
            in2 => \_gnd_net_\,
            in3 => \N__4834\,
            lcout => \VPP_VDDQ.countZ0Z_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_1_cry_12\,
            clk => \N__10633\,
            ce => 'H',
            sr => \N__6110\
        );

    \VPP_VDDQ.count_13_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9085\,
            in1 => \N__5271\,
            in2 => \_gnd_net_\,
            in3 => \N__4831\,
            lcout => \VPP_VDDQ.countZ0Z_13\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_1_cry_13\,
            clk => \N__10633\,
            ce => 'H',
            sr => \N__6110\
        );

    \VPP_VDDQ.count_14_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9089\,
            in1 => \N__5299\,
            in2 => \_gnd_net_\,
            in3 => \N__4828\,
            lcout => \VPP_VDDQ.countZ0Z_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14\,
            clk => \N__10633\,
            ce => 'H',
            sr => \N__6110\
        );

    \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10114\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_14\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_15_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5257\,
            in2 => \_gnd_net_\,
            in3 => \N__4825\,
            lcout => \VPP_VDDQ.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10617\,
            ce => \N__6082\,
            sr => \N__6118\
        );

    \VPP_VDDQ.slp_s3n_signal_i_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5152\,
            lcout => v5s_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.VCCST_EN_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5468\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4798\,
            lcout => vccst_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_7_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__6613\,
            in1 => \N__7192\,
            in2 => \N__6139\,
            in3 => \N__6455\,
            lcout => \PCH_PWRGD.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10494\,
            ce => \N__6972\,
            sr => \N__6786\
        );

    \PCH_PWRGD.count_5_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__6202\,
            in1 => \N__7191\,
            in2 => \N__6229\,
            in3 => \N__6454\,
            lcout => \PCH_PWRGD.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10494\,
            ce => \N__6972\,
            sr => \N__6786\
        );

    \PCH_PWRGD.count_RNI_3_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6203\,
            in1 => \N__4964\,
            in2 => \N__6256\,
            in3 => \N__6612\,
            lcout => \PCH_PWRGD.un12_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_c_RNITFQG1_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__6249\,
            in1 => \N__7189\,
            in2 => \N__4987\,
            in3 => \N__6449\,
            lcout => \PCH_PWRGD.count_rst_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_3_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__6447\,
            in1 => \N__6248\,
            in2 => \N__7201\,
            in3 => \N__4983\,
            lcout => \PCH_PWRGD.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10597\,
            ce => \N__6968\,
            sr => \N__6790\
        );

    \PCH_PWRGD.un2_count_1_cry_3_c_RNIUHRG1_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__4950\,
            in1 => \N__7184\,
            in2 => \N__4971\,
            in3 => \N__6446\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI3ME94_4_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__6887\,
            in1 => \_gnd_net_\,
            in2 => \N__4912\,
            in3 => \N__4906\,
            lcout => \PCH_PWRGD.countZ0Z_4\,
            ltout => \PCH_PWRGD.countZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_4_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__4951\,
            in1 => \N__7185\,
            in2 => \N__4909\,
            in3 => \N__6448\,
            lcout => \PCH_PWRGD.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10597\,
            ce => \N__6968\,
            sr => \N__6790\
        );

    \PCH_PWRGD.count_RNI5PF94_5_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4900\,
            in1 => \N__6181\,
            in2 => \_gnd_net_\,
            in3 => \N__6886\,
            lcout => \PCH_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4892\,
            in2 => \N__4874\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_6_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_RNISDPG1_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7135\,
            in1 => \N__5827\,
            in2 => \_gnd_net_\,
            in3 => \N__4840\,
            lcout => \PCH_PWRGD.count_rst_12\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_1\,
            carryout => \PCH_PWRGD.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6247\,
            in2 => \_gnd_net_\,
            in3 => \N__4975\,
            lcout => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_2\,
            carryout => \PCH_PWRGD.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4972\,
            in3 => \N__4942\,
            lcout => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_3\,
            carryout => \PCH_PWRGD.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6210\,
            in3 => \N__4939\,
            lcout => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_4\,
            carryout => \PCH_PWRGD.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_5_c_RNI0MTG1_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7136\,
            in1 => \N__5866\,
            in2 => \_gnd_net_\,
            in3 => \N__4936\,
            lcout => \PCH_PWRGD.count_rst_8\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_5\,
            carryout => \PCH_PWRGD.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6611\,
            in2 => \_gnd_net_\,
            in3 => \N__4933\,
            lcout => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_6\,
            carryout => \PCH_PWRGD.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6552\,
            in2 => \_gnd_net_\,
            in3 => \N__4930\,
            lcout => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_7\,
            carryout => \PCH_PWRGD.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6515\,
            in2 => \_gnd_net_\,
            in3 => \N__4927\,
            lcout => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_5_7_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_9_c_RNI4U1H1_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7183\,
            in1 => \N__4999\,
            in2 => \_gnd_net_\,
            in3 => \N__4924\,
            lcout => \PCH_PWRGD.count_rst_4\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_9\,
            carryout => \PCH_PWRGD.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_10_c_RNI84N7_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6165\,
            in2 => \_gnd_net_\,
            in3 => \N__4921\,
            lcout => \PCH_PWRGD.un2_count_1_cry_10_c_RNI84NZ0Z7\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_10\,
            carryout => \PCH_PWRGD.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_11_c_RNI96O7_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6358\,
            in2 => \_gnd_net_\,
            in3 => \N__5047\,
            lcout => \PCH_PWRGD.un2_count_1_cry_11_c_RNI96OZ0Z7\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_11\,
            carryout => \PCH_PWRGD.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8P7_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5176\,
            in2 => \_gnd_net_\,
            in3 => \N__5044\,
            lcout => \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8PZ0Z7\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_12\,
            carryout => \PCH_PWRGD.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4993\,
            in2 => \_gnd_net_\,
            in3 => \N__5041\,
            lcout => \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_13\,
            carryout => \PCH_PWRGD.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_14_c_RNICCR7_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5037\,
            in2 => \_gnd_net_\,
            in3 => \N__5023\,
            lcout => \PCH_PWRGD.un2_count_1_cry_14_c_RNICCRZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_e_0_RNIG9DT_1_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5227\,
            in1 => \N__5170\,
            in2 => \_gnd_net_\,
            in3 => \N__5069\,
            lcout => \PCH_PWRGD.count_m2_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI1N0D1_10_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6636\,
            in1 => \N__5187\,
            in2 => \N__6991\,
            in3 => \N__7032\,
            lcout => \PCH_PWRGD.count_RNI1N0D1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIMH4I4_10_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__6916\,
            in1 => \N__6990\,
            in2 => \N__7017\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.un2_count_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_1_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__7213\,
            in1 => \N__9033\,
            in2 => \N__5467\,
            in3 => \N__8096\,
            lcout => rsmrstn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI53QC4_14_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__6915\,
            in1 => \_gnd_net_\,
            in2 => \N__7036\,
            in3 => \N__5118\,
            lcout => \PCH_PWRGD.un2_count_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_vccin_ok_1_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5226\,
            in1 => \N__5169\,
            in2 => \_gnd_net_\,
            in3 => \N__5433\,
            lcout => \PCH_PWRGD.N_3_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_12_c_RNIE9MB1_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7160\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5200\,
            lcout => \PCH_PWRGD.count_rst_1\,
            ltout => \PCH_PWRGD.count_rst_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI30PC4_13_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5188\,
            in2 => \N__5179\,
            in3 => \N__6917\,
            lcout => \PCH_PWRGD.un2_count_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8481\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8587\,
            lcout => \clk_100Khz_signalkeep\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10571\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNIBDBV2_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5463\,
            in1 => \N__5083\,
            in2 => \_gnd_net_\,
            in3 => \N__5153\,
            lcout => pch_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_9_c_RNIEQ4K5_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6370\,
            in1 => \N__5119\,
            in2 => \N__5107\,
            in3 => \N__7018\,
            lcout => \PCH_PWRGD.un2_count_1_cry_9_c_RNIEQ4KZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_RNIBJDJ_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8567\,
            in2 => \_gnd_net_\,
            in3 => \N__8474\,
            lcout => \tmp_1_RNIBJDJ\,
            ltout => \tmp_1_RNIBJDJ_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNI45EG2_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000101010"
        )
    port map (
            in0 => \N__5653\,
            in1 => \N__5053\,
            in2 => \N__5086\,
            in3 => \N__5690\,
            lcout => \PCH_PWRGD.delayed_vccin_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_e_0_RNILRFU_0_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101111111"
        )
    port map (
            in0 => \N__6305\,
            in1 => \N__5077\,
            in2 => \N__5699\,
            in3 => \N__5509\,
            lcout => \PCH_PWRGD.delayed_vccin_ok_e_1\,
            ltout => \PCH_PWRGD.delayed_vccin_ok_e_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111010101010"
        )
    port map (
            in0 => \N__5652\,
            in1 => \N__5689\,
            in2 => \N__5656\,
            in3 => \N__9419\,
            lcout => \PCH_PWRGD.delayed_vccin_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10627\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5634\,
            in1 => \N__5614\,
            in2 => \N__5588\,
            in3 => \N__5544\,
            lcout => \RSMRST_PWRGD.N_3_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_e_0_RNI41T31_0_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5524\,
            in1 => \N__5505\,
            in2 => \N__8503\,
            in3 => \N__5462\,
            lcout => \PCH_PWRGD.count_m2_0_a2_iso\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIVJP51_3_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5400\,
            in1 => \N__5388\,
            in2 => \N__5377\,
            in3 => \N__5361\,
            lcout => \VPP_VDDQ.un6_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI63141_10_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5349\,
            in1 => \N__5337\,
            in2 => \N__5326\,
            in3 => \N__5310\,
            lcout => \VPP_VDDQ.un6_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNI7CQO_15_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5298\,
            in1 => \N__5286\,
            in2 => \N__5275\,
            in3 => \N__5256\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un6_count_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNIRFM64_15_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5245\,
            in1 => \N__5755\,
            in2 => \N__5236\,
            in3 => \N__5233\,
            lcout => \VPP_VDDQ_un6_count\,
            ltout => \VPP_VDDQ_un6_count_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.G_24_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__5818\,
            in1 => \N__5724\,
            in2 => \N__5821\,
            in3 => \N__8949\,
            lcout => \G_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNID2IU_0_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__6059\,
            in1 => \_gnd_net_\,
            in2 => \N__6040\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ_curr_state12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFC141_11_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5811\,
            in1 => \N__5797\,
            in2 => \N__5782\,
            in3 => \N__5766\,
            lcout => \VPP_VDDQ.un6_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNIT4VK1_0_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101011111010"
        )
    port map (
            in0 => \N__6034\,
            in1 => \N__9612\,
            in2 => \N__6069\,
            in3 => \N__5973\,
            lcout => \VPP_VDDQ.un1_curr_state13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_1_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110100000"
        )
    port map (
            in0 => \N__8950\,
            in1 => \N__5734\,
            in2 => \N__5728\,
            in3 => \N__6035\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__6067\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6038\,
            lcout => \VPP_VDDQ.curr_state11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNIT4VK1_0_0_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6036\,
            in1 => \N__6063\,
            in2 => \_gnd_net_\,
            in3 => \N__6001\,
            lcout => \VPP_VDDQ_delayed_vddq_pwrgd_1_sqmuxa\,
            ltout => \VPP_VDDQ_delayed_vddq_pwrgd_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011001110"
        )
    port map (
            in0 => \N__9020\,
            in1 => \N__5988\,
            in2 => \N__5716\,
            in3 => \N__6010\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5713\,
            in1 => \N__6004\,
            in2 => \N__5707\,
            in3 => \N__9021\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10616\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNO_0_15_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9019\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6100\,
            lcout => \VPP_VDDQ.N_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_0_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__6039\,
            in1 => \N__6068\,
            in2 => \N__9103\,
            in3 => \N__6003\,
            lcout => \VPP_VDDQ.curr_stateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10616\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_2_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110101"
        )
    port map (
            in0 => \N__6002\,
            in1 => \_gnd_net_\,
            in2 => \N__6070\,
            in3 => \N__6037\,
            lcout => \VPP_VDDQ.un1_curr_state12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_vddq_pwrgd_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9602\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5964\,
            lcout => \VPP_VDDQ.un1_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNI32MH_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5989\,
            in2 => \_gnd_net_\,
            in3 => \N__5965\,
            lcout => vpp_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNIVKCF4_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8218\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5909\,
            lcout => vccst_pwrgd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI7SG94_6_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5856\,
            in1 => \N__5838\,
            in2 => \_gnd_net_\,
            in3 => \N__6881\,
            lcout => \PCH_PWRGD.un2_count_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_6_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5855\,
            lcout => \PCH_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10450\,
            ce => \N__6965\,
            sr => \N__6791\
        );

    \PCH_PWRGD.count_RNIVFC94_2_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6350\,
            in1 => \N__6333\,
            in2 => \_gnd_net_\,
            in3 => \N__6882\,
            lcout => \PCH_PWRGD.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_2_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6351\,
            lcout => \PCH_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10450\,
            ce => \N__6965\,
            sr => \N__6791\
        );

    \PCH_PWRGD.curr_state_e_0_RNI4GQL2_0_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000100"
        )
    port map (
            in0 => \N__6322\,
            in1 => \N__9444\,
            in2 => \N__6310\,
            in3 => \N__7194\,
            lcout => \PCH_PWRGD.curr_state_e_0_RNI4GQL2Z0Z_0\,
            ltout => \PCH_PWRGD.curr_state_e_0_RNI4GQL2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI1JD94_3_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__6271\,
            in1 => \_gnd_net_\,
            in2 => \N__6265\,
            in3 => \N__6262\,
            lcout => \PCH_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_c_RNIVJSG1_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__6478\,
            in1 => \N__6222\,
            in2 => \N__6211\,
            in3 => \N__7196\,
            lcout => \PCH_PWRGD.count_rst_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_10_c_RNIC5KB1_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__7195\,
            in1 => \N__6154\,
            in2 => \_gnd_net_\,
            in3 => \N__6477\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIVPMC4_11_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6145\,
            in2 => \N__6175\,
            in3 => \N__6879\,
            lcout => \PCH_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_11_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__7198\,
            in1 => \N__6153\,
            in2 => \_gnd_net_\,
            in3 => \N__6480\,
            lcout => \PCH_PWRGD.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10455\,
            ce => \N__6932\,
            sr => \N__6792\
        );

    \PCH_PWRGD.un2_count_1_cry_6_c_RNI1OUG1_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__6479\,
            in1 => \N__6610\,
            in2 => \N__6135\,
            in3 => \N__7197\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI9VH94_7_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__6880\,
            in1 => \_gnd_net_\,
            in2 => \N__6625\,
            in3 => \N__6622\,
            lcout => \PCH_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_8_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__7199\,
            in1 => \N__6550\,
            in2 => \N__6586\,
            in3 => \N__6481\,
            lcout => \PCH_PWRGD.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10455\,
            ce => \N__6932\,
            sr => \N__6792\
        );

    \PCH_PWRGD.un2_count_1_cry_7_c_RNI2QVG1_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__7179\,
            in1 => \N__6551\,
            in2 => \N__6585\,
            in3 => \N__6482\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIB2J94_8_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__6919\,
            in1 => \_gnd_net_\,
            in2 => \N__6568\,
            in3 => \N__6565\,
            lcout => \PCH_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_c_RNI3S0H1_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__7180\,
            in1 => \N__6495\,
            in2 => \N__6519\,
            in3 => \N__6483\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNID5K94_9_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6967\,
            in2 => \N__6529\,
            in3 => \N__6379\,
            lcout => \PCH_PWRGD.countZ0Z_9\,
            ltout => \PCH_PWRGD.countZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_9_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__7181\,
            in1 => \N__6496\,
            in2 => \N__6487\,
            in3 => \N__6484\,
            lcout => \PCH_PWRGD.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10545\,
            ce => \N__6966\,
            sr => \N__6789\
        );

    \PCH_PWRGD.un2_count_1_cry_11_c_RNID7LB1_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6646\,
            in2 => \_gnd_net_\,
            in3 => \N__7178\,
            lcout => \PCH_PWRGD.count_rst_2\,
            ltout => \PCH_PWRGD.count_rst_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI1TNC4_12_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6637\,
            in2 => \N__6361\,
            in3 => \N__6918\,
            lcout => \PCH_PWRGD.un2_count_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_12_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6645\,
            in2 => \_gnd_net_\,
            in3 => \N__7182\,
            lcout => \PCH_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10545\,
            ce => \N__6966\,
            sr => \N__6789\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIMO1Q2_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__8166\,
            in1 => \N__8586\,
            in2 => \N__7323\,
            in3 => \N__8332\,
            lcout => \VPP_VDDQ.g0_3_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIR9731_0_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__10841\,
            in1 => \N__11054\,
            in2 => \_gnd_net_\,
            in3 => \N__8165\,
            lcout => \VPP_VDDQ.count_2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_6_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10842\,
            in2 => \N__11099\,
            in3 => \N__8281\,
            lcout => \VPP_VDDQ.count_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10550\,
            ce => \N__10278\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_4_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__8167\,
            in1 => \N__11055\,
            in2 => \N__10852\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10550\,
            ce => \N__10278\,
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6664\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => \COUNTER.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6655\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_0\,
            carryout => \COUNTER.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6706\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_1\,
            carryout => \COUNTER.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6694\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_2\,
            carryout => \COUNTER.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6682\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_3\,
            carryout => \COUNTER.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7252\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_4\,
            carryout => \COUNTER.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7225\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_5\,
            carryout => \COUNTER.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7240\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_6\,
            carryout => \COUNTER_un4_counter_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER_un4_counter_7_THRU_LUT4_0_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6670\,
            lcout => \COUNTER_un4_counter_7_THRU_CO\,
            ltout => \COUNTER_un4_counter_7_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_3_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000000110"
        )
    port map (
            in0 => \N__7575\,
            in1 => \N__7561\,
            in2 => \N__6667\,
            in3 => \_gnd_net_\,
            lcout => \COUNTER.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10554\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_RNIBJDJ_0_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8568\,
            in2 => \_gnd_net_\,
            in3 => \N__8496\,
            lcout => \tmp_1_RNIBJDJ_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_RNO_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7574\,
            in1 => \N__7618\,
            in2 => \N__7552\,
            in3 => \N__7601\,
            lcout => \COUNTER.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_RNO_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__7458\,
            in1 => \N__7637\,
            in2 => \N__7519\,
            in3 => \N__7487\,
            lcout => \COUNTER.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_0_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__8569\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7619\,
            lcout => \COUNTER.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10554\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNINUSC_1_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__9502\,
            in1 => \N__9658\,
            in2 => \N__9613\,
            in3 => \N__8495\,
            lcout => \VPP_VDDQ.curr_state_2_e_0_RNINUSCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__8570\,
            in1 => \_gnd_net_\,
            in2 => \N__7642\,
            in3 => \N__7620\,
            lcout => \COUNTER.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10554\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_6_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__7489\,
            in1 => \_gnd_net_\,
            in2 => \N__7471\,
            in3 => \N__8580\,
            lcout => \COUNTER.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_RNO_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7749\,
            in1 => \N__7764\,
            in2 => \N__7783\,
            in3 => \N__7443\,
            lcout => \COUNTER.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_4_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__8577\,
            in1 => \_gnd_net_\,
            in2 => \N__7531\,
            in3 => \N__7551\,
            lcout => \COUNTER.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_5_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__8578\,
            in1 => \N__7498\,
            in2 => \_gnd_net_\,
            in3 => \N__7518\,
            lcout => \COUNTER.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_2_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7585\,
            in1 => \N__7603\,
            in2 => \_gnd_net_\,
            in3 => \N__8579\,
            lcout => \COUNTER.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10615\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_RNO_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7719\,
            in1 => \N__7686\,
            in2 => \N__7705\,
            in3 => \N__7734\,
            lcout => \COUNTER.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_RNO_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7671\,
            in1 => \N__7656\,
            in2 => \N__7894\,
            in3 => \N__7908\,
            lcout => \COUNTER.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_RNO_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7860\,
            in1 => \N__7827\,
            in2 => \N__7846\,
            in3 => \N__7875\,
            lcout => \COUNTER.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIIJV1_4_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7414\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7389\,
            lcout => \VPP_VDDQ.un9_clk_100khz_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNO_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7971\,
            in1 => \N__7956\,
            in2 => \N__7924\,
            in3 => \N__7941\,
            lcout => \COUNTER.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_RNO_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7812\,
            in1 => \N__7797\,
            in2 => \N__7990\,
            in3 => \N__8004\,
            lcout => \COUNTER.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_1_RNO_0_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8065\,
            in2 => \_gnd_net_\,
            in3 => \N__8034\,
            lcout => \RSMRST_PWRGD.curr_state10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_14_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7200\,
            in2 => \_gnd_net_\,
            in3 => \N__7051\,
            lcout => \PCH_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10454\,
            ce => \N__6962\,
            sr => \N__6793\
        );

    \PCH_PWRGD.count_10_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7016\,
            lcout => \PCH_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10454\,
            ce => \N__6962\,
            sr => \N__6793\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__10812\,
            in1 => \N__11106\,
            in2 => \N__10022\,
            in3 => \N__8241\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIES131_10_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__10274\,
            in1 => \_gnd_net_\,
            in2 => \N__6709\,
            in3 => \N__7423\,
            lcout => \VPP_VDDQ.count_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIB5TR_4_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7382\,
            in1 => \N__10271\,
            in2 => \_gnd_net_\,
            in3 => \N__7347\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNITC831_5_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10272\,
            in1 => \N__11140\,
            in2 => \_gnd_net_\,
            in3 => \N__7429\,
            lcout => \VPP_VDDQ.count_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIVF931_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__10811\,
            in1 => \N__11105\,
            in2 => \_gnd_net_\,
            in3 => \N__8276\,
            lcout => \VPP_VDDQ.count_2_1_6\,
            ltout => \VPP_VDDQ.count_2_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNID7TR_6_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__10273\,
            in1 => \_gnd_net_\,
            in2 => \N__7282\,
            in3 => \N__7413\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNI98JR5_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__9256\,
            in1 => \N__7270\,
            in2 => \N__7279\,
            in3 => \N__8277\,
            lcout => \VPP_VDDQ.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNIJCTQ_0_1_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__11107\,
            in1 => \N__8585\,
            in2 => \N__7324\,
            in3 => \N__10813\,
            lcout => \VPP_VDDQ.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__9975\,
            in1 => \N__10808\,
            in2 => \N__11060\,
            in3 => \N__8253\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI5PC31_9_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7258\,
            in2 => \N__7264\,
            in3 => \N__10205\,
            lcout => \VPP_VDDQ.count_2Z0Z_9\,
            ltout => \VPP_VDDQ.count_2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_9_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__11005\,
            in1 => \N__10810\,
            in2 => \N__7261\,
            in3 => \N__8254\,
            lcout => \VPP_VDDQ.count_2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10407\,
            ce => \N__10260\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_8_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100000000000"
        )
    port map (
            in0 => \N__10809\,
            in1 => \N__9901\,
            in2 => \N__8395\,
            in3 => \N__11004\,
            lcout => \VPP_VDDQ.count_2_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10407\,
            ce => \N__10260\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__11193\,
            in1 => \N__10807\,
            in2 => \N__11059\,
            in3 => \N__11151\,
            lcout => \VPP_VDDQ.count_2_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_10_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__8242\,
            in1 => \N__10011\,
            in2 => \N__11084\,
            in3 => \N__10840\,
            lcout => \VPP_VDDQ.count_2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10407\,
            ce => \N__10260\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI25V3_1_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7412\,
            in1 => \N__8720\,
            in2 => \N__7390\,
            in3 => \N__9228\,
            lcout => \VPP_VDDQ.count_2_RNI25V3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI82TR_1_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10729\,
            in2 => \N__11052\,
            in3 => \N__8324\,
            lcout => \VPP_VDDQ.count_2_1_1\,
            ltout => \VPP_VDDQ.count_2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNI_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7363\,
            in1 => \N__9241\,
            in2 => \N__7354\,
            in3 => \N__7351\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNILHSU_0_1_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110111111111"
        )
    port map (
            in0 => \N__7336\,
            in1 => \N__10187\,
            in2 => \N__7330\,
            in3 => \N__8416\,
            lcout => \VPP_VDDQ.m4_1\,
            ltout => \VPP_VDDQ.m4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_1_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__10730\,
            in1 => \_gnd_net_\,
            in2 => \N__7327\,
            in3 => \N__8328\,
            lcout => \VPP_VDDQ.count_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10564\,
            ce => \N__10267\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI82TR_1_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__8721\,
            in1 => \N__8566\,
            in2 => \N__7313\,
            in3 => \N__7288\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_c_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7641\,
            in2 => \N__7624\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \COUNTER.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7602\,
            in2 => \_gnd_net_\,
            in3 => \N__7579\,
            lcout => \COUNTER.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_1\,
            carryout => \COUNTER.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7576\,
            in2 => \_gnd_net_\,
            in3 => \N__7555\,
            lcout => \COUNTER.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_2\,
            carryout => \COUNTER.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7550\,
            in2 => \_gnd_net_\,
            in3 => \N__7522\,
            lcout => \COUNTER.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_3\,
            carryout => \COUNTER.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7517\,
            in2 => \_gnd_net_\,
            in3 => \N__7492\,
            lcout => \COUNTER.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_4\,
            carryout => \COUNTER.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7488\,
            in2 => \_gnd_net_\,
            in3 => \N__7462\,
            lcout => \COUNTER.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_5\,
            carryout => \COUNTER.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_7_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7459\,
            in2 => \_gnd_net_\,
            in3 => \N__7447\,
            lcout => \COUNTER.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_6\,
            carryout => \COUNTER.counter_1_cry_7\,
            clk => \N__10613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_8_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7444\,
            in2 => \_gnd_net_\,
            in3 => \N__7432\,
            lcout => \COUNTER.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_7\,
            carryout => \COUNTER.counter_1_cry_8\,
            clk => \N__10613\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_9_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7782\,
            in2 => \_gnd_net_\,
            in3 => \N__7768\,
            lcout => \COUNTER.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \COUNTER.counter_1_cry_9\,
            clk => \N__10610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_10_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7765\,
            in2 => \_gnd_net_\,
            in3 => \N__7753\,
            lcout => \COUNTER.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_9\,
            carryout => \COUNTER.counter_1_cry_10\,
            clk => \N__10610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_11_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7750\,
            in2 => \_gnd_net_\,
            in3 => \N__7738\,
            lcout => \COUNTER.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_10\,
            carryout => \COUNTER.counter_1_cry_11\,
            clk => \N__10610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_12_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7735\,
            in2 => \_gnd_net_\,
            in3 => \N__7723\,
            lcout => \COUNTER.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_11\,
            carryout => \COUNTER.counter_1_cry_12\,
            clk => \N__10610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_13_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7720\,
            in2 => \_gnd_net_\,
            in3 => \N__7708\,
            lcout => \COUNTER.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_12\,
            carryout => \COUNTER.counter_1_cry_13\,
            clk => \N__10610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_14_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7704\,
            in2 => \_gnd_net_\,
            in3 => \N__7690\,
            lcout => \COUNTER.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_13\,
            carryout => \COUNTER.counter_1_cry_14\,
            clk => \N__10610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_15_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7687\,
            in2 => \_gnd_net_\,
            in3 => \N__7675\,
            lcout => \COUNTER.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_14\,
            carryout => \COUNTER.counter_1_cry_15\,
            clk => \N__10610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_16_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7672\,
            in2 => \_gnd_net_\,
            in3 => \N__7660\,
            lcout => \COUNTER.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_15\,
            carryout => \COUNTER.counter_1_cry_16\,
            clk => \N__10610\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_17_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7657\,
            in2 => \_gnd_net_\,
            in3 => \N__7645\,
            lcout => \COUNTER.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \COUNTER.counter_1_cry_17\,
            clk => \N__10614\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_18_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7909\,
            in2 => \_gnd_net_\,
            in3 => \N__7897\,
            lcout => \COUNTER.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_17\,
            carryout => \COUNTER.counter_1_cry_18\,
            clk => \N__10614\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_19_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7893\,
            in2 => \_gnd_net_\,
            in3 => \N__7879\,
            lcout => \COUNTER.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_18\,
            carryout => \COUNTER.counter_1_cry_19\,
            clk => \N__10614\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_20_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7876\,
            in2 => \_gnd_net_\,
            in3 => \N__7864\,
            lcout => \COUNTER.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_19\,
            carryout => \COUNTER.counter_1_cry_20\,
            clk => \N__10614\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_21_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7861\,
            in2 => \_gnd_net_\,
            in3 => \N__7849\,
            lcout => \COUNTER.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_20\,
            carryout => \COUNTER.counter_1_cry_21\,
            clk => \N__10614\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_22_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7845\,
            in2 => \_gnd_net_\,
            in3 => \N__7831\,
            lcout => \COUNTER.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_21\,
            carryout => \COUNTER.counter_1_cry_22\,
            clk => \N__10614\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_23_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7828\,
            in2 => \_gnd_net_\,
            in3 => \N__7816\,
            lcout => \COUNTER.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_22\,
            carryout => \COUNTER.counter_1_cry_23\,
            clk => \N__10614\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_24_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7813\,
            in2 => \_gnd_net_\,
            in3 => \N__7801\,
            lcout => \COUNTER.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_23\,
            carryout => \COUNTER.counter_1_cry_24\,
            clk => \N__10614\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_25_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7798\,
            in2 => \_gnd_net_\,
            in3 => \N__7786\,
            lcout => \COUNTER.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \COUNTER.counter_1_cry_25\,
            clk => \N__10611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_26_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8005\,
            in2 => \_gnd_net_\,
            in3 => \N__7993\,
            lcout => \COUNTER.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_25\,
            carryout => \COUNTER.counter_1_cry_26\,
            clk => \N__10611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_27_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7989\,
            in2 => \_gnd_net_\,
            in3 => \N__7975\,
            lcout => \COUNTER.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_26\,
            carryout => \COUNTER.counter_1_cry_27\,
            clk => \N__10611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_28_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7972\,
            in2 => \_gnd_net_\,
            in3 => \N__7960\,
            lcout => \COUNTER.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_27\,
            carryout => \COUNTER.counter_1_cry_28\,
            clk => \N__10611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_29_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7957\,
            in2 => \_gnd_net_\,
            in3 => \N__7945\,
            lcout => \COUNTER.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_28\,
            carryout => \COUNTER.counter_1_cry_29\,
            clk => \N__10611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_30_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7942\,
            in2 => \_gnd_net_\,
            in3 => \N__7930\,
            lcout => \COUNTER.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_29\,
            carryout => \COUNTER.counter_1_cry_30\,
            clk => \N__10611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_31_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7923\,
            in2 => \_gnd_net_\,
            in3 => \N__7927\,
            lcout => \COUNTER.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10611\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNISEFS1_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__8118\,
            in1 => \N__8062\,
            in2 => \_gnd_net_\,
            in3 => \N__8030\,
            lcout => \RSMRST_PWRGD.un1_curr_state10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI9RLK1_3_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8787\,
            in1 => \N__8802\,
            in2 => \N__8773\,
            in3 => \N__8832\,
            lcout => \RSMRST_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI4MLK1_1_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8817\,
            in1 => \N__8847\,
            in2 => \N__9187\,
            in3 => \N__8862\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.un4_count_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIR8OP4_10_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8146\,
            in1 => \N__8206\,
            in2 => \N__8140\,
            in3 => \N__8125\,
            lcout => \RSMRST_PWRGD.N_1_i\,
            ltout => \RSMRST_PWRGD.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m5_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__8117\,
            in1 => \_gnd_net_\,
            in2 => \N__8137\,
            in3 => \N__8063\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_1_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__8064\,
            in1 => \N__8035\,
            in2 => \N__8134\,
            in3 => \N__9102\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10591\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNINN7M6_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101111"
        )
    port map (
            in0 => \N__8060\,
            in1 => \N__8031\,
            in2 => \N__8119\,
            in3 => \N__8073\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.G_10_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8131\,
            in3 => \N__9053\,
            lcout => \G_10\,
            ltout => \G_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNO_0_15_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9054\,
            in1 => \_gnd_net_\,
            in2 => \N__8128\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.N_9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNISRRR_15_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8901\,
            in1 => \N__8601\,
            in2 => \N__8884\,
            in3 => \N__9117\,
            lcout => \RSMRST_PWRGD.un4_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m3_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8113\,
            in1 => \N__8032\,
            in2 => \_gnd_net_\,
            in3 => \N__8074\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.i3_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_0_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000010101010"
        )
    port map (
            in0 => \N__8033\,
            in1 => \N__8061\,
            in2 => \N__8038\,
            in3 => \N__9055\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNIK71G1_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__9608\,
            in1 => \N__8199\,
            in2 => \N__8368\,
            in3 => \N__8308\,
            lcout => \VPP_VDDQ_delayed_vddq_ok\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIIRGK_10_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9150\,
            in1 => \N__9165\,
            in2 => \N__9136\,
            in3 => \N__8754\,
            lcout => \RSMRST_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__9601\,
            in1 => \N__8364\,
            in2 => \N__8200\,
            in3 => \N__8307\,
            lcout => \VPP_VDDQ.delayed_vddq_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10541\,
            ce => 'H',
            sr => \N__8404\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__9861\,
            in1 => \N__11053\,
            in2 => \N__10839\,
            in3 => \N__10053\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIP6631_3_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10042\,
            in2 => \N__8185\,
            in3 => \N__10270\,
            lcout => \VPP_VDDQ.count_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8698\,
            in2 => \N__8350\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_cZ0_THRU_LUT4_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9801\,
            in2 => \_gnd_net_\,
            in3 => \N__8182\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_1_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_1_cZ0\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_cZ0_THRU_LUT4_0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9862\,
            in3 => \N__8179\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_2_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_2_cZ0\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIR9731_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8176\,
            in3 => \N__8149\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIRZ0Z9731\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_3_cZ0\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_4_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_cZ0_THRU_LUT4_0_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11197\,
            in3 => \N__8293\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_4_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_4_cZ0\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIVF931_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8290\,
            in3 => \N__8263\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNIVFZ0Z931\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_5_cZ0\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNI1JA31_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9202\,
            in2 => \_gnd_net_\,
            in3 => \N__8260\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNI1JAZ0Z31\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_6_cZ0\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_cZ0_THRU_LUT4_0_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9910\,
            in3 => \N__8257\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_7_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_7_cZ0\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_cZ0_THRU_LUT4_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9964\,
            in2 => \_gnd_net_\,
            in3 => \N__8245\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_8_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_THRU_LUT4_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10018\,
            in3 => \N__8230\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_THRU_LUT4_0_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9937\,
            in3 => \N__8227\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_THRU_LUT4_0_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10885\,
            in3 => \N__8224\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_THRU_LUT4_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9764\,
            in3 => \N__8221\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_THRU_LUT4_0_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9713\,
            in3 => \N__8410\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_THRU_LUT4_0_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8407\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__9946\,
            in1 => \N__11015\,
            in2 => \N__10846\,
            in3 => \N__9276\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNO_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__10780\,
            in1 => \N__8505\,
            in2 => \N__9500\,
            in3 => \N__9594\,
            lcout => \VPP_VDDQ.delayed_vddq_ok_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__11014\,
            in1 => \N__10777\,
            in2 => \N__9909\,
            in3 => \N__8394\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI3MB31_8_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8377\,
            in2 => \N__8371\,
            in3 => \N__10204\,
            lcout => \VPP_VDDQ.count_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNI8PF7_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9486\,
            in1 => \_gnd_net_\,
            in2 => \N__9606\,
            in3 => \N__10778\,
            lcout => \VPP_VDDQ.un1_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI82TR_0_1_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8346\,
            in2 => \_gnd_net_\,
            in3 => \N__8697\,
            lcout => \VPP_VDDQ.count_2_RNI82TR_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNIJCTQ_1_1_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__9487\,
            in1 => \N__9445\,
            in2 => \N__9607\,
            in3 => \N__10779\,
            lcout => \VPP_VDDQ.delayed_vddq_ok_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI8PF7_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9587\,
            in2 => \_gnd_net_\,
            in3 => \N__9485\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_en_0_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNIJCTQ_1_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__8504\,
            in1 => \N__9641\,
            in2 => \N__8590\,
            in3 => \N__8581\,
            lcout => \VPP_VDDQ.count_2_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_2_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9900\,
            in2 => \_gnd_net_\,
            in3 => \N__9794\,
            lcout => \VPP_VDDQ.g0_2_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNISBBC7_0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8623\,
            in2 => \N__8506\,
            in3 => \N__9664\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_0_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8512\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.curr_state_2_RNIZ0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2_RNIZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m6_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__9652\,
            in1 => \N__9573\,
            in2 => \N__8509\,
            in3 => \N__11030\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.m6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNIIOCG_1_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8502\,
            in2 => \N__8422\,
            in3 => \N__9454\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_1\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_RNI_1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8419\,
            in3 => \N__9484\,
            lcout => \VPP_VDDQ.un5_clk_100khz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_0_2_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__9826\,
            in1 => \N__8696\,
            in2 => \_gnd_net_\,
            in3 => \N__9793\,
            lcout => \VPP_VDDQ.count_2_RNI_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_0_10_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__9863\,
            in1 => \N__9974\,
            in2 => \N__10030\,
            in3 => \N__9945\,
            lcout => \VPP_VDDQ.g0_2_a2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNILHSU_1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9229\,
            in1 => \N__8740\,
            in2 => \N__8731\,
            in3 => \N__10231\,
            lcout => \VPP_VDDQ.N_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_0_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__10728\,
            in1 => \N__8695\,
            in2 => \_gnd_net_\,
            in3 => \N__11051\,
            lcout => \VPP_VDDQ.count_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10631\,
            ce => \N__10269\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_1_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10727\,
            in2 => \_gnd_net_\,
            in3 => \N__11034\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.g0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI71TR_0_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__10230\,
            in1 => \N__8707\,
            in2 => \N__8701\,
            in3 => \N__8694\,
            lcout => \VPP_VDDQ.count_2Z0Z_0\,
            ltout => \VPP_VDDQ.count_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_5_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8665\,
            in1 => \N__8659\,
            in2 => \N__8653\,
            in3 => \N__11205\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.g0_2_a2_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIUPFQ6_1_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__8650\,
            in1 => \N__8641\,
            in2 => \N__8629\,
            in3 => \N__9688\,
            lcout => \VPP_VDDQ.count_2_RNIUPFQ6Z0Z_1\,
            ltout => \VPP_VDDQ.count_2_RNIUPFQ6Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__9580\,
            in1 => \N__9682\,
            in2 => \N__8626\,
            in3 => \N__9656\,
            lcout => \VPP_VDDQ.m4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9098\,
            in1 => \N__8602\,
            in2 => \N__8617\,
            in3 => \N__8616\,
            lcout => \RSMRST_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_0\,
            clk => \N__10592\,
            ce => 'H',
            sr => \N__9309\
        );

    \RSMRST_PWRGD.count_1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9094\,
            in1 => \N__8863\,
            in2 => \_gnd_net_\,
            in3 => \N__8851\,
            lcout => \RSMRST_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_0\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_1\,
            clk => \N__10592\,
            ce => 'H',
            sr => \N__9309\
        );

    \RSMRST_PWRGD.count_2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9099\,
            in1 => \N__8848\,
            in2 => \_gnd_net_\,
            in3 => \N__8836\,
            lcout => \RSMRST_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_1\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_2\,
            clk => \N__10592\,
            ce => 'H',
            sr => \N__9309\
        );

    \RSMRST_PWRGD.count_3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9095\,
            in1 => \N__8833\,
            in2 => \_gnd_net_\,
            in3 => \N__8821\,
            lcout => \RSMRST_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_2\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_3\,
            clk => \N__10592\,
            ce => 'H',
            sr => \N__9309\
        );

    \RSMRST_PWRGD.count_4_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9100\,
            in1 => \N__8818\,
            in2 => \_gnd_net_\,
            in3 => \N__8806\,
            lcout => \RSMRST_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_3\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_4\,
            clk => \N__10592\,
            ce => 'H',
            sr => \N__9309\
        );

    \RSMRST_PWRGD.count_5_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9096\,
            in1 => \N__8803\,
            in2 => \_gnd_net_\,
            in3 => \N__8791\,
            lcout => \RSMRST_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_4\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_5\,
            clk => \N__10592\,
            ce => 'H',
            sr => \N__9309\
        );

    \RSMRST_PWRGD.count_6_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9101\,
            in1 => \N__8788\,
            in2 => \_gnd_net_\,
            in3 => \N__8776\,
            lcout => \RSMRST_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_5\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_6\,
            clk => \N__10592\,
            ce => 'H',
            sr => \N__9309\
        );

    \RSMRST_PWRGD.count_7_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9097\,
            in1 => \N__8772\,
            in2 => \_gnd_net_\,
            in3 => \N__8758\,
            lcout => \RSMRST_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_6\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_7\,
            clk => \N__10592\,
            ce => 'H',
            sr => \N__9309\
        );

    \RSMRST_PWRGD.count_8_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9080\,
            in1 => \N__8755\,
            in2 => \_gnd_net_\,
            in3 => \N__8743\,
            lcout => \RSMRST_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_8\,
            clk => \N__10546\,
            ce => 'H',
            sr => \N__9297\
        );

    \RSMRST_PWRGD.count_9_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9076\,
            in1 => \N__9183\,
            in2 => \_gnd_net_\,
            in3 => \N__9169\,
            lcout => \RSMRST_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_8\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_9\,
            clk => \N__10546\,
            ce => 'H',
            sr => \N__9297\
        );

    \RSMRST_PWRGD.count_10_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9077\,
            in1 => \N__9166\,
            in2 => \_gnd_net_\,
            in3 => \N__9154\,
            lcout => \RSMRST_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_9\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_10\,
            clk => \N__10546\,
            ce => 'H',
            sr => \N__9297\
        );

    \RSMRST_PWRGD.count_11_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9074\,
            in1 => \N__9151\,
            in2 => \_gnd_net_\,
            in3 => \N__9139\,
            lcout => \RSMRST_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_10\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_11\,
            clk => \N__10546\,
            ce => 'H',
            sr => \N__9297\
        );

    \RSMRST_PWRGD.count_12_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9078\,
            in1 => \N__9135\,
            in2 => \_gnd_net_\,
            in3 => \N__9121\,
            lcout => \RSMRST_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_11\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_12\,
            clk => \N__10546\,
            ce => 'H',
            sr => \N__9297\
        );

    \RSMRST_PWRGD.count_13_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9075\,
            in1 => \N__9118\,
            in2 => \_gnd_net_\,
            in3 => \N__9106\,
            lcout => \RSMRST_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_12\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_13\,
            clk => \N__10546\,
            ce => 'H',
            sr => \N__9297\
        );

    \RSMRST_PWRGD.count_14_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9079\,
            in1 => \N__8902\,
            in2 => \_gnd_net_\,
            in3 => \N__8890\,
            lcout => \RSMRST_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_13\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14\,
            clk => \N__10546\,
            ce => 'H',
            sr => \N__9297\
        );

    \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10113\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_14\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_15_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8883\,
            in2 => \_gnd_net_\,
            in3 => \N__8887\,
            lcout => \RSMRST_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10593\,
            ce => \N__8869\,
            sr => \N__9313\
        );

    \VPP_VDDQ.count_2_RNINQ791_11_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9262\,
            in1 => \N__10276\,
            in2 => \_gnd_net_\,
            in3 => \N__9283\,
            lcout => \VPP_VDDQ.count_2Z0Z_11\,
            ltout => \VPP_VDDQ.count_2Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_11_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__9277\,
            in1 => \N__11101\,
            in2 => \N__9265\,
            in3 => \N__10819\,
            lcout => \VPP_VDDQ.count_2_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10618\,
            ce => \N__10282\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_7_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__10818\,
            in1 => \_gnd_net_\,
            in2 => \N__11115\,
            in3 => \N__9255\,
            lcout => \VPP_VDDQ.count_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10618\,
            ce => \N__10282\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIPT891_12_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10645\,
            in2 => \N__9196\,
            in3 => \N__10277\,
            lcout => \VPP_VDDQ.count_2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNI1JA31_0_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9254\,
            in1 => \N__11100\,
            in2 => \_gnd_net_\,
            in3 => \N__10817\,
            lcout => \VPP_VDDQ.count_2_1_7\,
            ltout => \VPP_VDDQ.count_2_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIE8TR_7_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9221\,
            in2 => \N__9205\,
            in3 => \N__10275\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__10884\,
            in1 => \N__11088\,
            in2 => \N__10847\,
            in3 => \N__11127\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_15_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000010000000"
        )
    port map (
            in0 => \N__10850\,
            in1 => \N__9343\,
            in2 => \N__11114\,
            in3 => \N__9737\,
            lcout => \VPP_VDDQ.count_2_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10625\,
            ce => \N__10280\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__9712\,
            in1 => \N__11092\,
            in2 => \N__10848\,
            in3 => \N__9378\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIT3B91_14_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__10207\,
            in1 => \_gnd_net_\,
            in2 => \N__9385\,
            in3 => \N__9370\,
            lcout => \VPP_VDDQ.count_2Z0Z_14\,
            ltout => \VPP_VDDQ.count_2Z0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_14_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__10828\,
            in1 => \N__11093\,
            in2 => \N__9382\,
            in3 => \N__9379\,
            lcout => \VPP_VDDQ.count_2_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10625\,
            ce => \N__10280\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__9763\,
            in1 => \N__10823\,
            in2 => \N__11113\,
            in3 => \N__9357\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIR0A91_13_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9349\,
            in2 => \N__9364\,
            in3 => \N__10206\,
            lcout => \VPP_VDDQ.count_2Z0Z_13\,
            ltout => \VPP_VDDQ.count_2Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_13_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__11094\,
            in1 => \N__10827\,
            in2 => \N__9361\,
            in3 => \N__9358\,
            lcout => \VPP_VDDQ.count_2_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10625\,
            ce => \N__10280\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__9738\,
            in1 => \N__11078\,
            in2 => \N__10829\,
            in3 => \N__9342\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIV6C91_15_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9331\,
            in2 => \N__9325\,
            in3 => \N__10186\,
            lcout => \VPP_VDDQ.count_2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIN3531_2_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9319\,
            in2 => \N__9775\,
            in3 => \N__10185\,
            lcout => \VPP_VDDQ.count_2Z0Z_2\,
            ltout => \VPP_VDDQ.count_2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_2_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__9816\,
            in1 => \N__11079\,
            in2 => \N__9322\,
            in3 => \N__10793\,
            lcout => \VPP_VDDQ.count_2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10612\,
            ce => \N__10268\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_3_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100000000000"
        )
    port map (
            in0 => \N__10792\,
            in1 => \N__9864\,
            in2 => \N__10063\,
            in3 => \N__11083\,
            lcout => \VPP_VDDQ.count_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10612\,
            ce => \N__10268\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_15_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9736\,
            in1 => \N__9766\,
            in2 => \N__10893\,
            in3 => \N__9715\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.N_1_i_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_10_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10029\,
            in1 => \N__9979\,
            in2 => \N__9949\,
            in3 => \N__9944\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un9_clk_100khz_14_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_3_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__11206\,
            in1 => \N__9905\,
            in2 => \N__9871\,
            in3 => \N__9868\,
            lcout => \VPP_VDDQ.count_2_RNIZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000000000"
        )
    port map (
            in0 => \N__11116\,
            in1 => \N__9820\,
            in2 => \N__9802\,
            in3 => \N__10726\,
            lcout => \VPP_VDDQ.count_2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_0_15_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10886\,
            in1 => \N__9765\,
            in2 => \N__9739\,
            in3 => \N__9714\,
            lcout => \VPP_VDDQ.g0_2_a2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011100000001000"
        )
    port map (
            in0 => \N__9551\,
            in1 => \N__9681\,
            in2 => \N__9657\,
            in3 => \N__9670\,
            lcout => \VPP_VDDQ.curr_state_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10632\,
            ce => \N__9448\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_e_0_1_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__9648\,
            in1 => \N__9552\,
            in2 => \N__9501\,
            in3 => \N__11108\,
            lcout => \VPP_VDDQ.curr_state_2_e_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10632\,
            ce => \N__9448\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_5_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__11201\,
            in1 => \N__11109\,
            in2 => \N__11158\,
            in3 => \N__10851\,
            lcout => \VPP_VDDQ.count_2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10608\,
            ce => \N__10281\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_12_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__11131\,
            in1 => \N__11098\,
            in2 => \N__10897\,
            in3 => \N__10849\,
            lcout => \VPP_VDDQ.count_2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10493\,
            ce => \N__10279\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
